-- Version: 7.3 7.3.0.29

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity PDL_INTERF is

    port( PULSE         : in    std_logic_vector(8 to 8);
          P_PDL_c       : out   std_logic_vector(7 downto 1);
          PDL_RDATA     : out   std_logic_vector(7 downto 0);
          PDL_RADDR     : in    std_logic_vector(5 downto 0);
          PDLCFG_RAD    : out   std_logic_vector(5 downto 0);
          PDLCFG_DT     : in    std_logic_vector(7 downto 0);
          PDLCFG_DT_0_0 : in    std_logic_vector(0 to 0);
          PDLCFG_DT_3   : in    std_logic_vector(0 to 0);
          PDLCFG_DT_1   : in    std_logic_vector(0 to 0);
          PDLCFG_DT_2   : in    std_logic_vector(0 to 0);
          PDLCFG_DT_0   : in    std_logic_vector(0 to 0);
          P0            : out   std_logic_vector(47 downto 0);
          AE_PDL_c      : out   std_logic_vector(47 downto 0);
          SP_PDL_in     : in    std_logic_vector(47 downto 0);
          REG_0         : in    std_logic_vector(127 downto 124);
          REG_i_0       : in    std_logic_vector(121 to 121);
          REG_32        : in    std_logic;
          REG_33        : in    std_logic;
          REG_34        : in    std_logic;
          REG_35        : in    std_logic;
          REG_36        : in    std_logic;
          REG_37        : in    std_logic;
          REG_38        : in    std_logic;
          REG_39        : in    std_logic;
          REG_40        : in    std_logic;
          REG_41        : in    std_logic;
          REG_42        : in    std_logic;
          REG_43        : in    std_logic;
          REG_44        : in    std_logic;
          REG_45        : in    std_logic;
          REG_46        : in    std_logic;
          REG_47        : in    std_logic;
          REG_48        : in    std_logic;
          REG_49        : in    std_logic;
          REG_50        : in    std_logic;
          REG_51        : in    std_logic;
          REG_52        : in    std_logic;
          REG_53        : in    std_logic;
          REG_54        : in    std_logic;
          REG_55        : in    std_logic;
          REG_56        : in    std_logic;
          REG_57        : in    std_logic;
          REG_58        : in    std_logic;
          REG_59        : in    std_logic;
          REG_60        : in    std_logic;
          REG_61        : in    std_logic;
          REG_62        : in    std_logic;
          REG_63        : in    std_logic;
          REG_64        : in    std_logic;
          REG_65        : in    std_logic;
          REG_66        : in    std_logic;
          REG_67        : in    std_logic;
          REG_68        : in    std_logic;
          REG_69        : in    std_logic;
          REG_70        : in    std_logic;
          REG_71        : in    std_logic;
          REG_72        : in    std_logic;
          REG_73        : in    std_logic;
          REG_74        : in    std_logic;
          REG_75        : in    std_logic;
          REG_76        : in    std_logic;
          REG_77        : in    std_logic;
          REG_78        : in    std_logic;
          REG_79        : in    std_logic;
          REG_3         : in    std_logic;
          REG_6         : in    std_logic;
          REG_5         : in    std_logic;
          REG_4         : in    std_logic;
          REG_2         : in    std_logic;
          REG_1         : in    std_logic;
          REG_24        : out   std_logic;
          REG_9         : in    std_logic;
          REG_16        : out   std_logic;
          REG_10        : in    std_logic;
          REG_17        : out   std_logic;
          REG_11        : in    std_logic;
          REG_18        : out   std_logic;
          REG_12        : in    std_logic;
          REG_19        : out   std_logic;
          REG_13        : in    std_logic;
          REG_20        : out   std_logic;
          REG_14        : in    std_logic;
          REG_21        : out   std_logic;
          REG_15        : in    std_logic;
          REG_22        : out   std_logic;
          REG_23        : out   std_logic;
          REG_0_d0      : in    std_logic;
          REG_8         : in    std_logic;
          MD_PDL_c      : out   std_logic;
          PDL_RACK      : out   std_logic;
          PDL_RREQ      : in    std_logic;
          SI_PDL_c      : out   std_logic;
          PDLCFG_nRD    : out   std_logic;
          SCLK_PDL_c    : out   std_logic;
          HWRES_c_2     : in    std_logic;
          HWRES_c_1     : in    std_logic;
          MD_PDL_c_0    : out   std_logic;
          MD_PDL_c_1    : out   std_logic;
          MD_PDL_c_2    : out   std_logic;
          MD_PDL_c_3    : out   std_logic;
          LOAD_RES      : in    std_logic;
          HWRES_c_0_3   : in    std_logic;
          HWRES_c_0_2   : in    std_logic;
          LOAD_RES_3    : in    std_logic;
          CLK_c_c       : in    std_logic;
          HWRES_c_23_0  : in    std_logic;
          HWRES_c_0     : in    std_logic;
          LOAD_RES_0    : in    std_logic
        );

end PDL_INTERF;

architecture DEF_ARCH of PDL_INTERF is 

  component NAND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NAND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OAI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \un1_load_res_0_0\, \sstate_2[6]_net_1\, 
        un2_load_res_i, \sstate_19_1[6]\, \sstate_1[6]_net_1\, 
        \sstate_0[6]_net_1\, \sstate_8[9]_net_1\, 
        \sstate[10]_net_1\, \sstate_7[9]_net_1\, 
        \sstate_6[9]_net_1\, \sstate_5[9]_net_1\, 
        \sstate_4[9]_net_1\, \sstate_3[9]_net_1\, 
        \sstate_2[9]_net_1\, \sstate_1[9]_net_1\, 
        \sstate_0[9]_net_1\, \un1_load_res\, \un1_load_res_11\, 
        \un1_load_res_10\, \un1_load_res_9\, \un1_load_res_8\, 
        \un1_load_res_7\, \un1_load_res_6\, \un1_load_res_5\, 
        \un1_load_res_4\, \un1_load_res_3\, \un1_load_res_2\, 
        \un1_load_res_1\, \un1_load_res_0\, un1_hwres_1_i, 
        \un1_reg_1_i\, \MODE_0\, \AE_1_sqmuxa_2\, \MD_PDL_c_0\, 
        \AE_1_sqmuxa_1\, \AE_1_sqmuxa_0\, \un1_sstate_2_3\, 
        \un1_sstate_2_2\, \un1_sstate_2_1\, \un1_sstate_2_0\, 
        \un1_sstate_14_2\, \un1_sstate_5\, \sstate[11]_net_1\, 
        \un1_sstate_14_1\, \un1_sstate_14_0\, \REG_m_i_2[129]\, 
        \REG_m_i_1[129]\, \REG_m_i_0[129]\, AE_0_sqmuxa_i_2, 
        AE_0_sqmuxa_i_1, AE_0_sqmuxa_i_0, N_6864_2, 
        \sstate[12]_net_1\, N_6864_1, N_6864_0, 
        \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \BITCNT[1]_net_1\, \DWACT_ADD_CI_0_TMP_0[0]\, 
        \CNT[1]_net_1\, \DWACT_ADD_CI_0_g_array_12_1[0]\, 
        \CNT[4]_net_1\, \DWACT_ADD_CI_0_g_array_12[0]\, 
        \CNT[2]_net_1\, LOAD_RES_i_0, un1_reg_1_i_i, 
        \PDLCFG_RAD_0_sqmuxa_1_i\, \PDLCFG_RAD_0_sqmuxa_1\, 
        \sstate_19_1[11]_net_1\, \sstate[8]_net_1\, \SBYTE_136\, 
        \SBYTE_5[7]_net_1\, \un1_sstate_20\, \SBYTE_135\, 
        \SBYTE_5[6]_net_1\, \REG[143]\, \SBYTE_134\, 
        \SBYTE_5[5]_net_1\, \REG[142]\, \SBYTE_133\, 
        \SBYTE_5[4]_net_1\, \REG[141]\, \SBYTE_132\, 
        \SBYTE_5[3]_net_1\, \REG[140]\, \SBYTE_131\, 
        \SBYTE_5[2]_net_1\, \REG[139]\, \SBYTE_130\, 
        \SBYTE_5[1]_net_1\, \REG[138]\, \SBYTE_129\, 
        \SBYTE_5[0]_net_1\, \REG[137]\, \sstate[3]_net_1\, 
        \ISI_1_sqmuxa_1\, \SO\, un4_so, N_474, N_497, N_462, 
        N_473, N_456_i, N_461_i, N_456_i_i, N_453, N_458, N_452, 
        N_457, N_461_i_i, N_455, N_460, N_454, N_459, N_467_i, 
        N_472_i, N_467_i_i, N_464, N_469, N_463, N_468, N_472_i_i, 
        N_466, N_471, N_465, N_470, N_485, N_496, N_479_i, 
        N_484_i, N_479_i_i, N_476, N_481, N_475, N_480, N_484_i_i, 
        N_478, N_483, N_477, N_482, N_490_i, N_495_i, N_490_i_i, 
        N_487, N_492, N_486, N_491, N_495_i_i, N_489, N_494, 
        N_488, N_493, \ISCK_128\, \un1_sstate_13\, \un1_sstate_1\, 
        \un1_sstate_13_0\, \sstate[2]_net_1\, \AE_127\, 
        \AE_7[47]\, \AE_i_m[47]_net_1\, \REG_i_m[200]_net_1\, 
        \AE_0_sqmuxa_188\, \AE_0_sqmuxa_190\, \AE_PDL_c[47]\, 
        \un69_ae_3[47]\, \un69_ae_4[47]\, \AE_126\, \AE_7[46]\, 
        \AE_i_m[46]_net_1\, \REG_i_m[199]_net_1\, 
        \AE_0_sqmuxa_184\, \AE_0_sqmuxa_186\, \AE_PDL_c[46]\, 
        \un69_ae_1[38]\, \AE_125\, \AE_7[45]\, \AE_i_m[45]_net_1\, 
        \REG_i_m[198]_net_1\, \AE_0_sqmuxa_180\, 
        \AE_0_sqmuxa_182\, \AE_PDL_c[45]\, un69_ae_37_0, \AE_124\, 
        \AE_7[44]\, \AE_i_m[44]_net_1\, \REG_i_m[197]_net_1\, 
        \AE_0_sqmuxa_176\, \AE_0_sqmuxa_178\, \AE_PDL_c[44]\, 
        \un69_ae_1[44]\, \AE_123\, \AE_7[43]\, \AE_i_m[43]_net_1\, 
        \REG_i_m[196]_net_1\, \AE_0_sqmuxa_172\, 
        \AE_0_sqmuxa_174\, \AE_PDL_c[43]\, \un69_ae_2[43]\, 
        \AE_122\, \AE_7[42]\, \AE_i_m[42]_net_1\, 
        \REG_i_m[195]_net_1\, \AE_0_sqmuxa_168\, 
        \AE_0_sqmuxa_170\, \AE_PDL_c[42]\, \un69_ae_1[42]\, 
        \AE_121\, \AE_7[41]\, \AE_i_m[41]_net_1\, 
        \REG_i_m[194]_net_1\, \AE_0_sqmuxa_164\, 
        \AE_0_sqmuxa_166\, \AE_PDL_c[41]\, \un69_ae_1[33]\, 
        \AE_120\, \AE_7[40]\, \AE_i_m[40]_net_1\, 
        \REG_i_m[193]_net_1\, \AE_0_sqmuxa_160\, 
        \AE_0_sqmuxa_162\, \AE_PDL_c[40]\, \un69_ae_1[40]\, 
        \AE_119\, \AE_7[39]\, \AE_i_m[39]_net_1\, 
        \REG_i_m[192]_net_1\, \AE_0_sqmuxa_156\, 
        \AE_0_sqmuxa_158\, \AE_PDL_c[39]\, \un69_ae_1[39]\, 
        \un69_ae_1_i[47]\, \un69_ae_2[47]\, \AE_118\, \AE_7[38]\, 
        \AE_i_m[38]_net_1\, \REG_i_m[191]_net_1\, 
        \AE_0_sqmuxa_152\, \AE_0_sqmuxa_154\, \AE_PDL_c[38]\, 
        \un69_ae_1_i[46]\, \AE_117\, \AE_7[37]\, 
        \AE_i_m[37]_net_1\, \REG_i_m[190]_net_1\, 
        \AE_0_sqmuxa_148\, \AE_0_sqmuxa_150\, \AE_PDL_c[37]\, 
        \un69_ae_1[45]\, \AE_116\, \AE_7[36]\, \AE_i_m[36]_net_1\, 
        \REG_i_m[189]_net_1\, \AE_0_sqmuxa_144\, 
        \AE_0_sqmuxa_146\, \AE_PDL_c[36]\, \AE_115\, \AE_7[35]\, 
        \AE_i_m[35]_net_1\, \REG_i_m[188]_net_1\, 
        \AE_0_sqmuxa_140\, \AE_0_sqmuxa_142\, \AE_PDL_c[35]\, 
        \un69_ae_1[43]\, \AE_114\, \AE_7[34]\, \AE_i_m[34]_net_1\, 
        \REG_i_m[187]_net_1\, \AE_0_sqmuxa_136\, 
        \AE_0_sqmuxa_138\, \AE_PDL_c[34]\, \AE_113\, \AE_7[33]\, 
        \AE_i_m[33]_net_1\, \REG_i_m[186]_net_1\, 
        \AE_0_sqmuxa_132\, \AE_0_sqmuxa_134\, \AE_PDL_c[33]\, 
        \un69_ae_1[41]\, \AE_112\, \AE_7[32]\, \AE_i_m[32]_net_1\, 
        \REG_i_m[185]_net_1\, \AE_0_sqmuxa_128\, 
        \AE_0_sqmuxa_130\, \AE_PDL_c[32]\, \AE_111\, \AE_7[31]\, 
        \AE_i_m[31]_net_1\, \REG_i_m[184]_net_1\, 
        \AE_0_sqmuxa_124\, \AE_0_sqmuxa_126\, \AE_PDL_c[31]\, 
        \un69_ae_2[31]\, \un69_ae_3[31]\, \AE_110\, \AE_7[30]\, 
        \AE_i_m[30]_net_1\, \REG_i_m[183]_net_1\, 
        \AE_0_sqmuxa_120\, \AE_0_sqmuxa_122\, \AE_PDL_c[30]\, 
        un69_ae_30_0, \AE_109\, \AE_7[29]\, \AE_i_m[29]_net_1\, 
        \REG_i_m[182]_net_1\, \AE_0_sqmuxa_116\, 
        \AE_0_sqmuxa_118\, \AE_PDL_c[29]\, \un69_ae_1[29]\, 
        \AE_108\, \AE_7[28]\, \AE_i_m[28]_net_1\, 
        \REG_i_m[181]_net_1\, \AE_0_sqmuxa_112\, 
        \AE_0_sqmuxa_114\, \AE_PDL_c[28]\, \un69_ae_1[28]\, 
        \AE_107\, \AE_7[27]\, \AE_i_m[27]_net_1\, 
        \REG_i_m[180]_net_1\, \AE_0_sqmuxa_108\, 
        \AE_0_sqmuxa_110\, \AE_PDL_c[27]\, \un69_ae_1[27]\, 
        \AE_106\, \AE_7[26]\, \AE_i_m[26]_net_1\, 
        \REG_i_m[179]_net_1\, \AE_0_sqmuxa_104\, 
        \AE_0_sqmuxa_106\, \AE_PDL_c[26]\, \un69_ae_1[26]\, 
        \AE_105\, \AE_7[25]\, \AE_i_m[25]_net_1\, 
        \REG_i_m[178]_net_1\, \AE_0_sqmuxa_100\, 
        \AE_0_sqmuxa_102\, \AE_PDL_c[25]\, \un69_ae_1[25]\, 
        \AE_104\, \AE_7[24]\, \AE_i_m[24]_net_1\, 
        \REG_i_m[177]_net_1\, \AE_0_sqmuxa_96\, \AE_0_sqmuxa_98\, 
        \AE_PDL_c[24]\, \un69_ae_1[24]\, \AE_103\, \AE_7[23]\, 
        \AE_i_m[23]_net_1\, \REG_i_m[176]_net_1\, 
        \AE_0_sqmuxa_92\, \AE_0_sqmuxa_94\, \AE_PDL_c[23]\, 
        \un69_ae_1[23]\, \un69_ae_1_i[31]\, \AE_102\, \AE_7[22]\, 
        \AE_i_m[22]_net_1\, \REG_i_m[175]_net_1\, 
        \AE_0_sqmuxa_88\, \AE_0_sqmuxa_90\, \AE_PDL_c[22]\, 
        \un69_ae_1_i[30]\, \AE_101\, \AE_7[21]\, 
        \AE_i_m[21]_net_1\, \REG_i_m[174]_net_1\, 
        \AE_0_sqmuxa_84\, \AE_0_sqmuxa_86\, \AE_PDL_c[21]\, 
        \AE_100\, \AE_7[20]\, \AE_i_m[20]_net_1\, 
        \REG_i_m[173]_net_1\, \AE_0_sqmuxa_80\, \AE_0_sqmuxa_82\, 
        \AE_PDL_c[20]\, \AE_99\, \AE_7[19]\, \AE_i_m[19]_net_1\, 
        \REG_i_m[172]_net_1\, \AE_0_sqmuxa_76\, \AE_0_sqmuxa_78\, 
        \AE_PDL_c[19]\, \AE_98\, \AE_7[18]\, \AE_i_m[18]_net_1\, 
        \REG_i_m[171]_net_1\, \AE_0_sqmuxa_72\, \AE_0_sqmuxa_74\, 
        \AE_PDL_c[18]\, \AE_1_sqmuxa\, \AE_97\, \AE_7[17]\, 
        \AE_i_m[17]_net_1\, \REG_i_m[170]_net_1\, 
        \AE_0_sqmuxa_68\, \AE_0_sqmuxa_70\, \AE_PDL_c[17]\, 
        \AE_96\, \AE_7[16]\, \AE_i_m[16]_net_1\, 
        \REG_i_m[169]_net_1\, \AE_0_sqmuxa_64\, \AE_0_sqmuxa_66\, 
        \AE_PDL_c[16]\, \AE_95\, \AE_7[15]\, \AE_i_m[15]_net_1\, 
        \REG_i_m[168]_net_1\, \AE_0_sqmuxa_60\, \AE_0_sqmuxa_62\, 
        \AE_PDL_c[15]\, \un69_ae_2[7]\, \un69_ae_2[15]\, \AE_94\, 
        \AE_7[14]\, \AE_i_m[14]_net_1\, \REG_i_m[167]_net_1\, 
        \AE_0_sqmuxa_56\, \AE_0_sqmuxa_58\, \AE_PDL_c[14]\, 
        \un69_ae_1[14]\, \AE_93\, \AE_7[13]\, \AE_i_m[13]_net_1\, 
        \REG_i_m[166]_net_1\, \AE_0_sqmuxa_52\, \AE_0_sqmuxa_54\, 
        \AE_PDL_c[13]\, \un69_ae_13_0\, \un69_ae_1[15]\, \AE_92\, 
        \AE_7[12]\, \AE_i_m[12]_net_1\, \REG_i_m[165]_net_1\, 
        \AE_0_sqmuxa_48\, \AE_0_sqmuxa_50\, \AE_PDL_c[12]\, 
        \un69_ae_12_0\, \AE_91\, \AE_7[11]\, \un1_sstate_14\, 
        \AE_i_m[11]_net_1\, \REG_i_m[164]_net_1\, 
        \AE_7_r_i[47]_net_1\, AE_0_sqmuxa_i, \AE_0_sqmuxa_44\, 
        \AE_0_sqmuxa_46\, \AE_PDL_c[11]\, \un69_ae_1[11]\, 
        \AE_90\, \AE_7[10]\, \AE_i_m[10]_net_1\, 
        \REG_i_m[163]_net_1\, \AE_0_sqmuxa_40\, \AE_0_sqmuxa_42\, 
        \AE_PDL_c[10]\, \AE_89\, \AE_7[9]\, \AE_i_m[9]_net_1\, 
        \REG_i_m[162]_net_1\, \AE_0_sqmuxa_36\, \AE_0_sqmuxa_38\, 
        \AE_PDL_c[9]\, \un69_ae_1[9]\, \AE_88\, \AE_7[8]\, 
        \AE_i_m[8]_net_1\, \REG_i_m[161]_net_1\, \AE_0_sqmuxa_32\, 
        \AE_0_sqmuxa_34\, \AE_PDL_c[8]\, \AE_87\, \AE_7[7]\, 
        \AE_i_m[7]_net_1\, \REG_i_m[160]_net_1\, \AE_0_sqmuxa_28\, 
        \AE_0_sqmuxa_30\, \AE_PDL_c[7]\, \un69_ae_1[7]\, \AE_86\, 
        \AE_7[6]\, \AE_i_m[6]_net_1\, \REG_i_m[159]_net_1\, 
        \AE_0_sqmuxa_24\, \AE_0_sqmuxa_26\, \AE_PDL_c[6]\, 
        \un69_ae_1[6]\, \AE_85\, \AE_7[5]\, \AE_i_m[5]_net_1\, 
        \REG_i_m[158]_net_1\, \AE_0_sqmuxa_20\, \AE_0_sqmuxa_22\, 
        \AE_PDL_c[5]\, \un69_ae_1[5]\, \AE_84\, \AE_7[4]\, 
        \AE_i_m[4]_net_1\, \REG_i_m[157]_net_1\, \AE_0_sqmuxa_16\, 
        \AE_0_sqmuxa_18\, \AE_PDL_c[4]\, \un69_ae_1[4]\, \AE_83\, 
        \AE_7[3]\, \AE_i_m[3]_net_1\, \REG_i_m[156]_net_1\, 
        \AE_0_sqmuxa_12\, \AE_0_sqmuxa_14\, \AE_PDL_c[3]\, 
        \AE_82\, \AE_7[2]\, \AE_i_m[2]_net_1\, 
        \REG_i_m[155]_net_1\, \AE_0_sqmuxa_8\, \AE_0_sqmuxa_10\, 
        \AE_PDL_c[2]\, \AE_81\, \AE_7[1]\, \AE_i_m[1]_net_1\, 
        \REG_i_m[154]_net_1\, \AE_0_sqmuxa_4\, \AE_0_sqmuxa_6\, 
        \AE_PDL_c[1]\, \AE_80\, \AE_7[0]\, \AE_i_m[0]_net_1\, 
        \REG_i_m[153]_net_1\, \AE_0_sqmuxa_0\, \AE_0_sqmuxa_2\, 
        \AE_PDL_c[0]\, \un69_ae_0_0\, \PDLCFG_nRD_79\, 
        \un1_sstate_29_1\, \un1_sstate_27\, un1_sstate_27_2_i, 
        un1_sstate_27_3_i, \sstate[1]_net_1\, \sstate_i_i[0]\, 
        un1_sstate_27_0_i, \sstate_i[7]\, \PDLCFG_RAD_0_sqmuxa\, 
        \ISI_78\, ISI_5, \un1_sstate_18\, \ISI_0_sqmuxa\, 
        \REG_m_i[136]\, \SBYTE_m_i[7]\, \un1_sstate_22\, 
        \REG[144]\, \P0_77\, \P0_50[47]\, \P0_m_i[47]\, 
        \PDLCFG_DT_m_7[0]_net_1\, \P0[47]_net_1\, \un3_ae[47]\, 
        \un3_ae_3[47]\, \un3_ae_4[47]\, \P0_76\, \P0_50[46]\, 
        \P0_m_i[46]\, \PDLCFG_DT_m_6[0]_net_1\, \P0[46]_net_1\, 
        \un3_ae[46]\, \un3_ae_2[46]\, \P0_75\, \P0_50[45]\, 
        \PDLCFG_DT_m_5[0]_net_1\, \P0_m[45]_net_1\, 
        \P0[45]_net_1\, \un3_ae[45]\, un3_ae_45_0, \P0_74\, 
        \P0_50[44]\, \PDLCFG_DT_m_4[0]_net_1\, \P0_m[44]_net_1\, 
        \P0[44]_net_1\, \un3_ae[44]\, \un3_ae_1[44]\, \P0_73\, 
        \P0_50[43]\, \P0_m_i[43]\, \PDLCFG_DT_m_3[0]_net_1\, 
        \P0[43]_net_1\, \un3_ae[43]\, \un3_ae_2[43]\, \P0_72\, 
        \P0_50[42]\, \P0_m_i[42]\, \PDLCFG_DT_m_2[0]_net_1\, 
        \P0[42]_net_1\, \un3_ae[42]\, \un3_ae_1[42]\, \P0_71\, 
        \P0_50[41]\, \P0_m_i[41]\, \PDLCFG_DT_m_1[0]_net_1\, 
        \P0[41]_net_1\, \un3_ae[41]\, \un3_ae_1[33]\, \P0_70\, 
        \P0_50[40]\, \P0_m_i[40]\, \PDLCFG_DT_m_0[0]_net_1\, 
        \P0[40]_net_1\, \un3_ae[40]\, \un3_ae_1[40]\, 
        \CNT[3]_net_1\, \CNT[5]_net_1\, \P0_69\, \P0_50[39]\, 
        \P0_m_i[39]\, \PDLCFG_DT_m_i[0]\, \un3_ae[39]\, 
        \P0[39]_net_1\, \un3_ae_1[39]\, \un3_ae_1_i[47]\, 
        \un3_ae_2[47]\, \P0_68\, \P0_50[38]\, \P0_m_i[38]\, 
        \PDLCFG_DT_m_22_i[0]\, \un3_ae[38]\, \P0[38]_net_1\, 
        \un3_ae_1_i[46]\, \P0_67\, \P0_50[37]\, 
        \PDLCFG_DT_m_21_i[0]\, \P0_m[37]_net_1\, \un3_ae[37]\, 
        \P0[37]_net_1\, \un3_ae_1[45]\, \P0_66\, \P0_50[36]\, 
        \PDLCFG_DT_m_20_i[0]\, \P0_m[36]_net_1\, \un3_ae[36]\, 
        \P0[36]_net_1\, \P0_65\, \P0_50[35]\, \P0_m_i[35]\, 
        \PDLCFG_DT_m_19_i[0]\, \un3_ae[35]\, \P0[35]_net_1\, 
        \un3_ae_1_i[43]\, \P0_64\, \P0_50[34]\, \P0_m_i[34]\, 
        \PDLCFG_DT_m_18_i[0]\, \un3_ae[34]\, \P0[34]_net_1\, 
        \P0_63\, \P0_50[33]\, \P0_m_i[33]\, \PDLCFG_DT_m_17_i[0]\, 
        \un3_ae[33]\, \P0[33]_net_1\, \un3_ae_1[41]\, 
        \CNT[0]_net_1\, \P0_62\, \P0_50[32]\, \P0_m_i[32]\, 
        \PDLCFG_DT_m_16_i[0]\, \un3_ae[32]\, \P0[32]_net_1\, 
        \P0_61\, \P0_50[31]\, \P0_m_i[31]\, 
        \PDLCFG_DT_m_15[0]_net_1\, \P0[31]_net_1\, \un3_ae[31]\, 
        \un3_ae_2[31]\, \un3_ae_3[31]\, \P0_60\, \P0_50[30]\, 
        \P0_m_i[30]\, \PDLCFG_DT_m_14[0]_net_1\, \P0[30]_net_1\, 
        \un3_ae[30]\, \un3_ae_1[30]\, \P0_59\, \P0_50[29]\, 
        \PDLCFG_DT_m_13[0]_net_1\, \P0_m[29]_net_1\, 
        \P0[29]_net_1\, \un3_ae[29]\, un3_ae_21_0, \P0_58\, 
        \P0_50[28]\, \P0_m_i[28]\, \PDLCFG_DT_m_12[0]_net_1\, 
        \P0[28]_net_1\, \un3_ae[28]\, \P0_57\, \P0_50[27]\, 
        \P0_m_i[27]\, \PDLCFG_DT_m_11[0]_net_1\, \P0[27]_net_1\, 
        \un3_ae[27]\, \un3_ae_1[27]\, \P0_56\, \P0_50[26]\, 
        \P0_m_i[26]\, \PDLCFG_DT_m_10[0]_net_1\, \P0[26]_net_1\, 
        \un3_ae[26]\, \un3_ae_1[26]\, \P0_55\, \P0_50[25]\, 
        \P0_m_i[25]\, \PDLCFG_DT_m_9[0]_net_1\, \P0[25]_net_1\, 
        \un3_ae[25]\, \un3_ae_1[25]\, \P0_54\, \P0_50[24]\, 
        \P0_m_i[24]\, \PDLCFG_DT_m_8[0]_net_1\, \P0[24]_net_1\, 
        \un3_ae[24]\, \un3_ae_1[24]\, \P0_53\, \P0_50[23]\, 
        \P0_m_i[23]\, \PDLCFG_DT_m_37_i[0]\, \un3_ae[23]\, 
        \P0[23]_net_1\, \un3_ae_1[23]\, \un3_ae_1_i[31]\, \P0_52\, 
        \P0_50[22]\, \P0_m[22]_net_1\, \PDLCFG_DT_m_36[0]_net_1\, 
        \un3_ae[22]\, \P0[22]_net_1\, \un3_ae_1[22]\, \P0_51\, 
        \P0_50[21]\, \PDLCFG_DT_m_35_i[0]\, \P0_m[21]_net_1\, 
        \un3_ae[21]\, \P0[21]_net_1\, \P0_50\, \P0_50[20]\, 
        \P0_m[20]_net_1\, \PDLCFG_DT_m_34[0]_net_1\, \un3_ae[20]\, 
        \P0[20]_net_1\, \P0_49\, \P0_50[19]\, \P0_m_i[19]\, 
        \PDLCFG_DT_m_33_i[0]\, \un3_ae[19]\, \P0[19]_net_1\, 
        \P0_48\, \P0_50[18]\, \PDLCFG_DT_m_32_i[0]\, \P0_m_i[18]\, 
        \P0[18]_net_1\, \un3_ae[18]\, \P0_47\, \P0_50[17]\, 
        \P0_m_i[17]\, \PDLCFG_DT_m_31_i[0]\, \un3_ae[17]\, 
        \P0[17]_net_1\, \P0_46\, \P0_50[16]\, 
        \PDLCFG_DT_m_30_i[0]\, \P0_m_i[16]\, \P0[16]_net_1\, 
        \un3_ae[16]\, \P0_45\, \P0_50[15]\, \P0_m[15]_net_1\, 
        \PDLCFG_DT_m_29[0]_net_1\, \un3_ae[15]\, \P0[15]_net_1\, 
        \un3_ae_2[7]\, \un3_ae_2[15]\, \P0_44\, \P0_50[14]\, 
        \P0_m[14]_net_1\, \PDLCFG_DT_m_28[0]_net_1\, \un3_ae[14]\, 
        \P0[14]_net_1\, \un3_ae_1[14]\, \P0_43\, \P0_50[13]\, 
        \PDLCFG_DT_m_27_i[0]\, \P0_m_i[13]\, \P0[13]_net_1\, 
        \un3_ae[13]\, \un3_ae_1[15]\, \P0_42\, \P0_50[12]\, 
        \PDLCFG_DT_m_26_i[0]\, \P0_m_i[12]\, \P0[12]_net_1\, 
        \un3_ae[12]\, \P0_41\, \P0_50[11]\, \P0_m_i[11]\, 
        \PDLCFG_DT_m_25[0]_net_1\, \REG_m_i[129]\, \P0[11]_net_1\, 
        \un3_ae[11]\, \un3_ae_1[11]\, \P0_40\, \P0_50[10]\, 
        \PDLCFG_DT_m_24_i[0]\, \P0_m_i[10]\, \P0[10]_net_1\, 
        \un3_ae[10]\, \P0_39\, \P0_50[9]\, \P0_m_i[9]\, 
        \PDLCFG_DT_m_23[0]_net_1\, \P0[9]_net_1\, \un3_ae[9]\, 
        \un3_ae_1[9]\, \P0_38\, \P0_50[8]\, \PDLCFG_DT_m_46_i[0]\, 
        \P0_m[8]_net_1\, \un3_ae[8]\, \P0[8]_net_1\, \P0_37\, 
        \P0_50[7]\, \P0_m[7]_net_1\, \PDLCFG_DT_m_45[0]_net_1\, 
        \un3_ae[7]\, \P0[7]_net_1\, \un3_ae_1[7]\, \P0_36\, 
        \P0_50[6]\, \P0_m[6]_net_1\, \PDLCFG_DT_m_44[0]_net_1\, 
        \un3_ae[6]\, \P0[6]_net_1\, \un3_ae_1[6]\, \P0_35\, 
        \P0_50[5]\, \PDLCFG_DT_m_43[0]_net_1\, \P0_m[5]_net_1\, 
        \P0[5]_net_1\, \un3_ae[5]\, \un3_ae_1[5]\, \P0_34\, 
        \P0_50[4]\, \PDLCFG_DT_m_42_i[0]\, \P0_m[4]_net_1\, 
        \un3_ae[4]\, \P0[4]_net_1\, \un3_ae_1[2]\, \P0_33\, 
        \P0_50[3]\, \un1_sstate_2\, \PDLCFG_DT_m_41_i[0]\, 
        \P0_m[3]_net_1\, \un3_ae[3]\, \P0[3]_net_1\, \P0_32\, 
        \P0_50[2]\, \PDLCFG_DT_m_40[0]_net_1\, \P0_m[2]_net_1\, 
        \P0[2]_net_1\, \un3_ae[2]\, \P0_31\, \P0_50[1]\, 
        \PDLCFG_DT_m_39_i[0]\, \P0_m[1]_net_1\, \un3_ae[1]\, 
        \P0[1]_net_1\, \P0_30\, \P0_50[0]\, \PDLCFG_DT_m_38_i[0]\, 
        \P0_m_i[0]\, \P0[0]_net_1\, \un3_ae[0]\, \VALID_29\, 
        \REG[145]\, \PDLCFG_RAD_28\, \PDLCFG_RAD_6[5]_net_1\, 
        \un1_sstate_25\, N_506, \PDLCFG_RAD_1_sqmuxa\, 
        \PDLCFG_RAD_27\, \PDLCFG_RAD_6[4]_net_1\, N_505, 
        \sstate[6]_net_1\, \PDLCFG_RAD_26\, 
        \PDLCFG_RAD_6[3]_net_1\, N_504, \PDLCFG_RAD_25\, 
        \PDLCFG_RAD_6[2]_net_1\, N_503, \PDLCFG_RAD_24\, 
        \PDLCFG_RAD_6[1]_net_1\, N_502, \PDLCFG_RAD_23\, 
        \PDLCFG_RAD_6[0]_net_1\, \un1_cnt\, N_501, \PDL_RACK_22\, 
        \un1_sstate_15\, \un1_sstate_16\, \un1_sstate_3_0\, 
        \PDL_RACK_1_sqmuxa\, \sstate[4]_net_1\, \PDL_RDATA_21\, 
        \PDL_RDATA_20\, \PDL_RDATA_19\, \PDL_RDATA_18\, 
        \PDL_RDATA_17\, \PDL_RDATA_16\, \PDL_RDATA_15\, 
        \PDL_RDATA_14\, \P_13\, \P_4[7]_net_1\, \P_12\, 
        \P_4[6]_net_1\, \P_11\, \P_4[5]_net_1\, \P_10\, 
        \P_4[4]_net_1\, \sstate[9]_net_1\, \P_9\, \P_4[3]_net_1\, 
        \P_8\, \P_4[2]_net_1\, \P_7\, \P_4[1]_net_1\, \MODE_2\, 
        \BITCNT_5[2]\, N_389, I_14_1, \sstate_0_sqmuxa\, 
        \BITCNT_5[1]\, I_13_5, \BITCNT_5[0]\, 
        \DWACT_ADD_CI_0_partial_sum[0]\, 
        \sstate_19_1_1_iv_0_i[6]\, \sstate_2_sqmuxa\, 
        \un5_bitcnt\, \sstate_19[0]\, \sstate_19[3]\, 
        \BITCNT[0]_net_1\, \BITCNT[2]_net_1\, \un3_pulse\, 
        \un1_sstate_21\, \sstate_19_1[10]\, \un1_cnt_0\, 
        \sstate_19[5]\, \SCLK_PDL_c\, PDLCFG_nRD_net_1, 
        \SI_PDL_c\, PDL_RACK_net_1, \PDLCFG_RAD[0]_net_1\, 
        \PDLCFG_RAD[1]_net_1\, \PDLCFG_RAD[2]_net_1\, 
        \PDLCFG_RAD[3]_net_1\, \PDLCFG_RAD[4]_net_1\, 
        \PDLCFG_RAD[5]_net_1\, \PDL_RDATA[0]_net_1\, 
        \PDL_RDATA[1]_net_1\, \PDL_RDATA[2]_net_1\, 
        \PDL_RDATA[3]_net_1\, \PDL_RDATA[4]_net_1\, 
        \PDL_RDATA[5]_net_1\, \PDL_RDATA[6]_net_1\, 
        \PDL_RDATA[7]_net_1\, \P_PDL_c[1]\, \P_PDL_c[2]\, 
        \P_PDL_c[3]\, \P_PDL_c[4]\, \P_PDL_c[5]\, \P_PDL_c[6]\, 
        \P_PDL_c[7]\, \sstate[5]_net_1\, 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, \CNT_2[1]\, \CNT_2[2]\, 
        \CNT_2[3]\, \CNT_2[4]\, \CNT_2[5]\, \GND\, \VCC\
         : std_logic;

begin 

    P_PDL_c(7) <= \P_PDL_c[7]\;
    P_PDL_c(6) <= \P_PDL_c[6]\;
    P_PDL_c(5) <= \P_PDL_c[5]\;
    P_PDL_c(4) <= \P_PDL_c[4]\;
    P_PDL_c(3) <= \P_PDL_c[3]\;
    P_PDL_c(2) <= \P_PDL_c[2]\;
    P_PDL_c(1) <= \P_PDL_c[1]\;
    PDL_RDATA(7) <= \PDL_RDATA[7]_net_1\;
    PDL_RDATA(6) <= \PDL_RDATA[6]_net_1\;
    PDL_RDATA(5) <= \PDL_RDATA[5]_net_1\;
    PDL_RDATA(4) <= \PDL_RDATA[4]_net_1\;
    PDL_RDATA(3) <= \PDL_RDATA[3]_net_1\;
    PDL_RDATA(2) <= \PDL_RDATA[2]_net_1\;
    PDL_RDATA(1) <= \PDL_RDATA[1]_net_1\;
    PDL_RDATA(0) <= \PDL_RDATA[0]_net_1\;
    PDLCFG_RAD(5) <= \PDLCFG_RAD[5]_net_1\;
    PDLCFG_RAD(4) <= \PDLCFG_RAD[4]_net_1\;
    PDLCFG_RAD(3) <= \PDLCFG_RAD[3]_net_1\;
    PDLCFG_RAD(2) <= \PDLCFG_RAD[2]_net_1\;
    PDLCFG_RAD(1) <= \PDLCFG_RAD[1]_net_1\;
    PDLCFG_RAD(0) <= \PDLCFG_RAD[0]_net_1\;
    P0(47) <= \P0[47]_net_1\;
    P0(46) <= \P0[46]_net_1\;
    P0(45) <= \P0[45]_net_1\;
    P0(44) <= \P0[44]_net_1\;
    P0(43) <= \P0[43]_net_1\;
    P0(42) <= \P0[42]_net_1\;
    P0(41) <= \P0[41]_net_1\;
    P0(40) <= \P0[40]_net_1\;
    P0(39) <= \P0[39]_net_1\;
    P0(38) <= \P0[38]_net_1\;
    P0(37) <= \P0[37]_net_1\;
    P0(36) <= \P0[36]_net_1\;
    P0(35) <= \P0[35]_net_1\;
    P0(34) <= \P0[34]_net_1\;
    P0(33) <= \P0[33]_net_1\;
    P0(32) <= \P0[32]_net_1\;
    P0(31) <= \P0[31]_net_1\;
    P0(30) <= \P0[30]_net_1\;
    P0(29) <= \P0[29]_net_1\;
    P0(28) <= \P0[28]_net_1\;
    P0(27) <= \P0[27]_net_1\;
    P0(26) <= \P0[26]_net_1\;
    P0(25) <= \P0[25]_net_1\;
    P0(24) <= \P0[24]_net_1\;
    P0(23) <= \P0[23]_net_1\;
    P0(22) <= \P0[22]_net_1\;
    P0(21) <= \P0[21]_net_1\;
    P0(20) <= \P0[20]_net_1\;
    P0(19) <= \P0[19]_net_1\;
    P0(18) <= \P0[18]_net_1\;
    P0(17) <= \P0[17]_net_1\;
    P0(16) <= \P0[16]_net_1\;
    P0(15) <= \P0[15]_net_1\;
    P0(14) <= \P0[14]_net_1\;
    P0(13) <= \P0[13]_net_1\;
    P0(12) <= \P0[12]_net_1\;
    P0(11) <= \P0[11]_net_1\;
    P0(10) <= \P0[10]_net_1\;
    P0(9) <= \P0[9]_net_1\;
    P0(8) <= \P0[8]_net_1\;
    P0(7) <= \P0[7]_net_1\;
    P0(6) <= \P0[6]_net_1\;
    P0(5) <= \P0[5]_net_1\;
    P0(4) <= \P0[4]_net_1\;
    P0(3) <= \P0[3]_net_1\;
    P0(2) <= \P0[2]_net_1\;
    P0(1) <= \P0[1]_net_1\;
    P0(0) <= \P0[0]_net_1\;
    AE_PDL_c(47) <= \AE_PDL_c[47]\;
    AE_PDL_c(46) <= \AE_PDL_c[46]\;
    AE_PDL_c(45) <= \AE_PDL_c[45]\;
    AE_PDL_c(44) <= \AE_PDL_c[44]\;
    AE_PDL_c(43) <= \AE_PDL_c[43]\;
    AE_PDL_c(42) <= \AE_PDL_c[42]\;
    AE_PDL_c(41) <= \AE_PDL_c[41]\;
    AE_PDL_c(40) <= \AE_PDL_c[40]\;
    AE_PDL_c(39) <= \AE_PDL_c[39]\;
    AE_PDL_c(38) <= \AE_PDL_c[38]\;
    AE_PDL_c(37) <= \AE_PDL_c[37]\;
    AE_PDL_c(36) <= \AE_PDL_c[36]\;
    AE_PDL_c(35) <= \AE_PDL_c[35]\;
    AE_PDL_c(34) <= \AE_PDL_c[34]\;
    AE_PDL_c(33) <= \AE_PDL_c[33]\;
    AE_PDL_c(32) <= \AE_PDL_c[32]\;
    AE_PDL_c(31) <= \AE_PDL_c[31]\;
    AE_PDL_c(30) <= \AE_PDL_c[30]\;
    AE_PDL_c(29) <= \AE_PDL_c[29]\;
    AE_PDL_c(28) <= \AE_PDL_c[28]\;
    AE_PDL_c(27) <= \AE_PDL_c[27]\;
    AE_PDL_c(26) <= \AE_PDL_c[26]\;
    AE_PDL_c(25) <= \AE_PDL_c[25]\;
    AE_PDL_c(24) <= \AE_PDL_c[24]\;
    AE_PDL_c(23) <= \AE_PDL_c[23]\;
    AE_PDL_c(22) <= \AE_PDL_c[22]\;
    AE_PDL_c(21) <= \AE_PDL_c[21]\;
    AE_PDL_c(20) <= \AE_PDL_c[20]\;
    AE_PDL_c(19) <= \AE_PDL_c[19]\;
    AE_PDL_c(18) <= \AE_PDL_c[18]\;
    AE_PDL_c(17) <= \AE_PDL_c[17]\;
    AE_PDL_c(16) <= \AE_PDL_c[16]\;
    AE_PDL_c(15) <= \AE_PDL_c[15]\;
    AE_PDL_c(14) <= \AE_PDL_c[14]\;
    AE_PDL_c(13) <= \AE_PDL_c[13]\;
    AE_PDL_c(12) <= \AE_PDL_c[12]\;
    AE_PDL_c(11) <= \AE_PDL_c[11]\;
    AE_PDL_c(10) <= \AE_PDL_c[10]\;
    AE_PDL_c(9) <= \AE_PDL_c[9]\;
    AE_PDL_c(8) <= \AE_PDL_c[8]\;
    AE_PDL_c(7) <= \AE_PDL_c[7]\;
    AE_PDL_c(6) <= \AE_PDL_c[6]\;
    AE_PDL_c(5) <= \AE_PDL_c[5]\;
    AE_PDL_c(4) <= \AE_PDL_c[4]\;
    AE_PDL_c(3) <= \AE_PDL_c[3]\;
    AE_PDL_c(2) <= \AE_PDL_c[2]\;
    AE_PDL_c(1) <= \AE_PDL_c[1]\;
    AE_PDL_c(0) <= \AE_PDL_c[0]\;
    REG_24 <= \REG[145]\;
    REG_16 <= \REG[137]\;
    REG_17 <= \REG[138]\;
    REG_18 <= \REG[139]\;
    REG_19 <= \REG[140]\;
    REG_20 <= \REG[141]\;
    REG_21 <= \REG[142]\;
    REG_22 <= \REG[143]\;
    REG_23 <= \REG[144]\;
    PDL_RACK <= PDL_RACK_net_1;
    SI_PDL_c <= \SI_PDL_c\;
    PDLCFG_nRD <= PDLCFG_nRD_net_1;
    SCLK_PDL_c <= \SCLK_PDL_c\;
    MD_PDL_c_0 <= \MD_PDL_c_0\;

    \P0_50_iv[30]\ : NAND3FTT
      port map(A => \P0_m_i[30]\, B => \PDLCFG_DT_m_14[0]_net_1\, 
        C => \REG_m_i_1[129]\, Y => \P0_50[30]\);
    
    \CNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, CLR => 
        \un1_load_res_4\, Q => \CNT[0]_net_1\);
    
    AE_0_sqmuxa_90 : AO21
      port map(A => \un69_ae_1[23]\, B => un69_ae_30_0, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_90\);
    
    un4_so_39_0_i : INV
      port map(A => N_490_i_i, Y => N_490_i);
    
    \PDLCFG_RAD_6[3]\ : MUX2H
      port map(A => \CNT[3]_net_1\, B => PDL_RADDR(3), S => 
        \sstate[6]_net_1\, Y => N_504);
    
    \BITCNT_5_r[0]\ : OA21
      port map(A => N_389, B => \DWACT_ADD_CI_0_partial_sum[0]\, 
        C => \sstate_0_sqmuxa\, Y => \BITCNT_5[0]\);
    
    un69_ae_14_1 : NOR2FT
      port map(A => REG_0(125), B => REG_1, Y => \un69_ae_1[14]\);
    
    \REG_i_m[182]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_61, Y => 
        \REG_i_m[182]_net_1\);
    
    \REG_i_m[166]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_45, Y => 
        \REG_i_m[166]_net_1\);
    
    \AE[36]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_116\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[36]\);
    
    \REG_i_m[155]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_34, Y => 
        \REG_i_m[155]_net_1\);
    
    un69_ae_46_1 : OR2
      port map(A => REG_1, B => REG_0(126), Y => 
        \un69_ae_1_i[46]\);
    
    AE_0_sqmuxa_16 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[4]\, Y => 
        \AE_0_sqmuxa_16\);
    
    un4_so_24_0 : MUX2H
      port map(A => SP_PDL_in(1), B => SP_PDL_in(33), S => REG_6, 
        Y => N_475);
    
    \P0_m[41]\ : AND2FT
      port map(A => \AE_0_sqmuxa_164\, B => \P0[41]_net_1\, Y => 
        \P0_m_i[41]\);
    
    \sstate_7[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_7[9]_net_1\);
    
    \REG_i_m[176]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_55, Y => 
        \REG_i_m[176]_net_1\);
    
    \P0[39]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_69\, CLR => 
        \un1_load_res_7\, Q => \P0[39]_net_1\);
    
    \AE_7_r[8]\ : AND3FFT
      port map(A => \AE_i_m[8]_net_1\, B => \REG_i_m[161]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[8]\);
    
    \REG_i_m[180]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_59, Y => 
        \REG_i_m[180]_net_1\);
    
    MODE_2 : OR2
      port map(A => REG_0_d0, B => \sstate[12]_net_1\, Y => 
        \MODE_2\);
    
    ISCK_128 : MUX2H
      port map(A => \SCLK_PDL_c\, B => \sstate[3]_net_1\, S => 
        \un1_sstate_13\, Y => \ISCK_128\);
    
    \AE_7_r[24]\ : AND3FFT
      port map(A => \AE_i_m[24]_net_1\, B => \REG_i_m[177]_net_1\, 
        C => N_6864_1, Y => \AE_7[24]\);
    
    \AE_7_r[2]\ : AND3FFT
      port map(A => \AE_i_m[2]_net_1\, B => \REG_i_m[155]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[2]\);
    
    \AE_i_m[41]\ : AOI21
      port map(A => \AE_0_sqmuxa_164\, B => \AE_0_sqmuxa_166\, C
         => \AE_PDL_c[41]\, Y => \AE_i_m[41]_net_1\);
    
    AE_0_sqmuxa_26 : AO21
      port map(A => \un69_ae_1[6]\, B => \un69_ae_2[7]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_26\);
    
    un3_ae_47_3 : AND2
      port map(A => \CNT[3]_net_1\, B => \CNT[5]_net_1\, Y => 
        \un3_ae_3[47]\);
    
    un1_sstate_22 : OR2FT
      port map(A => \ISI_1_sqmuxa_1\, B => \sstate[12]_net_1\, Y
         => \un1_sstate_22\);
    
    \REG_i_m[189]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_68, Y => 
        \REG_i_m[189]_net_1\);
    
    AE_0_sqmuxa_72 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[18]\, Y => 
        \AE_0_sqmuxa_72\);
    
    un3_ae_32 : AND2
      port map(A => \un3_ae_1[39]\, B => \un3_ae_1[40]\, Y => 
        \un3_ae[32]\);
    
    un1_cnt_0 : OR2FT
      port map(A => \CNT[5]_net_1\, B => \CNT[0]_net_1\, Y => 
        \un1_cnt_0\);
    
    un3_ae_26 : NAND2
      port map(A => \un3_ae_1[26]\, B => \un3_ae_2[31]\, Y => 
        \un3_ae[26]\);
    
    un1_load_res_0 : OR2FT
      port map(A => LOAD_RES, B => HWRES_c_0_3, Y => 
        \un1_load_res_0\);
    
    un3_ae_46 : NAND2
      port map(A => \un3_ae_2[46]\, B => \un3_ae_3[47]\, Y => 
        \un3_ae[46]\);
    
    un69_ae_13_0 : NOR2FT
      port map(A => \un69_ae_2[15]\, B => \un69_ae_1[45]\, Y => 
        \un69_ae_13_0\);
    
    \PDLCFG_RAD[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDLCFG_RAD_27\, CLR => 
        \un1_load_res_9\, Q => \PDLCFG_RAD[4]_net_1\);
    
    un1_sstate_2_3 : OR2
      port map(A => \sstate_0[9]_net_1\, B => \sstate_0[6]_net_1\, 
        Y => \un1_sstate_2_3\);
    
    \sstate_19_1[11]\ : OR2
      port map(A => \sstate[8]_net_1\, B => \sstate[12]_net_1\, Y
         => \sstate_19_1[11]_net_1\);
    
    un4_so_42_0 : MUX2H
      port map(A => SP_PDL_in(43), B => SP_PDL_in(47), S => REG_3, 
        Y => N_493);
    
    \AE_i_m[38]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_152\, B => \AE_0_sqmuxa_154\, C
         => \AE_PDL_c[38]\, Y => \AE_i_m[38]_net_1\);
    
    \P_4[5]\ : MUX2H
      port map(A => REG_13, B => PDLCFG_DT(5), S => 
        \sstate_8[9]_net_1\, Y => \P_4[5]_net_1\);
    
    P_11 : MUX2H
      port map(A => \P_PDL_c[5]\, B => \P_4[5]_net_1\, S => 
        \un1_sstate_2\, Y => \P_11\);
    
    \P0_50_iv[40]\ : NAND3FTT
      port map(A => \P0_m_i[40]\, B => \PDLCFG_DT_m_0[0]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[40]\);
    
    un3_ae_19 : NOR2FT
      port map(A => \un3_ae_1[27]\, B => \un3_ae_1[23]\, Y => 
        \un3_ae[19]\);
    
    \AE_7_r[18]\ : AND3FFT
      port map(A => \AE_i_m[18]_net_1\, B => \REG_i_m[171]_net_1\, 
        C => N_6864_2, Y => \AE_7[18]\);
    
    un3_ae_30 : OR3FTT
      port map(A => \un3_ae_2[31]\, B => \un3_ae_1[30]\, C => 
        \un3_ae_2[47]\, Y => \un3_ae[30]\);
    
    \P[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \P_7\, CLR => 
        \un1_load_res_10\, Q => \P_PDL_c[1]\);
    
    \PDLCFG_DT_m_11[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[27]\, Y => \PDLCFG_DT_m_11[0]_net_1\);
    
    \P0_m[38]\ : AND2
      port map(A => \AE_0_sqmuxa_152\, B => \P0[38]_net_1\, Y => 
        \P0_m_i[38]\);
    
    AE_0_sqmuxa_144 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[36]\, Y => 
        \AE_0_sqmuxa_144\);
    
    \AE[37]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_117\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[37]\);
    
    \REG_i_m[200]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_79, Y => 
        \REG_i_m[200]_net_1\);
    
    AE_0_sqmuxa_12 : NOR2FT
      port map(A => \sstate_0[9]_net_1\, B => \un3_ae[3]\, Y => 
        \AE_0_sqmuxa_12\);
    
    un4_so_28_0_i : INV
      port map(A => N_479_i_i, Y => N_479_i);
    
    \REG_i_m[154]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_33, Y => 
        \REG_i_m[154]_net_1\);
    
    AE_0_sqmuxa_182 : AO21
      port map(A => \un69_ae_3[47]\, B => un69_ae_37_0, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_182\);
    
    \P0_50_iv[37]\ : NAND3FTT
      port map(A => \PDLCFG_DT_m_21_i[0]\, B => \P0_m[37]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[37]\);
    
    un4_so_40_0 : MUX2H
      port map(A => SP_PDL_in(7), B => SP_PDL_in(39), S => REG_6, 
        Y => N_491);
    
    \PDLCFG_DT_m_26[0]\ : AND3
      port map(A => PDLCFG_DT_0_0(0), B => \un3_ae[12]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_26_i[0]\);
    
    \PDLCFG_DT_m_46[0]\ : AND3
      port map(A => PDLCFG_DT_0_0(0), B => \un3_ae[8]\, C => 
        \sstate_8[9]_net_1\, Y => \PDLCFG_DT_m_46_i[0]\);
    
    \REG_i_m[153]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_32, Y => 
        \REG_i_m[153]_net_1\);
    
    \P0[41]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_71\, CLR => 
        \un1_load_res_7\, Q => \P0[41]_net_1\);
    
    AE_0_sqmuxa_36 : NAND2
      port map(A => \sstate_7[9]_net_1\, B => \un3_ae[9]\, Y => 
        \AE_0_sqmuxa_36\);
    
    \sstate_6[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_6[9]_net_1\);
    
    AE_1_sqmuxa_1 : OR2FT
      port map(A => \sstate_0[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        \AE_1_sqmuxa_1\);
    
    un3_ae_23 : NOR2FT
      port map(A => \un3_ae_3[31]\, B => \un3_ae_1[23]\, Y => 
        \un3_ae[23]\);
    
    \AE[45]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_125\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[45]\);
    
    \sstate_3[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_3[9]_net_1\);
    
    MODE_1 : DFFB
      port map(CLK => CLK_c_c, D => \MODE_0\, CLR => 
        un1_hwres_1_i, SET => \un1_reg_1_i\, Q => MD_PDL_c_1);
    
    AE_0_sqmuxa_0_0 : NAND2
      port map(A => \sstate_1[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        AE_0_sqmuxa_i_0);
    
    un3_ae_43 : NAND2
      port map(A => \un3_ae_2[43]\, B => \un3_ae_3[47]\, Y => 
        \un3_ae[43]\);
    
    \PDLCFG_DT_m_7[0]\ : OR3FFT
      port map(A => \sstate_2[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[47]\, Y => \PDLCFG_DT_m_7[0]_net_1\);
    
    un1_BITCNT_I_14 : XOR2
      port map(A => \BITCNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, Y => I_14_1);
    
    un3_ae_2 : OR2
      port map(A => \un3_ae_1[2]\, B => \un3_ae_1_i[43]\, Y => 
        \un3_ae[2]\);
    
    \AE[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_82\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[2]\);
    
    \REG_i_m[187]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_66, Y => 
        \REG_i_m[187]_net_1\);
    
    \PDLCFG_DT_m_29[0]\ : NAND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[15]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_29[0]_net_1\);
    
    AE_0_sqmuxa_22 : OAI21FTF
      port map(A => \un69_ae_1[5]\, B => \un69_ae_1[45]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_22\);
    
    \P0[40]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_70\, CLR => 
        \un1_load_res_7\, Q => \P0[40]_net_1\);
    
    un3_ae_4 : NOR2
      port map(A => \un3_ae_1[2]\, B => \un3_ae_1[45]\, Y => 
        \un3_ae[4]\);
    
    un69_ae_23_2 : NOR2
      port map(A => \un69_ae_1_i[31]\, B => \un69_ae_2[47]\, Y
         => \un69_ae_3[31]\);
    
    P_7 : MUX2H
      port map(A => \P_PDL_c[1]\, B => \P_4[1]_net_1\, S => 
        \un1_sstate_2\, Y => \P_7\);
    
    un3_ae_36_1 : NOR2
      port map(A => \un3_ae_1[45]\, B => \un3_ae_1_i[46]\, Y => 
        \un3_ae_1[44]\);
    
    \PDL_RDATA[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_18\, CLR => 
        \un1_load_res_9\, Q => \PDL_RDATA[4]_net_1\);
    
    \AE_7_r[37]\ : AND3FFT
      port map(A => \AE_i_m[37]_net_1\, B => \REG_i_m[190]_net_1\, 
        C => N_6864_0, Y => \AE_7[37]\);
    
    \PDLCFG_DT_m_15[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[31]\, Y => \PDLCFG_DT_m_15[0]_net_1\);
    
    un1_sstate_14_0 : OR3
      port map(A => \un1_sstate_5\, B => \sstate_0[9]_net_1\, C
         => \sstate[11]_net_1\, Y => \un1_sstate_14_0\);
    
    \PDLCFG_RAD_6[1]\ : MUX2H
      port map(A => \CNT[1]_net_1\, B => PDL_RADDR(1), S => 
        \sstate[6]_net_1\, Y => N_502);
    
    AE_0_sqmuxa_0 : NOR2FT
      port map(A => \sstate_0[9]_net_1\, B => \un3_ae[0]\, Y => 
        \AE_0_sqmuxa_0\);
    
    P0_36 : MUX2H
      port map(A => \P0[6]_net_1\, B => \P0_50[6]\, S => 
        \un1_sstate_2_3\, Y => \P0_36\);
    
    AE_1_sqmuxa_2 : OR2FT
      port map(A => \sstate_0[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        \AE_1_sqmuxa_2\);
    
    \SBYTE[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_135\, CLR => 
        \un1_load_res_11\, Q => \REG[143]\);
    
    AE_93 : MUX2H
      port map(A => \AE_PDL_c[13]\, B => \AE_7[13]\, S => 
        \un1_sstate_14_2\, Y => \AE_93\);
    
    P0_39 : MUX2H
      port map(A => \P0[9]_net_1\, B => \P0_50[9]\, S => 
        \un1_sstate_2_3\, Y => \P0_39\);
    
    \AE_7_r[35]\ : AND3FFT
      port map(A => \AE_i_m[35]_net_1\, B => \REG_i_m[188]_net_1\, 
        C => N_6864_1, Y => \AE_7[35]\);
    
    \P0_50_iv[24]\ : NAND3FTT
      port map(A => \P0_m_i[24]\, B => \PDLCFG_DT_m_8[0]_net_1\, 
        C => \REG_m_i_1[129]\, Y => \P0_50[24]\);
    
    AE_0_sqmuxa_178 : AO21
      port map(A => \un69_ae_1[44]\, B => \un69_ae_3[47]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_178\);
    
    un3_ae_33_1 : NOR2
      port map(A => \un3_ae_1[41]\, B => \un3_ae_1_i[47]\, Y => 
        \un3_ae_1[33]\);
    
    un4_so_3_0 : MUX2H
      port map(A => SP_PDL_in(8), B => SP_PDL_in(40), S => 
        REG_0(127), Y => N_454);
    
    \sstate[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_19[3]\, CLR => 
        \un1_load_res\, Q => \sstate[3]_net_1\);
    
    \P0_m[9]\ : AND2FT
      port map(A => \AE_0_sqmuxa_36\, B => \P0[9]_net_1\, Y => 
        \P0_m_i[9]\);
    
    un69_ae_45_0 : NOR2
      port map(A => \un69_ae_1[45]\, B => \un69_ae_1_i[47]\, Y
         => un69_ae_37_0);
    
    un69_ae_17_1 : NOR2
      port map(A => \un69_ae_1_i[31]\, B => \un69_ae_1[41]\, Y
         => \un69_ae_1[25]\);
    
    un4_so_44_0 : MUX2H
      port map(A => N_489, B => N_494, S => REG_5, Y => N_495_i_i);
    
    \P0[32]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_62\, CLR => 
        \un1_load_res_7\, Q => \P0[32]_net_1\);
    
    \AE[33]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_113\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[33]\);
    
    AE_86 : MUX2H
      port map(A => \AE_PDL_c[6]\, B => \AE_7[6]\, S => 
        \un1_sstate_14\, Y => \AE_86\);
    
    P0_76 : MUX2H
      port map(A => \P0[46]_net_1\, B => \P0_50[46]\, S => 
        \un1_sstate_2_0\, Y => \P0_76\);
    
    AE_89 : MUX2H
      port map(A => \AE_PDL_c[9]\, B => \AE_7[9]\, S => 
        \un1_sstate_14\, Y => \AE_89\);
    
    un3_ae_24 : NAND2
      port map(A => \un3_ae_1[24]\, B => \un3_ae_2[31]\, Y => 
        \un3_ae[24]\);
    
    P0_45 : MUX2H
      port map(A => \P0[15]_net_1\, B => \P0_50[15]\, S => 
        \un1_sstate_2_2\, Y => \P0_45\);
    
    un3_ae_44 : NAND2
      port map(A => \un3_ae_1[44]\, B => \un3_ae_3[47]\, Y => 
        \un3_ae[44]\);
    
    un3_ae_31 : NAND2
      port map(A => \un3_ae_2[31]\, B => \un3_ae_3[31]\, Y => 
        \un3_ae[31]\);
    
    \PDLCFG_DT_m_31[0]\ : AND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[17]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_31_i[0]\);
    
    AE_0_sqmuxa_186 : AO21
      port map(A => \un69_ae_1[38]\, B => \un69_ae_3[47]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_186\);
    
    \PDLCFG_DT_m_0[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[40]\, Y => \PDLCFG_DT_m_0[0]_net_1\);
    
    AE_0_sqmuxa_8 : NAND2
      port map(A => \sstate_8[9]_net_1\, B => \un3_ae[2]\, Y => 
        \AE_0_sqmuxa_8\);
    
    P0_55 : MUX2H
      port map(A => \P0[25]_net_1\, B => \P0_50[25]\, S => 
        \un1_sstate_2_2\, Y => \P0_55\);
    
    \P0_50_iv[47]\ : NAND3FTT
      port map(A => \P0_m_i[47]\, B => \PDLCFG_DT_m_7[0]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[47]\);
    
    AE_0_sqmuxa_32 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[8]\, Y => 
        \AE_0_sqmuxa_32\);
    
    sstate_0_sqmuxa : OR2FT
      port map(A => \sstate_1[6]_net_1\, B => \un3_pulse\, Y => 
        \sstate_0_sqmuxa\);
    
    PDL_RDATA_14 : MUX2H
      port map(A => \PDL_RDATA[0]_net_1\, B => PDLCFG_DT(0), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_14\);
    
    P_13 : MUX2H
      port map(A => \P_PDL_c[7]\, B => \P_4[7]_net_1\, S => 
        \un1_sstate_2\, Y => \P_13\);
    
    P0_65 : MUX2H
      port map(A => \P0[35]_net_1\, B => \P0_50[35]\, S => 
        \un1_sstate_2_1\, Y => \P0_65\);
    
    un3_ae_35 : AND2
      port map(A => \un3_ae_1[39]\, B => \un3_ae_2[43]\, Y => 
        \un3_ae[35]\);
    
    \CNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_2[3]\, CLR => 
        \un1_load_res_4\, Q => \CNT[3]_net_1\);
    
    \PDLCFG_RAD_6[5]\ : MUX2H
      port map(A => \CNT[5]_net_1\, B => PDL_RADDR(5), S => 
        \sstate_2[6]_net_1\, Y => N_506);
    
    PDLCFG_RAD_28 : MUX2H
      port map(A => \PDLCFG_RAD_6[5]_net_1\, B => 
        \PDLCFG_RAD[5]_net_1\, S => \un1_sstate_25\, Y => 
        \PDLCFG_RAD_28\);
    
    AE_0_sqmuxa_158 : AOI21
      port map(A => \un69_ae_1[39]\, B => \un69_ae_4[47]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_158\);
    
    PDL_RDATA_21 : MUX2H
      port map(A => \PDL_RDATA[7]_net_1\, B => PDLCFG_DT(7), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_21\);
    
    un1_sstate_2_0 : OR2
      port map(A => \sstate_0[9]_net_1\, B => \sstate_0[6]_net_1\, 
        Y => \un1_sstate_2_0\);
    
    \P0_50_iv[21]\ : NAND3FTT
      port map(A => \PDLCFG_DT_m_35_i[0]\, B => \P0_m[21]_net_1\, 
        C => \REG_m_i_2[129]\, Y => \P0_50[21]\);
    
    SBYTE_133 : MUX2H
      port map(A => \SBYTE_5[4]_net_1\, B => \REG[141]\, S => 
        \un1_sstate_20\, Y => \SBYTE_133\);
    
    \P0[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_55\, CLR => 
        \un1_load_res_6\, Q => \P0[25]_net_1\);
    
    \PDLCFG_DT_m_35[0]\ : AND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[21]\, C => 
        \sstate_6[9]_net_1\, Y => \PDLCFG_DT_m_35_i[0]\);
    
    \P0[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_45\, CLR => 
        \un1_load_res_5\, Q => \P0[15]_net_1\);
    
    \PDLCFG_DT_m_18[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[34]\, C => 
        \sstate_5[9]_net_1\, Y => \PDLCFG_DT_m_18_i[0]\);
    
    un3_ae_1_1 : NOR2
      port map(A => \un3_ae_1[15]\, B => \un3_ae_1[41]\, Y => 
        \un3_ae_1[9]\);
    
    P0_40 : MUX2H
      port map(A => \P0[10]_net_1\, B => \P0_50[10]\, S => 
        \un1_sstate_2_3\, Y => \P0_40\);
    
    un3_ae_18 : NOR2FT
      port map(A => \un3_ae_1[26]\, B => \un3_ae_1[23]\, Y => 
        \un3_ae[18]\);
    
    CNT_2_I_21 : XOR2
      port map(A => \CNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP_0[0]\, Y => \CNT_2[1]\);
    
    P0_50 : MUX2H
      port map(A => \P0[20]_net_1\, B => \P0_50[20]\, S => 
        \un1_sstate_2_2\, Y => \P0_50\);
    
    \AE_i_m[34]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_136\, B => \AE_0_sqmuxa_138\, C
         => \AE_PDL_c[34]\, Y => \AE_i_m[34]_net_1\);
    
    \AE_7_r[21]\ : AND3FFT
      port map(A => \AE_i_m[21]_net_1\, B => \REG_i_m[174]_net_1\, 
        C => N_6864_2, Y => \AE_7[21]\);
    
    \PDLCFG_RAD[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDLCFG_RAD_24\, CLR => 
        \un1_load_res_9\, Q => \PDLCFG_RAD[1]_net_1\);
    
    \PDLCFG_DT_m_10[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[26]\, Y => \PDLCFG_DT_m_10[0]_net_1\);
    
    un3_ae_39_1 : NOR2FT
      port map(A => \CNT[5]_net_1\, B => \CNT[3]_net_1\, Y => 
        \un3_ae_1[39]\);
    
    \P0_m[2]\ : NAND2FT
      port map(A => \AE_0_sqmuxa_8\, B => \P0[2]_net_1\, Y => 
        \P0_m[2]_net_1\);
    
    \AE_i_m[23]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_92\, B => \AE_0_sqmuxa_94\, C
         => \AE_PDL_c[23]\, Y => \AE_i_m[23]_net_1\);
    
    \AE_7_r[14]\ : AND3FFT
      port map(A => \AE_i_m[14]_net_1\, B => \REG_i_m[167]_net_1\, 
        C => N_6864_2, Y => \AE_7[14]\);
    
    AE_0_sqmuxa_58 : AOI21
      port map(A => \un69_ae_1[14]\, B => \un69_ae_2[7]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_58\);
    
    un69_ae_36_1 : NOR2
      port map(A => \un69_ae_1[45]\, B => \un69_ae_1_i[46]\, Y
         => \un69_ae_1[44]\);
    
    P0_60 : MUX2H
      port map(A => \P0[30]_net_1\, B => \P0_50[30]\, S => 
        \un1_sstate_2_1\, Y => \P0_60\);
    
    AE_0_sqmuxa_48 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[12]\, Y => 
        \AE_0_sqmuxa_48\);
    
    \P0[44]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_74\, CLR => 
        \un1_load_res_8\, Q => \P0[44]_net_1\);
    
    PDL_RDATA_17 : MUX2H
      port map(A => \PDL_RDATA[3]_net_1\, B => PDLCFG_DT(3), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_17\);
    
    PDLCFG_RAD_24 : MUX2H
      port map(A => \PDLCFG_RAD_6[1]_net_1\, B => 
        \PDLCFG_RAD[1]_net_1\, S => \un1_sstate_25\, Y => 
        \PDLCFG_RAD_24\);
    
    un1_reg_1_i : INV
      port map(A => un1_reg_1_i_i, Y => \un1_reg_1_i\);
    
    AE_119 : MUX2H
      port map(A => \AE_PDL_c[39]\, B => \AE_7[39]\, S => 
        \un1_sstate_14_0\, Y => \AE_119\);
    
    \PDLCFG_DT_m_17[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[33]\, C => 
        \sstate_5[9]_net_1\, Y => \PDLCFG_DT_m_17_i[0]\);
    
    un69_ae_43_1 : OR2FT
      port map(A => REG_2, B => REG_0(124), Y => \un69_ae_1[43]\);
    
    \sstate[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_19_1[11]_net_1\, CLR
         => \un1_load_res_11\, Q => \sstate[11]_net_1\);
    
    \P0_m[45]\ : NAND2FT
      port map(A => \AE_0_sqmuxa_180\, B => \P0[45]_net_1\, Y => 
        \P0_m[45]_net_1\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    AE_0_sqmuxa_60 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[15]\, Y => 
        \AE_0_sqmuxa_60\);
    
    \PDLCFG_RAD_6_r[2]\ : AND2
      port map(A => N_503, B => \PDLCFG_RAD_1_sqmuxa\, Y => 
        \PDLCFG_RAD_6[2]_net_1\);
    
    un4_so_16_0_i : INV
      port map(A => N_467_i_i, Y => N_467_i);
    
    un1_sstate_13 : OR3
      port map(A => \un1_sstate_1\, B => \un1_sstate_13_0\, C => 
        \sstate[3]_net_1\, Y => \un1_sstate_13\);
    
    un1_load_res_7 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_3, Y => 
        \un1_load_res_7\);
    
    \PDLCFG_nRD\ : DFFS
      port map(CLK => CLK_c_c, D => \PDLCFG_nRD_79\, SET => 
        \un1_load_res_9\, Q => PDLCFG_nRD_net_1);
    
    un1_load_res_3 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_3, Y => 
        \un1_load_res_3\);
    
    \P0_50_iv[4]\ : NAND3FTT
      port map(A => \PDLCFG_DT_m_42_i[0]\, B => \P0_m[4]_net_1\, 
        C => \REG_m_i[129]\, Y => \P0_50[4]\);
    
    un4_so_21_0_i : INV
      port map(A => N_472_i_i, Y => N_472_i);
    
    un69_ae_31_2 : AND2
      port map(A => REG_4, B => REG_5, Y => \un69_ae_2[31]\);
    
    \AE[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_95\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[15]\);
    
    \PDLCFG_DT_m_38[0]\ : AND3
      port map(A => PDLCFG_DT(0), B => \un3_ae[0]\, C => 
        \sstate_8[9]_net_1\, Y => \PDLCFG_DT_m_38_i[0]\);
    
    \P0_m[14]\ : NAND2
      port map(A => \AE_0_sqmuxa_56\, B => \P0[14]_net_1\, Y => 
        \P0_m[14]_net_1\);
    
    un3_ae_45_1 : OR2FT
      port map(A => \CNT[2]_net_1\, B => \CNT[1]_net_1\, Y => 
        \un3_ae_1[45]\);
    
    \AE_i_m[43]\ : AOI21
      port map(A => \AE_0_sqmuxa_172\, B => \AE_0_sqmuxa_174\, C
         => \AE_PDL_c[43]\, Y => \AE_i_m[43]_net_1\);
    
    un69_ae_41_1 : OR2
      port map(A => REG_0(124), B => REG_2, Y => \un69_ae_1[41]\);
    
    \PDLCFG_DT_m_14[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[30]\, Y => \PDLCFG_DT_m_14[0]_net_1\);
    
    AE_0_sqmuxa_148 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[37]\, Y => 
        \AE_0_sqmuxa_148\);
    
    \AE[44]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_124\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[44]\);
    
    \PDL_RDATA[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_15\, CLR => 
        \un1_load_res_9\, Q => \PDL_RDATA[1]_net_1\);
    
    \P0_50_iv[28]\ : NAND3FTT
      port map(A => \P0_m_i[28]\, B => \PDLCFG_DT_m_12[0]_net_1\, 
        C => \REG_m_i_1[129]\, Y => \P0_50[28]\);
    
    \PDLCFG_DT_m_30[0]\ : AND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[16]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_30_i[0]\);
    
    \AE_i_m[29]\ : AOI21
      port map(A => \AE_0_sqmuxa_116\, B => \AE_0_sqmuxa_118\, C
         => \AE_PDL_c[29]\, Y => \AE_i_m[29]_net_1\);
    
    un1_load_res_1 : OR2FT
      port map(A => LOAD_RES, B => HWRES_c_0_3, Y => 
        \un1_load_res_1\);
    
    \PDLCFG_DT_m_9[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[25]\, Y => \PDLCFG_DT_m_9[0]_net_1\);
    
    AE_0_sqmuxa_110 : AO21
      port map(A => \un69_ae_1[27]\, B => \un69_ae_2[31]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_110\);
    
    \P0_m[24]\ : AND2FT
      port map(A => \AE_0_sqmuxa_96\, B => \P0[24]_net_1\, Y => 
        \P0_m_i[24]\);
    
    \AE_7_r[1]\ : AND3FFT
      port map(A => \AE_i_m[1]_net_1\, B => \REG_i_m[154]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[1]\);
    
    \P0_50_iv[14]\ : NAND3
      port map(A => \P0_m[14]_net_1\, B => 
        \PDLCFG_DT_m_28[0]_net_1\, C => \REG_m_i_2[129]\, Y => 
        \P0_50[14]\);
    
    \P0_50_iv[2]\ : NAND3
      port map(A => \PDLCFG_DT_m_40[0]_net_1\, B => 
        \P0_m[2]_net_1\, C => \REG_m_i[129]\, Y => \P0_50[2]\);
    
    P0_33 : MUX2H
      port map(A => \P0[3]_net_1\, B => \P0_50[3]\, S => 
        \un1_sstate_2\, Y => \P0_33\);
    
    un69_ae_39_1 : NOR2FT
      port map(A => REG_0(127), B => REG_0(125), Y => 
        \un69_ae_1[39]\);
    
    \P0[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_32\, CLR => 
        \un1_load_res_6\, Q => \P0[2]_net_1\);
    
    un1_sstate_21 : AND2
      port map(A => \ISI_1_sqmuxa_1\, B => \un1_sstate_1\, Y => 
        \un1_sstate_21\);
    
    \sstate[6]\ : DFFB
      port map(CLK => CLK_c_c, D => \sstate_19_1[6]\, CLR => 
        un2_load_res_i, SET => HWRES_c_23_0, Q => 
        \sstate[6]_net_1\);
    
    \PDLCFG_DT_m_37[0]\ : AND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[23]\, C => 
        \sstate_6[9]_net_1\, Y => \PDLCFG_DT_m_37_i[0]\);
    
    P0_47 : MUX2H
      port map(A => \P0[17]_net_1\, B => \P0_50[17]\, S => 
        \un1_sstate_2_2\, Y => \P0_47\);
    
    un4_so_15_0 : MUX2H
      port map(A => N_465, B => SP_PDL_in(26), S => REG_5, Y => 
        N_466);
    
    \AE_i_m[20]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_80\, B => \AE_0_sqmuxa_82\, C
         => \AE_PDL_c[20]\, Y => \AE_i_m[20]_net_1\);
    
    MODE_3 : DFFB
      port map(CLK => CLK_c_c, D => \MODE_0\, CLR => 
        un1_hwres_1_i, SET => \un1_reg_1_i\, Q => MD_PDL_c_3);
    
    \AE_i_m[5]\ : AOI21
      port map(A => \AE_0_sqmuxa_20\, B => \AE_0_sqmuxa_22\, C
         => \AE_PDL_c[5]\, Y => \AE_i_m[5]_net_1\);
    
    \P0_50_iv[23]\ : NAND3FFT
      port map(A => \P0_m_i[23]\, B => \PDLCFG_DT_m_37_i[0]\, C
         => \REG_m_i_2[129]\, Y => \P0_50[23]\);
    
    P0_57 : MUX2H
      port map(A => \P0[27]_net_1\, B => \P0_50[27]\, S => 
        \un1_sstate_2_1\, Y => \P0_57\);
    
    un1_BITCNT_I_9 : XOR2
      port map(A => \BITCNT[0]_net_1\, B => \un1_sstate_21\, Y
         => \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \sstate_2[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_2[9]_net_1\);
    
    P0_73 : MUX2H
      port map(A => \P0[43]_net_1\, B => \P0_50[43]\, S => 
        \un1_sstate_2_0\, Y => \P0_73\);
    
    AE_118 : MUX2H
      port map(A => \AE_PDL_c[38]\, B => \AE_7[38]\, S => 
        \un1_sstate_14_0\, Y => \AE_118\);
    
    un3_ae_40_1 : NOR2
      port map(A => \un3_ae_1[41]\, B => \un3_ae_1_i[46]\, Y => 
        \un3_ae_1[40]\);
    
    \PDLCFG_RAD_6[0]\ : MUX2H
      port map(A => \CNT[0]_net_1\, B => PDL_RADDR(0), S => 
        \sstate[6]_net_1\, Y => N_501);
    
    AE_0_sqmuxa_160 : NAND2
      port map(A => \sstate_5[9]_net_1\, B => \un3_ae[40]\, Y => 
        \AE_0_sqmuxa_160\);
    
    un4_so_44_0_i : INV
      port map(A => N_495_i_i, Y => N_495_i);
    
    un1_sstate_5 : OR2
      port map(A => \sstate[12]_net_1\, B => \sstate_1[6]_net_1\, 
        Y => \un1_sstate_5\);
    
    \SBYTE_5[1]\ : MUX2H
      port map(A => \REG[137]\, B => REG_9, S => 
        \sstate_2[6]_net_1\, Y => \SBYTE_5[1]_net_1\);
    
    \REG_i_m[195]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_74, Y => 
        \REG_i_m[195]_net_1\);
    
    \P[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \P_12\, CLR => 
        \un1_load_res_10\, Q => \P_PDL_c[6]\);
    
    P0_67 : MUX2H
      port map(A => \P0[37]_net_1\, B => \P0_50[37]\, S => 
        \un1_sstate_2_0\, Y => \P0_67\);
    
    AE_0_sqmuxa_86 : AOI21
      port map(A => \un69_ae_1[23]\, B => \un69_ae_1[29]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_86\);
    
    un1_hwres_1 : NOR2FT
      port map(A => HWRES_c_0, B => REG_0_d0, Y => un1_hwres_1_i);
    
    un4_so_7_0 : MUX2H
      port map(A => N_457, B => SP_PDL_in(20), S => REG_0(126), Y
         => N_458);
    
    un3_ae_39 : AND2
      port map(A => \un3_ae_1[39]\, B => \un3_ae_4[47]\, Y => 
        \un3_ae[39]\);
    
    SBYTE_136 : MUX2H
      port map(A => \SBYTE_5[7]_net_1\, B => \REG[144]\, S => 
        \un1_sstate_20\, Y => \SBYTE_136\);
    
    \sstate_0[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res\, Q => \sstate_0[9]_net_1\);
    
    un69_ae_6_0_2 : NOR2
      port map(A => \un69_ae_1[15]\, B => \un69_ae_2[47]\, Y => 
        \un69_ae_2[7]\);
    
    \AE_i_m[12]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_48\, B => \AE_0_sqmuxa_50\, C
         => \AE_PDL_c[12]\, Y => \AE_i_m[12]_net_1\);
    
    \P0_m[13]\ : AND2
      port map(A => \AE_0_sqmuxa_52\, B => \P0[13]_net_1\, Y => 
        \P0_m_i[13]\);
    
    \P0_50_iv[7]\ : NAND3
      port map(A => \P0_m[7]_net_1\, B => 
        \PDLCFG_DT_m_45[0]_net_1\, C => \REG_m_i[129]\, Y => 
        \P0_50[7]\);
    
    \P0[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_61\, CLR => 
        \un1_load_res_6\, Q => \P0[31]_net_1\);
    
    SBYTE_134 : MUX2H
      port map(A => \SBYTE_5[5]_net_1\, B => \REG[142]\, S => 
        \un1_sstate_20\, Y => \SBYTE_134\);
    
    \AE[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_105\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[25]\);
    
    \PDLCFG_DT_m_34[0]\ : NAND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[20]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_34[0]_net_1\);
    
    \P0_m[32]\ : AND2
      port map(A => \AE_0_sqmuxa_128\, B => \P0[32]_net_1\, Y => 
        \P0_m_i[32]\);
    
    \P0_50_iv[11]\ : NAND3FTT
      port map(A => \P0_m_i[11]\, B => \PDLCFG_DT_m_25[0]_net_1\, 
        C => \REG_m_i[129]\, Y => \P0_50[11]\);
    
    un69_ae_22_0 : NOR2
      port map(A => \un69_ae_1_i[30]\, B => \un69_ae_2[47]\, Y
         => un69_ae_30_0);
    
    \PDLCFG_RAD[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDLCFG_RAD_25\, CLR => 
        \un1_load_res_9\, Q => \PDLCFG_RAD[2]_net_1\);
    
    \AE_7_r[42]\ : AND3FFT
      port map(A => \AE_i_m[42]_net_1\, B => \REG_i_m[195]_net_1\, 
        C => N_6864_0, Y => \AE_7[42]\);
    
    \sstate_4[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_4[9]_net_1\);
    
    \P0_50_iv[25]\ : NAND3FTT
      port map(A => \P0_m_i[25]\, B => \PDLCFG_DT_m_9[0]_net_1\, 
        C => \REG_m_i_1[129]\, Y => \P0_50[25]\);
    
    \sstate_19_1_1_iv[6]\ : NAND3FTT
      port map(A => \sstate_19_1_1_iv_0_i[6]\, B => 
        \sstate_2_sqmuxa\, C => \ISI_0_sqmuxa\, Y => 
        \sstate_19_1[6]\);
    
    \P0[46]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_76\, CLR => 
        \un1_load_res_8\, Q => \P0[46]_net_1\);
    
    \PDLCFG_RAD_6_r[1]\ : AND2
      port map(A => N_502, B => \PDLCFG_RAD_1_sqmuxa\, Y => 
        \PDLCFG_RAD_6[1]_net_1\);
    
    \AE_i_m[40]\ : AOI21
      port map(A => \AE_0_sqmuxa_160\, B => \AE_0_sqmuxa_162\, C
         => \AE_PDL_c[40]\, Y => \AE_i_m[40]_net_1\);
    
    \P0[30]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_60\, CLR => 
        \un1_load_res_6\, Q => \P0[30]_net_1\);
    
    \sstate_19_0_iv[3]\ : OAI21FTT
      port map(A => \sstate[1]_net_1\, B => \un5_bitcnt\, C => 
        \sstate_0_sqmuxa\, Y => \sstate_19[3]\);
    
    AE_0_sqmuxa_96 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[24]\, Y => 
        \AE_0_sqmuxa_96\);
    
    PDL_RACK_22 : MUX2H
      port map(A => \un1_sstate_15\, B => PDL_RACK_net_1, S => 
        \un1_sstate_16\, Y => \PDL_RACK_22\);
    
    \P0_m[10]\ : AND2
      port map(A => \AE_0_sqmuxa_40\, B => \P0[10]_net_1\, Y => 
        \P0_m_i[10]\);
    
    \P0_m[23]\ : AND2
      port map(A => \AE_0_sqmuxa_92\, B => \P0[23]_net_1\, Y => 
        \P0_m_i[23]\);
    
    un3_ae_14_1 : OR2FT
      port map(A => \CNT[3]_net_1\, B => \CNT[0]_net_1\, Y => 
        \un3_ae_1[14]\);
    
    un1_sstate_1 : OR2
      port map(A => \sstate[1]_net_1\, B => \sstate[6]_net_1\, Y
         => \un1_sstate_1\);
    
    PDL_RDATA_16 : MUX2H
      port map(A => \PDL_RDATA[2]_net_1\, B => PDLCFG_DT(2), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_16\);
    
    AE_1_sqmuxa_0 : OR2FT
      port map(A => \sstate_0[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        \AE_1_sqmuxa_0\);
    
    un1_load_res_10 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_2, Y => 
        \un1_load_res_10\);
    
    \SBYTE_m[7]\ : AND2
      port map(A => \sstate[1]_net_1\, B => \REG[144]\, Y => 
        \SBYTE_m_i[7]\);
    
    \P0_m[6]\ : NAND2FT
      port map(A => \AE_0_sqmuxa_24\, B => \P0[6]_net_1\, Y => 
        \P0_m[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    AE_0_sqmuxa_102 : AO21
      port map(A => \un69_ae_1[25]\, B => \un69_ae_2[31]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_102\);
    
    AE_114 : MUX2H
      port map(A => \AE_PDL_c[34]\, B => \AE_7[34]\, S => 
        \un1_sstate_14_1\, Y => \AE_114\);
    
    AE_0_sqmuxa_120 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[30]\, Y => 
        \AE_0_sqmuxa_120\);
    
    \AE_i_m[31]\ : AOI21
      port map(A => \AE_0_sqmuxa_124\, B => \AE_0_sqmuxa_126\, C
         => \AE_PDL_c[31]\, Y => \AE_i_m[31]_net_1\);
    
    un3_ae_7 : NOR2FT
      port map(A => \un3_ae_1[7]\, B => \un3_ae_2[7]\, Y => 
        \un3_ae[7]\);
    
    ISI_1_sqmuxa_1 : NAND2
      port map(A => \sstate[6]_net_1\, B => \un3_pulse\, Y => 
        \ISI_1_sqmuxa_1\);
    
    \P0_m[20]\ : NAND2
      port map(A => \AE_0_sqmuxa_80\, B => \P0[20]_net_1\, Y => 
        \P0_m[20]_net_1\);
    
    \PDL_RDATA[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_19\, CLR => 
        \un1_load_res_10\, Q => \PDL_RDATA[5]_net_1\);
    
    AE_83 : MUX2H
      port map(A => \AE_PDL_c[3]\, B => \AE_7[3]\, S => 
        \un1_sstate_14\, Y => \AE_83\);
    
    un2_load_res : NOR2
      port map(A => LOAD_RES, B => HWRES_c_1, Y => un2_load_res_i);
    
    \sstate_2[6]\ : DFFB
      port map(CLK => CLK_c_c, D => \sstate_19_1[6]\, CLR => 
        un2_load_res_i, SET => HWRES_c_23_0, Q => 
        \sstate_2[6]_net_1\);
    
    \AE_7_r[11]\ : AND3FFT
      port map(A => \AE_i_m[11]_net_1\, B => \REG_i_m[164]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[11]\);
    
    AE_110 : MUX2H
      port map(A => \AE_PDL_c[30]\, B => \AE_7[30]\, S => 
        \un1_sstate_14_1\, Y => \AE_110\);
    
    \sstate[12]\ : DFFB
      port map(CLK => CLK_c_c, D => \GND\, CLR => HWRES_c_23_0, 
        SET => LOAD_RES_i_0, Q => \sstate[12]_net_1\);
    
    AE_0_sqmuxa_82 : AOI21
      port map(A => \un69_ae_1[23]\, B => \un69_ae_1[28]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_82\);
    
    \REG_i_m[194]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_73, Y => 
        \REG_i_m[194]_net_1\);
    
    \REG_i_m[165]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_44, Y => 
        \REG_i_m[165]_net_1\);
    
    \AE_i_m[26]\ : AOI21
      port map(A => \AE_0_sqmuxa_104\, B => \AE_0_sqmuxa_106\, C
         => \AE_PDL_c[26]\, Y => \AE_i_m[26]_net_1\);
    
    P_9 : MUX2H
      port map(A => \P_PDL_c[3]\, B => \P_4[3]_net_1\, S => 
        \un1_sstate_2\, Y => \P_9\);
    
    \P0_m[36]\ : NAND2
      port map(A => \AE_0_sqmuxa_144\, B => \P0[36]_net_1\, Y => 
        \P0_m[36]_net_1\);
    
    \sstate[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_19[0]\, CLR => 
        \un1_load_res_11\, Q => \sstate_i_i[0]\);
    
    un4_so_37_0 : MUX2H
      port map(A => SP_PDL_in(11), B => SP_PDL_in(15), S => REG_3, 
        Y => N_488);
    
    \REG_i_m[193]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_72, Y => 
        \REG_i_m[193]_net_1\);
    
    \REG_i_m[175]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_54, Y => 
        \REG_i_m[175]_net_1\);
    
    AE_0_sqmuxa_184 : NAND2
      port map(A => \sstate_4[9]_net_1\, B => \un3_ae[46]\, Y => 
        \AE_0_sqmuxa_184\);
    
    un4_so_13_0 : MUX2H
      port map(A => N_463, B => SP_PDL_in(18), S => REG_0(126), Y
         => N_464);
    
    \P[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \P_11\, CLR => 
        \un1_load_res_10\, Q => \P_PDL_c[5]\);
    
    AE_0_sqmuxa_74 : AOI21
      port map(A => \un69_ae_1[23]\, B => \un69_ae_1[26]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_74\);
    
    un3_ae_22 : OR2
      port map(A => \un3_ae_1[22]\, B => \un3_ae_2[47]\, Y => 
        \un3_ae[22]\);
    
    \PDLCFG_DT_m_3[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[43]\, Y => \PDLCFG_DT_m_3[0]_net_1\);
    
    un69_ae_38_1 : NOR2
      port map(A => \un69_ae_1_i[46]\, B => \un69_ae_2[47]\, Y
         => \un69_ae_1[38]\);
    
    un3_ae_42 : NAND2
      port map(A => \un3_ae_1[42]\, B => \un3_ae_3[47]\, Y => 
        \un3_ae[42]\);
    
    AE_95 : MUX2H
      port map(A => \AE_PDL_c[15]\, B => \AE_7[15]\, S => 
        \un1_sstate_14_2\, Y => \AE_95\);
    
    AE_0_sqmuxa_6 : AOI21
      port map(A => \un69_ae_1[7]\, B => \un69_ae_1[9]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_6\);
    
    VALID : DFFS
      port map(CLK => CLK_c_c, D => \VALID_29\, SET => 
        \un1_load_res_11\, Q => \REG[145]\);
    
    \P0[47]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_77\, CLR => 
        \un1_load_res_8\, Q => \P0[47]_net_1\);
    
    AE_0_sqmuxa_92 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[23]\, Y => 
        \AE_0_sqmuxa_92\);
    
    un3_ae_15_1 : OR2
      port map(A => \CNT[4]_net_1\, B => \CNT[5]_net_1\, Y => 
        \un3_ae_1[15]\);
    
    \P0_50_iv[32]\ : NAND3FFT
      port map(A => \P0_m_i[32]\, B => \PDLCFG_DT_m_16_i[0]\, C
         => \REG_m_i_1[129]\, Y => \P0_50[32]\);
    
    un69_ae_33_1 : NOR2
      port map(A => \un69_ae_1[41]\, B => \un69_ae_1_i[47]\, Y
         => \un69_ae_1[33]\);
    
    SBYTE_132 : MUX2H
      port map(A => \SBYTE_5[3]_net_1\, B => \REG[140]\, S => 
        \un1_sstate_20\, Y => \SBYTE_132\);
    
    un4_so_31_0 : MUX2H
      port map(A => SP_PDL_in(13), B => SP_PDL_in(45), S => REG_6, 
        Y => N_482);
    
    \AE_7_r[0]\ : AND3FFT
      port map(A => \AE_i_m[0]_net_1\, B => \REG_i_m[153]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[0]\);
    
    \P0_50_iv[18]\ : NAND3FFT
      port map(A => \PDLCFG_DT_m_32_i[0]\, B => \P0_m_i[18]\, C
         => \REG_m_i_2[129]\, Y => \P0_50[18]\);
    
    un3_ae_20 : NOR2
      port map(A => \un3_ae_1[22]\, B => \un3_ae_1[45]\, Y => 
        \un3_ae[20]\);
    
    \AE_7_r[23]\ : AND3FFT
      port map(A => \AE_i_m[23]_net_1\, B => \REG_i_m[176]_net_1\, 
        C => N_6864_2, Y => \AE_7[23]\);
    
    AE_0_sqmuxa_106 : AO21
      port map(A => \un69_ae_1[26]\, B => \un69_ae_2[31]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_106\);
    
    \AE[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_94\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[14]\);
    
    \PDLCFG_RAD_6_r[5]\ : AND2
      port map(A => N_506, B => \PDLCFG_RAD_1_sqmuxa\, Y => 
        \PDLCFG_RAD_6[5]_net_1\);
    
    \AE_i_m[4]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_16\, B => \AE_0_sqmuxa_18\, C
         => \AE_PDL_c[4]\, Y => \AE_i_m[4]_net_1\);
    
    un3_ae_40 : NAND2
      port map(A => \un3_ae_1[40]\, B => \un3_ae_3[47]\, Y => 
        \un3_ae[40]\);
    
    un69_ae_39_2 : NOR2
      port map(A => \un69_ae_1_i[47]\, B => \un69_ae_2[47]\, Y
         => \un69_ae_4[47]\);
    
    SBYTE_129 : MUX2H
      port map(A => \SBYTE_5[0]_net_1\, B => \REG[137]\, S => 
        \un1_sstate_20\, Y => \SBYTE_129\);
    
    un1_sstate_16 : OAI21
      port map(A => \sstate[6]_net_1\, B => \un1_sstate_3_0\, C
         => \PDL_RACK_1_sqmuxa\, Y => \un1_sstate_16\);
    
    \sstate_i_0[12]\ : INV
      port map(A => LOAD_RES, Y => LOAD_RES_i_0);
    
    un3_ae_38 : AND2
      port map(A => \un3_ae_1[39]\, B => \un3_ae_2[46]\, Y => 
        \un3_ae[38]\);
    
    un1_sstate_29_1 : NOR2
      port map(A => \PDLCFG_RAD_0_sqmuxa\, B => 
        \sstate[11]_net_1\, Y => \un1_sstate_29_1\);
    
    \sstate_19_1_1_iv_0[6]\ : OAI21FTT
      port map(A => \sstate_i_i[0]\, B => PDL_RREQ, C => 
        \sstate_i[7]\, Y => \sstate_19_1_1_iv_0_i[6]\);
    
    AE_0_sqmuxa_14 : OA21FTF
      port map(A => \un69_ae_1[5]\, B => \un69_ae_1[43]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_14\);
    
    \PDLCFG_RAD[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDLCFG_RAD_26\, CLR => 
        \un1_load_res_9\, Q => \PDLCFG_RAD[3]_net_1\);
    
    \AE_i_m[46]\ : AOI21
      port map(A => \AE_0_sqmuxa_184\, B => \AE_0_sqmuxa_186\, C
         => \AE_PDL_c[46]\, Y => \AE_i_m[46]_net_1\);
    
    \REG_i_m[188]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_67, Y => 
        \REG_i_m[188]_net_1\);
    
    \AE_7_r[9]\ : AND3FFT
      port map(A => \AE_i_m[9]_net_1\, B => \REG_i_m[162]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[9]\);
    
    AE_0_sqmuxa_190 : AO21
      port map(A => \un69_ae_3[47]\, B => \un69_ae_4[47]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_190\);
    
    \AE_i_m[18]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_72\, B => \AE_0_sqmuxa_74\, C
         => \AE_PDL_c[18]\, Y => \AE_i_m[18]_net_1\);
    
    \P0_m[17]\ : AND2
      port map(A => \AE_0_sqmuxa_68\, B => \P0[17]_net_1\, Y => 
        \P0_m_i[17]\);
    
    sstate_2_sqmuxa : OR2
      port map(A => \ISI_1_sqmuxa_1\, B => PDL_RREQ, Y => 
        \sstate_2_sqmuxa\);
    
    \P0_50_iv[13]\ : NAND3FFT
      port map(A => \PDLCFG_DT_m_27_i[0]\, B => \P0_m_i[13]\, C
         => \REG_m_i_2[129]\, Y => \P0_50[13]\);
    
    \P0[34]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_64\, CLR => 
        \un1_load_res_7\, Q => \P0[34]_net_1\);
    
    \AE[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_98\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[18]\);
    
    \REG_i_m[164]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_43, Y => 
        \REG_i_m[164]_net_1\);
    
    \AE[40]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_120\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[40]\);
    
    AE_109 : MUX2H
      port map(A => \AE_PDL_c[29]\, B => \AE_7[29]\, S => 
        \un1_sstate_14_1\, Y => \AE_109\);
    
    un69_ae_31_1 : OR2FT
      port map(A => REG_1, B => REG_0(127), Y => 
        \un69_ae_1_i[31]\);
    
    un4_so_19_0 : MUX2H
      port map(A => SP_PDL_in(14), B => SP_PDL_in(46), S => REG_6, 
        Y => N_470);
    
    un3_ae_10_1 : NOR2
      port map(A => \un3_ae_1[15]\, B => \un3_ae_1_i[43]\, Y => 
        \un3_ae_1[11]\);
    
    \PDLCFG_DT_m_13[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[29]\, Y => \PDLCFG_DT_m_13[0]_net_1\);
    
    AE_0_sqmuxa_130 : AOI21
      port map(A => \un69_ae_1[39]\, B => \un69_ae_1[40]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_130\);
    
    \REG_i_m[163]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_42, Y => 
        \REG_i_m[163]_net_1\);
    
    AE_0_sqmuxa_24 : NAND2
      port map(A => \sstate_8[9]_net_1\, B => \un3_ae[6]\, Y => 
        \AE_0_sqmuxa_24\);
    
    \REG_i_m[174]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_53, Y => 
        \REG_i_m[174]_net_1\);
    
    \P0_m[27]\ : AND2FT
      port map(A => \AE_0_sqmuxa_108\, B => \P0[27]_net_1\, Y => 
        \P0_m_i[27]\);
    
    \AE_7_r[5]\ : AND3FFT
      port map(A => \AE_i_m[5]_net_1\, B => \REG_i_m[158]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[5]\);
    
    un4_so_16_0 : MUX2H
      port map(A => N_464, B => N_469, S => REG_0(124), Y => 
        N_467_i_i);
    
    \REG_i_m[173]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_52, Y => 
        \REG_i_m[173]_net_1\);
    
    PDLCFG_RAD_26 : MUX2H
      port map(A => \PDLCFG_RAD_6[3]_net_1\, B => 
        \PDLCFG_RAD[3]_net_1\, S => \un1_sstate_25\, Y => 
        \PDLCFG_RAD_26\);
    
    ISCK : DFFC
      port map(CLK => CLK_c_c, D => \ISCK_128\, CLR => 
        \un1_load_res_4\, Q => \SCLK_PDL_c\);
    
    \REG_i_m[186]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_65, Y => 
        \REG_i_m[186]_net_1\);
    
    \PDL_RDATA[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_20\, CLR => 
        \un1_load_res_10\, Q => \PDL_RDATA[6]_net_1\);
    
    \P0_50_iv[20]\ : NAND3
      port map(A => \P0_m[20]_net_1\, B => 
        \PDLCFG_DT_m_34[0]_net_1\, C => \REG_m_i_2[129]\, Y => 
        \P0_50[20]\);
    
    un4_so_6_0 : MUX2H
      port map(A => SP_PDL_in(4), B => SP_PDL_in(36), S => 
        REG_0(127), Y => N_457);
    
    un3_ae_15_2 : NAND2
      port map(A => \CNT[0]_net_1\, B => \CNT[3]_net_1\, Y => 
        \un3_ae_2[15]\);
    
    un69_ae_12_0 : NOR2FT
      port map(A => \un69_ae_1[14]\, B => \un69_ae_1[45]\, Y => 
        \un69_ae_12_0\);
    
    \AE_7_r[4]\ : AND3FFT
      port map(A => \AE_i_m[4]_net_1\, B => \REG_i_m[157]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[4]\);
    
    AE_0_sqmuxa_50 : OA21FTF
      port map(A => \un69_ae_12_0\, B => \un69_ae_1[15]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_50\);
    
    un1_sstate_25 : OAI21TTF
      port map(A => \sstate[11]_net_1\, B => \sstate_1[6]_net_1\, 
        C => \PDLCFG_RAD_0_sqmuxa_1\, Y => \un1_sstate_25\);
    
    AE_0_sqmuxa_40 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[10]\, Y => 
        \AE_0_sqmuxa_40\);
    
    un4_so_25_0 : MUX2H
      port map(A => N_475, B => SP_PDL_in(17), S => REG_5, Y => 
        N_476);
    
    \P0_50_iv[42]\ : NAND3FTT
      port map(A => \P0_m_i[42]\, B => \PDLCFG_DT_m_2[0]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[42]\);
    
    P0_44 : MUX2H
      port map(A => \P0[14]_net_1\, B => \P0_50[14]\, S => 
        \un1_sstate_2_3\, Y => \P0_44\);
    
    un4_so_32_0 : MUX2H
      port map(A => SP_PDL_in(25), B => SP_PDL_in(29), S => REG_3, 
        Y => N_483);
    
    \AE_7_r[29]\ : AND3FFT
      port map(A => \AE_i_m[29]_net_1\, B => \REG_i_m[182]_net_1\, 
        C => N_6864_1, Y => \AE_7[29]\);
    
    un3_ae_21 : NOR2FT
      port map(A => un3_ae_21_0, B => \un3_ae_1[23]\, Y => 
        \un3_ae[21]\);
    
    \P0_50_iv[15]\ : NAND3
      port map(A => \P0_m[15]_net_1\, B => 
        \PDLCFG_DT_m_29[0]_net_1\, C => \REG_m_i_2[129]\, Y => 
        \P0_50[15]\);
    
    P0_38 : MUX2H
      port map(A => \P0[8]_net_1\, B => \P0_50[8]\, S => 
        \un1_sstate_2_3\, Y => \P0_38\);
    
    \P0_50_iv[39]\ : NAND3FFT
      port map(A => \P0_m_i[39]\, B => \PDLCFG_DT_m_i[0]\, C => 
        \REG_m_i_0[129]\, Y => \P0_50[39]\);
    
    \AE_i_m[27]\ : AOI21
      port map(A => \AE_0_sqmuxa_108\, B => \AE_0_sqmuxa_110\, C
         => \AE_PDL_c[27]\, Y => \AE_i_m[27]_net_1\);
    
    P0_54 : MUX2H
      port map(A => \P0[24]_net_1\, B => \P0_50[24]\, S => 
        \un1_sstate_2_2\, Y => \P0_54\);
    
    \AE[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_104\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[24]\);
    
    un3_ae_41 : NAND2
      port map(A => \un3_ae_1[33]\, B => \un3_ae_3[47]\, Y => 
        \un3_ae[41]\);
    
    \AE_i_m[9]\ : AOI21
      port map(A => \AE_0_sqmuxa_36\, B => \AE_0_sqmuxa_38\, C
         => \AE_PDL_c[9]\, Y => \AE_i_m[9]_net_1\);
    
    \PDLCFG_DT_m_8[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[24]\, Y => \PDLCFG_DT_m_8[0]_net_1\);
    
    \P0[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_53\, CLR => 
        \un1_load_res_6\, Q => \P0[23]_net_1\);
    
    CNT_2_I_22 : XOR2
      port map(A => \CNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => \CNT_2[2]\);
    
    \AE_7_r[20]\ : AND3FFT
      port map(A => \AE_i_m[20]_net_1\, B => \REG_i_m[173]_net_1\, 
        C => N_6864_2, Y => \AE_7[20]\);
    
    un69_ae_47_1 : OR2FT
      port map(A => REG_1, B => REG_0(126), Y => 
        \un69_ae_1_i[47]\);
    
    CNT_2_I_23 : XOR2
      port map(A => \CNT[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => \CNT_2[3]\);
    
    \P0[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_43\, CLR => 
        \un1_load_res_5\, Q => \P0[13]_net_1\);
    
    \AE_i_m[25]\ : AOI21
      port map(A => \AE_0_sqmuxa_100\, B => \AE_0_sqmuxa_102\, C
         => \AE_PDL_c[25]\, Y => \AE_i_m[25]_net_1\);
    
    P0_64 : MUX2H
      port map(A => \P0[34]_net_1\, B => \P0_50[34]\, S => 
        \un1_sstate_2_1\, Y => \P0_64\);
    
    un4_so_30_0 : MUX2H
      port map(A => N_480, B => SP_PDL_in(21), S => REG_5, Y => 
        N_481);
    
    P0_41 : MUX2H
      port map(A => \P0[11]_net_1\, B => \P0_50[11]\, S => 
        \un1_sstate_2_3\, Y => \P0_41\);
    
    un1_sstate_14_2 : OR3
      port map(A => \un1_sstate_5\, B => \sstate_0[9]_net_1\, C
         => \sstate[11]_net_1\, Y => \un1_sstate_14_2\);
    
    \P0[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_34\, CLR => 
        \un1_load_res_8\, Q => \P0[4]_net_1\);
    
    AE_0_sqmuxa_34 : AOI21
      port map(A => \un69_ae_1[9]\, B => \un69_ae_1[14]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_34\);
    
    un3_ae_25 : NAND2
      port map(A => \un3_ae_1[25]\, B => \un3_ae_2[31]\, Y => 
        \un3_ae[25]\);
    
    P0_42 : MUX2H
      port map(A => \P0[12]_net_1\, B => \P0_50[12]\, S => 
        \un1_sstate_2_3\, Y => \P0_42\);
    
    \P0[28]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_58\, CLR => 
        \un1_load_res_6\, Q => \P0[28]_net_1\);
    
    un3_ae_45 : NAND2
      port map(A => \un3_ae_3[47]\, B => un3_ae_45_0, Y => 
        \un3_ae[45]\);
    
    PDLCFG_RAD_25 : MUX2H
      port map(A => \PDLCFG_RAD_6[2]_net_1\, B => 
        \PDLCFG_RAD[2]_net_1\, S => \un1_sstate_25\, Y => 
        \PDLCFG_RAD_25\);
    
    P0_51 : MUX2H
      port map(A => \P0[21]_net_1\, B => \P0_50[21]\, S => 
        \un1_sstate_2_2\, Y => \P0_51\);
    
    AE_117 : MUX2H
      port map(A => \AE_PDL_c[37]\, B => \AE_7[37]\, S => 
        \un1_sstate_14_0\, Y => \AE_117\);
    
    \P0[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_35\, CLR => 
        \un1_load_res_8\, Q => \P0[5]_net_1\);
    
    \AE[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_83\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[3]\);
    
    P0_52 : MUX2H
      port map(A => \P0[22]_net_1\, B => \P0_50[22]\, S => 
        \un1_sstate_2_2\, Y => \P0_52\);
    
    \AE[35]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_115\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[35]\);
    
    \AE[28]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_108\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[28]\);
    
    \P0[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_48\, CLR => 
        \un1_load_res_5\, Q => \P0[18]_net_1\);
    
    \P_4[4]\ : MUX2H
      port map(A => REG_12, B => PDLCFG_DT(4), S => 
        \sstate[9]_net_1\, Y => \P_4[4]_net_1\);
    
    \PDLCFG_DT_m_33[0]\ : AND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[19]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_33_i[0]\);
    
    \PDLCFG_DT_m_12[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[28]\, Y => \PDLCFG_DT_m_12[0]_net_1\);
    
    P0_61 : MUX2H
      port map(A => \P0[31]_net_1\, B => \P0_50[31]\, S => 
        \un1_sstate_2_1\, Y => \P0_61\);
    
    \P0[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_36\, CLR => 
        \un1_load_res_8\, Q => \P0[6]_net_1\);
    
    P0_62 : MUX2H
      port map(A => \P0[32]_net_1\, B => \P0_50[32]\, S => 
        \un1_sstate_2_1\, Y => \P0_62\);
    
    MODE : DFFB
      port map(CLK => CLK_c_c, D => \MODE_0\, CLR => 
        un1_hwres_1_i, SET => \un1_reg_1_i\, Q => MD_PDL_c);
    
    \P0_m[18]\ : AND2
      port map(A => \AE_0_sqmuxa_72\, B => \P0[18]_net_1\, Y => 
        \P0_m_i[18]\);
    
    \AE_i_m[0]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_0\, B => \AE_0_sqmuxa_2\, C => 
        \AE_PDL_c[0]\, Y => \AE_i_m[0]_net_1\);
    
    un4_so_38_0 : MUX2H
      port map(A => N_488, B => N_493, S => REG_6, Y => N_489);
    
    AE_108 : MUX2H
      port map(A => \AE_PDL_c[28]\, B => \AE_7[28]\, S => 
        \un1_sstate_14_1\, Y => \AE_108\);
    
    \SBYTE[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_133\, CLR => 
        \un1_load_res_11\, Q => \REG[141]\);
    
    un69_ae_30_1 : OR2
      port map(A => REG_1, B => REG_0(127), Y => 
        \un69_ae_1_i[30]\);
    
    \AE_7_r[32]\ : AND3FFT
      port map(A => \AE_i_m[32]_net_1\, B => \REG_i_m[185]_net_1\, 
        C => N_6864_1, Y => \AE_7[32]\);
    
    \sstate[7]\ : DFFS
      port map(CLK => CLK_c_c, D => \PDLCFG_RAD_0_sqmuxa_1_i\, 
        SET => \un1_load_res\, Q => \sstate_i[7]\);
    
    un69_ae_7_1 : NOR2FT
      port map(A => REG_1, B => REG_0(125), Y => \un69_ae_1[7]\);
    
    PDL_RDATA_19 : MUX2H
      port map(A => \PDL_RDATA[5]_net_1\, B => PDLCFG_DT(5), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_19\);
    
    \AE_i_m[47]\ : AOI21
      port map(A => \AE_0_sqmuxa_188\, B => \AE_0_sqmuxa_190\, C
         => \AE_PDL_c[47]\, Y => \AE_i_m[47]_net_1\);
    
    AE_91 : MUX2H
      port map(A => \AE_PDL_c[11]\, B => \AE_7[11]\, S => 
        \un1_sstate_14\, Y => \AE_91\);
    
    \REG_m_46_2[129]\ : NAND2
      port map(A => \sstate_0[6]_net_1\, B => REG_8, Y => 
        \REG_m_i_2[129]\);
    
    PDLCFG_RAD_0_sqmuxa : AND2
      port map(A => \sstate_1[6]_net_1\, B => PDL_RREQ, Y => 
        \PDLCFG_RAD_0_sqmuxa\);
    
    \PDL_RDATA[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_16\, CLR => 
        \un1_load_res_9\, Q => \PDL_RDATA[2]_net_1\);
    
    \PDLCFG_DT_m_6[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[46]\, Y => \PDLCFG_DT_m_6[0]_net_1\);
    
    \sstate[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[9]_net_1\, CLR => 
        \un1_load_res\, Q => \sstate[8]_net_1\);
    
    \P0_m[28]\ : AND2FT
      port map(A => \AE_0_sqmuxa_112\, B => \P0[28]_net_1\, Y => 
        \P0_m_i[28]\);
    
    un69_ae_0_0 : AND2FT
      port map(A => \un69_ae_1[41]\, B => \un69_ae_1[6]\, Y => 
        \un69_ae_0_0\);
    
    un4_so_34_0 : MUX2H
      port map(A => N_479_i, B => N_484_i, S => REG_4, Y => N_485);
    
    \AE_i_m[45]\ : AOI21
      port map(A => \AE_0_sqmuxa_180\, B => \AE_0_sqmuxa_182\, C
         => \AE_PDL_c[45]\, Y => \AE_i_m[45]_net_1\);
    
    AE_124 : MUX2H
      port map(A => \AE_PDL_c[44]\, B => \AE_7[44]\, S => 
        \un1_sstate_14_0\, Y => \AE_124\);
    
    \PDLCFG_DT_m_2[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[42]\, Y => \PDLCFG_DT_m_2[0]_net_1\);
    
    \P0_50_iv[27]\ : NAND3FTT
      port map(A => \P0_m_i[27]\, B => \PDLCFG_DT_m_11[0]_net_1\, 
        C => \REG_m_i_1[129]\, Y => \P0_50[27]\);
    
    un3_pulse : OR2FT
      port map(A => PULSE(8), B => \MD_PDL_c_0\, Y => \un3_pulse\);
    
    \REG_i_m[159]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_38, Y => 
        \REG_i_m[159]_net_1\);
    
    AE_120 : MUX2H
      port map(A => \AE_PDL_c[40]\, B => \AE_7[40]\, S => 
        \un1_sstate_14_0\, Y => \AE_120\);
    
    AE_0_sqmuxa_66 : AOI21
      port map(A => \un69_ae_1[23]\, B => \un69_ae_1[24]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_66\);
    
    \AE_i_m[14]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_56\, B => \AE_0_sqmuxa_58\, C
         => \AE_PDL_c[14]\, Y => \AE_i_m[14]_net_1\);
    
    un69_ae_34_1 : NOR2
      port map(A => \un69_ae_1[43]\, B => \un69_ae_1_i[46]\, Y
         => \un69_ae_1[42]\);
    
    \P0[29]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_59\, CLR => 
        \un1_load_res_6\, Q => \P0[29]_net_1\);
    
    AE_0_sqmuxa_188 : NAND2
      port map(A => \sstate_4[9]_net_1\, B => \un3_ae[47]\, Y => 
        \AE_0_sqmuxa_188\);
    
    \P[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \P_8\, CLR => 
        \un1_load_res_10\, Q => \P_PDL_c[2]\);
    
    \P0_m[31]\ : AND2FT
      port map(A => \AE_0_sqmuxa_124\, B => \P0[31]_net_1\, Y => 
        \P0_m_i[31]\);
    
    \P0[36]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_66\, CLR => 
        \un1_load_res_7\, Q => \P0[36]_net_1\);
    
    \P0[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_49\, CLR => 
        \un1_load_res_5\, Q => \P0[19]_net_1\);
    
    \AE_7_r[44]\ : AND3FFT
      port map(A => \AE_i_m[44]_net_1\, B => \REG_i_m[197]_net_1\, 
        C => N_6864_0, Y => \AE_7[44]\);
    
    AE_0_sqmuxa_170 : AO21
      port map(A => \un69_ae_1[42]\, B => \un69_ae_3[47]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_170\);
    
    \AE_i_m[33]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_132\, B => \AE_0_sqmuxa_134\, C
         => \AE_PDL_c[33]\, Y => \AE_i_m[33]_net_1\);
    
    PDLCFG_RAD_23 : MUX2H
      port map(A => \PDLCFG_RAD_6[0]_net_1\, B => 
        \PDLCFG_RAD[0]_net_1\, S => \un1_sstate_25\, Y => 
        \PDLCFG_RAD_23\);
    
    \PDL_RACK\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RACK_22\, CLR => 
        \un1_load_res_9\, Q => PDL_RACK_net_1);
    
    \AE[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_81\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[1]\);
    
    \P0_m[44]\ : NAND2FT
      port map(A => \AE_0_sqmuxa_176\, B => \P0[44]_net_1\, Y => 
        \P0_m[44]_net_1\);
    
    un4_so_23_0 : MUX2H
      port map(A => N_462, B => N_473, S => REG_2, Y => N_474);
    
    \AE_7_r[13]\ : AND3FFT
      port map(A => \AE_i_m[13]_net_1\, B => \REG_i_m[166]_net_1\, 
        C => N_6864_2, Y => \AE_7[13]\);
    
    \AE_7_r[26]\ : AND3FFT
      port map(A => \AE_i_m[26]_net_1\, B => \REG_i_m[179]_net_1\, 
        C => N_6864_1, Y => \AE_7[26]\);
    
    \PDLCFG_DT_m_32[0]\ : AND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[18]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_32_i[0]\);
    
    AE_104 : MUX2H
      port map(A => \AE_PDL_c[24]\, B => \AE_7[24]\, S => 
        \un1_sstate_14_1\, Y => \AE_104\);
    
    un3_ae_23_2 : NOR2
      port map(A => \un3_ae_1_i[31]\, B => \un3_ae_2[47]\, Y => 
        \un3_ae_3[31]\);
    
    \PDLCFG_RAD_6_r[0]\ : AND2
      port map(A => N_501, B => \PDLCFG_RAD_1_sqmuxa\, Y => 
        \PDLCFG_RAD_6[0]_net_1\);
    
    \P0[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_38\, CLR => 
        \un1_load_res_8\, Q => \P0[8]_net_1\);
    
    un3_ae_46_2 : NOR2
      port map(A => \un3_ae_1_i[46]\, B => \un3_ae_2[47]\, Y => 
        \un3_ae_2[46]\);
    
    un4_so_45_0 : MUX2H
      port map(A => N_490_i, B => N_495_i, S => REG_4, Y => N_496);
    
    un4_so_1_0 : MUX2H
      port map(A => SP_PDL_in(0), B => SP_PDL_in(32), S => 
        REG_0(127), Y => N_452);
    
    \P_4[6]\ : MUX2H
      port map(A => REG_14, B => PDLCFG_DT(6), S => 
        \sstate_8[9]_net_1\, Y => \P_4[6]_net_1\);
    
    \P0_50_iv[36]\ : NAND3FTT
      port map(A => \PDLCFG_DT_m_20_i[0]\, B => \P0_m[36]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[36]\);
    
    \BITCNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_5[1]\, CLR => 
        \un1_load_res_4\, Q => \BITCNT[1]_net_1\);
    
    AE_100 : MUX2H
      port map(A => \AE_PDL_c[20]\, B => \AE_7[20]\, S => 
        \un1_sstate_14_2\, Y => \AE_100\);
    
    \AE[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_90\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[10]\);
    
    MODE_2_0 : DFFB
      port map(CLK => CLK_c_c, D => \MODE_0\, CLR => 
        un1_hwres_1_i, SET => \un1_reg_1_i\, Q => MD_PDL_c_2);
    
    \AE[42]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_122\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[42]\);
    
    un3_ae_2_1 : OR2FT
      port map(A => \un3_ae_1[6]\, B => \un3_ae_1[15]\, Y => 
        \un3_ae_1[2]\);
    
    \PDLCFG_DT_m_16[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[32]\, C => 
        \sstate_6[9]_net_1\, Y => \PDLCFG_DT_m_16_i[0]\);
    
    \P0_m[3]\ : NAND2
      port map(A => \AE_0_sqmuxa_12\, B => \P0[3]_net_1\, Y => 
        \P0_m[3]_net_1\);
    
    un69_ae_3_0_1 : NOR2FT
      port map(A => \un69_ae_1[7]\, B => \un69_ae_1[15]\, Y => 
        \un69_ae_1[5]\);
    
    \SBYTE_5[3]\ : MUX2H
      port map(A => \REG[139]\, B => REG_11, S => 
        \sstate_2[6]_net_1\, Y => \SBYTE_5[3]_net_1\);
    
    \sstate_5[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_5[9]_net_1\);
    
    un3_ae_6 : OR2FT
      port map(A => \un3_ae_1[6]\, B => \un3_ae_2[7]\, Y => 
        \un3_ae[6]\);
    
    \REG_i_m[157]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_36, Y => 
        \REG_i_m[157]_net_1\);
    
    \P0_50_iv[10]\ : NAND3FFT
      port map(A => \PDLCFG_DT_m_24_i[0]\, B => \P0_m_i[10]\, C
         => \REG_m_i[129]\, Y => \P0_50[10]\);
    
    AE_0_sqmuxa_150 : AOI21
      port map(A => \un69_ae_1[39]\, B => un69_ae_37_0, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_150\);
    
    un69_ae_15_1 : OR2
      port map(A => REG_0(127), B => REG_0(126), Y => 
        \un69_ae_1[15]\);
    
    PDL_RACK_1_sqmuxa : NAND2
      port map(A => \sstate_i_i[0]\, B => PDL_RREQ, Y => 
        \PDL_RACK_1_sqmuxa\);
    
    un3_ae_39_2 : NOR2
      port map(A => \un3_ae_1_i[47]\, B => \un3_ae_2[47]\, Y => 
        \un3_ae_4[47]\);
    
    \PDLCFG_DT_m_19[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[35]\, C => 
        \sstate_5[9]_net_1\, Y => \PDLCFG_DT_m_19_i[0]\);
    
    \P0_m[39]\ : AND2
      port map(A => \AE_0_sqmuxa_156\, B => \P0[39]_net_1\, Y => 
        \P0_m_i[39]\);
    
    ISI : DFFC
      port map(CLK => CLK_c_c, D => \ISI_78\, CLR => 
        \un1_load_res_4\, Q => \SI_PDL_c\);
    
    AE_0_sqmuxa_62 : AOI21
      port map(A => \un69_ae_2[7]\, B => \un69_ae_2[15]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_62\);
    
    un3_ae_29_0 : NOR2
      port map(A => \un3_ae_1_i[31]\, B => \un3_ae_1[45]\, Y => 
        un3_ae_21_0);
    
    SO : NOR2
      port map(A => un4_so, B => \REG[145]\, Y => \SO\);
    
    \P0_m[7]\ : NAND2
      port map(A => \AE_0_sqmuxa_28\, B => \P0[7]_net_1\, Y => 
        \P0_m[7]_net_1\);
    
    sstate_1_sqmuxa : AND2
      port map(A => \PDLCFG_RAD_0_sqmuxa\, B => \un3_pulse\, Y
         => \sstate_19[5]\);
    
    \AE_7_r_i_2[47]\ : NOR2
      port map(A => \sstate[12]_net_1\, B => \sstate[11]_net_1\, 
        Y => N_6864_2);
    
    \P0[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_30\, CLR => 
        \un1_load_res_4\, Q => \P0[0]_net_1\);
    
    \P0[37]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_67\, CLR => 
        \un1_load_res_7\, Q => \P0[37]_net_1\);
    
    un4_so_29_0 : MUX2H
      port map(A => SP_PDL_in(5), B => SP_PDL_in(37), S => REG_6, 
        Y => N_480);
    
    \AE_7_r[3]\ : AND3FFT
      port map(A => \AE_i_m[3]_net_1\, B => \REG_i_m[156]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[3]\);
    
    \REG_m_46_0[129]\ : NAND2
      port map(A => \sstate_0[6]_net_1\, B => REG_8, Y => 
        \REG_m_i_0[129]\);
    
    \AE_i_m[39]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_156\, B => \AE_0_sqmuxa_158\, C
         => \AE_PDL_c[39]\, Y => \AE_i_m[39]_net_1\);
    
    un3_ae_29 : NAND2
      port map(A => \un3_ae_2[31]\, B => un3_ae_21_0, Y => 
        \un3_ae[29]\);
    
    AE_85 : MUX2H
      port map(A => \AE_PDL_c[5]\, B => \AE_7[5]\, S => 
        \un1_sstate_14\, Y => \AE_85\);
    
    \AE_7_r[38]\ : AND3FFT
      port map(A => \AE_i_m[38]_net_1\, B => \REG_i_m[191]_net_1\, 
        C => N_6864_0, Y => \AE_7[38]\);
    
    PDLCFG_nRD_79 : MUX2H
      port map(A => \un1_sstate_29_1\, B => PDLCFG_nRD_net_1, S
         => \un1_sstate_27\, Y => \PDLCFG_nRD_79\);
    
    \AE_7_r[19]\ : AND3FFT
      port map(A => \AE_i_m[19]_net_1\, B => \REG_i_m[172]_net_1\, 
        C => N_6864_2, Y => \AE_7[19]\);
    
    un4_so_26_0 : MUX2H
      port map(A => SP_PDL_in(9), B => SP_PDL_in(41), S => REG_6, 
        Y => N_477);
    
    \PDLCFG_RAD_6_r[4]\ : AND2
      port map(A => N_505, B => \PDLCFG_RAD_1_sqmuxa\, Y => 
        \PDLCFG_RAD_6[4]_net_1\);
    
    \P0_m[43]\ : AND2FT
      port map(A => \AE_0_sqmuxa_172\, B => \P0[43]_net_1\, Y => 
        \P0_m_i[43]\);
    
    P0_35 : MUX2H
      port map(A => \P0[5]_net_1\, B => \P0_50[5]\, S => 
        \un1_sstate_2_3\, Y => \P0_35\);
    
    un3_ae_17 : NOR2FT
      port map(A => \un3_ae_1[25]\, B => \un3_ae_1[23]\, Y => 
        \un3_ae[17]\);
    
    AE_113 : MUX2H
      port map(A => \AE_PDL_c[33]\, B => \AE_7[33]\, S => 
        \un1_sstate_14_1\, Y => \AE_113\);
    
    SBYTE_130 : MUX2H
      port map(A => \SBYTE_5[1]_net_1\, B => \REG[138]\, S => 
        \un1_sstate_20\, Y => \SBYTE_130\);
    
    AE_0_sqmuxa_4 : NOR2FT
      port map(A => \sstate_0[9]_net_1\, B => \un3_ae[1]\, Y => 
        \AE_0_sqmuxa_4\);
    
    \AE_i_m[30]\ : AOI21
      port map(A => \AE_0_sqmuxa_120\, B => \AE_0_sqmuxa_122\, C
         => \AE_PDL_c[30]\, Y => \AE_i_m[30]_net_1\);
    
    AE_0_sqmuxa_104 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[26]\, Y => 
        \AE_0_sqmuxa_104\);
    
    \sstate_0[6]\ : DFFB
      port map(CLK => CLK_c_c, D => \sstate_19_1[6]\, CLR => 
        un2_load_res_i, SET => HWRES_c_23_0, Q => 
        \sstate_0[6]_net_1\);
    
    un3_ae_37_0 : NOR2
      port map(A => \un3_ae_1[45]\, B => \un3_ae_1_i[47]\, Y => 
        un3_ae_45_0);
    
    \AE_7_r[10]\ : AND3FFT
      port map(A => \AE_i_m[10]_net_1\, B => \REG_i_m[163]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[10]\);
    
    \P0_50_iv[46]\ : NAND3FTT
      port map(A => \P0_m_i[46]\, B => \PDLCFG_DT_m_6[0]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[46]\);
    
    AE_0_sqmuxa_112 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[28]\, Y => 
        \AE_0_sqmuxa_112\);
    
    P0_75 : MUX2H
      port map(A => \P0[45]_net_1\, B => \P0_50[45]\, S => 
        \un1_sstate_2_0\, Y => \P0_75\);
    
    \AE_i_m[3]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_12\, B => \AE_0_sqmuxa_14\, C
         => \AE_PDL_c[3]\, Y => \AE_i_m[3]_net_1\);
    
    AE_116 : MUX2H
      port map(A => \AE_PDL_c[36]\, B => \AE_7[36]\, S => 
        \un1_sstate_14_0\, Y => \AE_116\);
    
    \P0_m[40]\ : AND2FT
      port map(A => \AE_0_sqmuxa_160\, B => \P0[40]_net_1\, Y => 
        \P0_m_i[40]\);
    
    \AE[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_100\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[20]\);
    
    \sstate_1[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_1[9]_net_1\);
    
    \P0_m[5]\ : NAND2FT
      port map(A => \AE_0_sqmuxa_20\, B => \P0[5]_net_1\, Y => 
        \P0_m[5]_net_1\);
    
    un1_sstate_2_1 : OR2
      port map(A => \sstate_0[9]_net_1\, B => \sstate_0[6]_net_1\, 
        Y => \un1_sstate_2_1\);
    
    \AE[34]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_114\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[34]\);
    
    \P0[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_52\, CLR => 
        \un1_load_res_6\, Q => \P0[22]_net_1\);
    
    \PDLCFG_DT_m_36[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[22]\, Y => \PDLCFG_DT_m_36[0]_net_1\);
    
    \SBYTE_5[0]\ : MUX2H
      port map(A => \SO\, B => REG_8, S => \sstate_2[6]_net_1\, Y
         => \SBYTE_5[0]_net_1\);
    
    \P0[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_42\, CLR => 
        \un1_load_res_5\, Q => \P0[12]_net_1\);
    
    un1_sstate_27_0 : NAND2FT
      port map(A => \sstate[8]_net_1\, B => \sstate_i[7]\, Y => 
        un1_sstate_27_0_i);
    
    un3_ae_41_1 : OR2
      port map(A => \CNT[2]_net_1\, B => \CNT[1]_net_1\, Y => 
        \un3_ae_1[41]\);
    
    un69_ae_2_0_1 : NOR2FT
      port map(A => \un69_ae_1[6]\, B => \un69_ae_1[15]\, Y => 
        \un69_ae_1[4]\);
    
    CNT_2_I_30 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \CNT[4]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    CNT_2_I_24 : XOR2
      port map(A => \CNT[4]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => \CNT_2[4]\);
    
    \PDLCFG_DT_m_39[0]\ : AND3
      port map(A => PDLCFG_DT(0), B => \un3_ae[1]\, C => 
        \sstate_8[9]_net_1\, Y => \PDLCFG_DT_m_39_i[0]\);
    
    AE_0_sqmuxa_162 : AO21
      port map(A => \un69_ae_1[40]\, B => \un69_ae_3[47]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_162\);
    
    \AE_7_r[27]\ : AND3FFT
      port map(A => \AE_i_m[27]_net_1\, B => \REG_i_m[180]_net_1\, 
        C => N_6864_1, Y => \AE_7[27]\);
    
    PDL_RDATA_15 : MUX2H
      port map(A => \PDL_RDATA[1]_net_1\, B => PDLCFG_DT(1), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_15\);
    
    PDL_RDATA_18 : MUX2H
      port map(A => \PDL_RDATA[4]_net_1\, B => PDLCFG_DT(4), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_18\);
    
    PDLCFG_RAD_0_sqmuxa_1_i : INV
      port map(A => \PDLCFG_RAD_0_sqmuxa_1\, Y => 
        \PDLCFG_RAD_0_sqmuxa_1_i\);
    
    P0_30 : MUX2H
      port map(A => \P0[0]_net_1\, B => \P0_50[0]\, S => 
        \un1_sstate_2\, Y => \P0_30\);
    
    \sstate_8[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res_0_0\, Q => \sstate_8[9]_net_1\);
    
    AE_0_sqmuxa_78 : AOI21
      port map(A => \un69_ae_1[23]\, B => \un69_ae_1[27]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_78\);
    
    un4_so_43_0 : MUX2H
      port map(A => SP_PDL_in(27), B => SP_PDL_in(31), S => REG_3, 
        Y => N_494);
    
    \AE[38]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_118\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[38]\);
    
    AE_127 : MUX2H
      port map(A => \AE_PDL_c[47]\, B => \AE_7[47]\, S => 
        \un1_sstate_14_0\, Y => \AE_127\);
    
    \P0_50_iv[17]\ : NAND3FFT
      port map(A => \P0_m_i[17]\, B => \PDLCFG_DT_m_31_i[0]\, C
         => \REG_m_i_2[129]\, Y => \P0_50[17]\);
    
    \CNT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_2[4]\, CLR => 
        \un1_load_res_4\, Q => \CNT[4]_net_1\);
    
    AE_0_sqmuxa_140 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[35]\, Y => 
        \AE_0_sqmuxa_140\);
    
    \AE_7_r[25]\ : AND3FFT
      port map(A => \AE_i_m[25]_net_1\, B => \REG_i_m[178]_net_1\, 
        C => N_6864_1, Y => \AE_7[25]\);
    
    un1_load_res_11 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_2, Y => 
        \un1_load_res_11\);
    
    un3_ae_20_1 : OR2
      port map(A => \un3_ae_1[30]\, B => \un3_ae_1[23]\, Y => 
        \un3_ae_1[22]\);
    
    \AE[41]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_121\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[41]\);
    
    un1_sstate_2_2 : OR2
      port map(A => \sstate_0[9]_net_1\, B => \sstate_0[6]_net_1\, 
        Y => \un1_sstate_2_2\);
    
    AE_0_sqmuxa_84 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[21]\, Y => 
        \AE_0_sqmuxa_84\);
    
    P0_70 : MUX2H
      port map(A => \P0[40]_net_1\, B => \P0_50[40]\, S => 
        \un1_sstate_2_0\, Y => \P0_70\);
    
    \CNT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_2[5]\, CLR => 
        \un1_load_res_4\, Q => \CNT[5]_net_1\);
    
    un5_bitcnt : AND3
      port map(A => \BITCNT[0]_net_1\, B => \BITCNT[1]_net_1\, C
         => \BITCNT[2]_net_1\, Y => \un5_bitcnt\);
    
    un69_ae_32_1 : NOR2
      port map(A => \un69_ae_1[41]\, B => \un69_ae_1_i[46]\, Y
         => \un69_ae_1[40]\);
    
    un4_so_5_0 : MUX2H
      port map(A => N_453, B => N_458, S => REG_0(124), Y => 
        N_456_i_i);
    
    \REG_i_m[191]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_70, Y => 
        \REG_i_m[191]_net_1\);
    
    \AE_i_m[11]\ : AOI21
      port map(A => \AE_0_sqmuxa_44\, B => \AE_0_sqmuxa_46\, C
         => \AE_PDL_c[11]\, Y => \AE_i_m[11]_net_1\);
    
    \SBYTE_5[4]\ : MUX2H
      port map(A => \REG[140]\, B => REG_12, S => 
        \sstate_2[6]_net_1\, Y => \SBYTE_5[4]_net_1\);
    
    AE_92 : MUX2H
      port map(A => \AE_PDL_c[12]\, B => \AE_7[12]\, S => 
        \un1_sstate_14_2\, Y => \AE_92\);
    
    \SBYTE[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_131\, CLR => 
        \un1_load_res_11\, Q => \REG[139]\);
    
    AE_0_sqmuxa_116 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[29]\, Y => 
        \AE_0_sqmuxa_116\);
    
    CNT_2_I_31 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \CNT[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    \P0[45]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_75\, CLR => 
        \un1_load_res_8\, Q => \P0[45]_net_1\);
    
    \AE_7_r_i[47]\ : NOR2
      port map(A => \sstate[12]_net_1\, B => \sstate[11]_net_1\, 
        Y => \AE_7_r_i[47]_net_1\);
    
    un1_load_res_5 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_3, Y => 
        \un1_load_res_5\);
    
    AE_0_sqmuxa_18 : OA21FTF
      port map(A => \un69_ae_1[4]\, B => \un69_ae_1[45]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_18\);
    
    un3_ae_31_2 : AND2
      port map(A => \CNT[3]_net_1\, B => \CNT[4]_net_1\, Y => 
        \un3_ae_2[31]\);
    
    AE_97 : MUX2H
      port map(A => \AE_PDL_c[17]\, B => \AE_7[17]\, S => 
        \un1_sstate_14_2\, Y => \AE_97\);
    
    \AE_7_r[41]\ : AND3FFT
      port map(A => \AE_i_m[41]_net_1\, B => \REG_i_m[194]_net_1\, 
        C => N_6864_0, Y => \AE_7[41]\);
    
    AE_107 : MUX2H
      port map(A => \AE_PDL_c[27]\, B => \AE_7[27]\, S => 
        \un1_sstate_14_1\, Y => \AE_107\);
    
    un69_ae_1_0_1 : NOR2
      port map(A => \un69_ae_1[15]\, B => \un69_ae_1[41]\, Y => 
        \un69_ae_1[9]\);
    
    \P0_50_iv[5]\ : NAND3
      port map(A => \PDLCFG_DT_m_43[0]_net_1\, B => 
        \P0_m[5]_net_1\, C => \REG_m_i[129]\, Y => \P0_50[5]\);
    
    \AE_i_m[36]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_144\, B => \AE_0_sqmuxa_146\, C
         => \AE_PDL_c[36]\, Y => \AE_i_m[36]_net_1\);
    
    \P0_50_iv[3]\ : NAND3FTT
      port map(A => \PDLCFG_DT_m_41_i[0]\, B => \P0_m[3]_net_1\, 
        C => \REG_m_i[129]\, Y => \P0_50[3]\);
    
    AE_0_sqmuxa_94 : AOI21
      port map(A => \un69_ae_1[23]\, B => \un69_ae_3[31]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_94\);
    
    AE_0_sqmuxa_166 : AO21
      port map(A => \un69_ae_1[33]\, B => \un69_ae_3[47]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_166\);
    
    \AE_7_r[16]\ : AND3FFT
      port map(A => \AE_i_m[16]_net_1\, B => \REG_i_m[169]_net_1\, 
        C => N_6864_2, Y => \AE_7[16]\);
    
    SBYTE_135 : MUX2H
      port map(A => \SBYTE_5[6]_net_1\, B => \REG[143]\, S => 
        \un1_sstate_20\, Y => \SBYTE_135\);
    
    P_8 : MUX2H
      port map(A => \P_PDL_c[2]\, B => \P_4[2]_net_1\, S => 
        \un1_sstate_2\, Y => \P_8\);
    
    \PDLCFG_DT_m[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[39]\, C => 
        \sstate_5[9]_net_1\, Y => \PDLCFG_DT_m_i[0]\);
    
    AE_0_sqmuxa_122 : AO21
      port map(A => \un69_ae_2[31]\, B => un69_ae_30_0, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_122\);
    
    AE_0_sqmuxa_28 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[7]\, Y => 
        \AE_0_sqmuxa_28\);
    
    \AE[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_92\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[12]\);
    
    \P0_m[47]\ : AND2FT
      port map(A => \AE_0_sqmuxa_188\, B => \P0[47]_net_1\, Y => 
        \P0_m_i[47]\);
    
    un3_ae_28 : OR3FTT
      port map(A => \un3_ae_2[31]\, B => \un3_ae_1[30]\, C => 
        \un3_ae_1[45]\, Y => \un3_ae[28]\);
    
    \AE_i_m[1]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_4\, B => \AE_0_sqmuxa_6\, C => 
        \AE_PDL_c[1]\, Y => \AE_i_m[1]_net_1\);
    
    AE_1_sqmuxa : OR2FT
      port map(A => \sstate_1[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        \AE_1_sqmuxa\);
    
    \P0_m[35]\ : AND2
      port map(A => \AE_0_sqmuxa_140\, B => \P0[35]_net_1\, Y => 
        \P0_m_i[35]\);
    
    AE_90 : MUX2H
      port map(A => \AE_PDL_c[10]\, B => \AE_7[10]\, S => 
        \un1_sstate_14\, Y => \AE_90\);
    
    un4_so_46_0 : MUX2H
      port map(A => N_485, B => N_496, S => REG_2, Y => N_497);
    
    \sstate[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[5]_net_1\, CLR => 
        \un1_load_res\, Q => \sstate[4]_net_1\);
    
    \P0_m[12]\ : AND2
      port map(A => \AE_0_sqmuxa_48\, B => \P0[12]_net_1\, Y => 
        \P0_m_i[12]\);
    
    \AE_7_r[34]\ : AND3FFT
      port map(A => \AE_i_m[34]_net_1\, B => \REG_i_m[187]_net_1\, 
        C => N_6864_1, Y => \AE_7[34]\);
    
    \PDLCFG_RAD[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDLCFG_RAD_28\, CLR => 
        \un1_load_res_9\, Q => \PDLCFG_RAD[5]_net_1\);
    
    un69_ae_15_2 : AND2
      port map(A => REG_1, B => REG_4, Y => \un69_ae_2[15]\);
    
    un1_load_res : OR2FT
      port map(A => LOAD_RES, B => HWRES_c_0, Y => \un1_load_res\);
    
    AE_81 : MUX2H
      port map(A => \AE_PDL_c[1]\, B => \AE_7[1]\, S => 
        \un1_sstate_14\, Y => \AE_81\);
    
    un3_ae_0 : NOR3FTT
      port map(A => \un3_ae_1[6]\, B => \un3_ae_1[15]\, C => 
        \un3_ae_1[41]\, Y => \un3_ae[0]\);
    
    AE_94 : MUX2H
      port map(A => \AE_PDL_c[14]\, B => \AE_7[14]\, S => 
        \un1_sstate_14_2\, Y => \AE_94\);
    
    un4_so_2_0 : MUX2H
      port map(A => N_452, B => SP_PDL_in(16), S => REG_0(126), Y
         => N_453);
    
    un3_ae_34_1 : NOR2
      port map(A => \un3_ae_1_i[43]\, B => \un3_ae_1_i[46]\, Y
         => \un3_ae_1[42]\);
    
    \SBYTE[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_134\, CLR => 
        \un1_load_res_11\, Q => \REG[142]\);
    
    \P0_m[22]\ : NAND2FT
      port map(A => \AE_0_sqmuxa_88\, B => \P0[22]_net_1\, Y => 
        \P0_m[22]_net_1\);
    
    \REG_i_m[161]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_40, Y => 
        \REG_i_m[161]_net_1\);
    
    P0_37 : MUX2H
      port map(A => \P0[7]_net_1\, B => \P0_50[7]\, S => 
        \un1_sstate_2_3\, Y => \P0_37\);
    
    \BITCNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_5[2]\, CLR => 
        \un1_load_res_4\, Q => \BITCNT[2]_net_1\);
    
    AE_98 : MUX2H
      port map(A => \AE_PDL_c[18]\, B => \AE_7[18]\, S => 
        \un1_sstate_14_2\, Y => \AE_98\);
    
    \AE[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_85\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[5]\);
    
    \REG_i_m[171]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_50, Y => 
        \REG_i_m[171]_net_1\);
    
    \AE_7_r_i_0[47]\ : NOR2
      port map(A => \sstate[12]_net_1\, B => \sstate[11]_net_1\, 
        Y => N_6864_0);
    
    un3_ae_16 : NOR2FT
      port map(A => \un3_ae_1[24]\, B => \un3_ae_1[23]\, Y => 
        \un3_ae[16]\);
    
    \sstate_1[6]\ : DFFB
      port map(CLK => CLK_c_c, D => \sstate_19_1[6]\, CLR => 
        un2_load_res_i, SET => HWRES_c_23_0, Q => 
        \sstate_1[6]_net_1\);
    
    \SBYTE[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_136\, CLR => 
        \un1_load_res_11\, Q => \REG[144]\);
    
    AE_0_sqmuxa_38 : AO21
      port map(A => \un69_ae_1[9]\, B => \un69_ae_2[15]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_38\);
    
    ISI_5_r : OA21TTF
      port map(A => \REG_m_i[136]\, B => \SBYTE_m_i[7]\, C => 
        \un1_sstate_22\, Y => ISI_5);
    
    AE_0_sqmuxa_56 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[14]\, Y => 
        \AE_0_sqmuxa_56\);
    
    P0_77 : MUX2H
      port map(A => \P0[47]_net_1\, B => \P0_50[47]\, S => 
        \un1_sstate_2_0\, Y => \P0_77\);
    
    \sstate[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[2]_net_1\, CLR => 
        \un1_load_res_11\, Q => \sstate[1]_net_1\);
    
    \REG_i_m[192]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_71, Y => 
        \REG_i_m[192]_net_1\);
    
    \sstate[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[10]_net_1\, CLR => 
        \un1_load_res\, Q => \sstate[9]_net_1\);
    
    AE_0_sqmuxa_46 : AO21
      port map(A => \un69_ae_1[11]\, B => \un69_ae_2[15]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_46\);
    
    PDL_RDATA_20 : MUX2H
      port map(A => \PDL_RDATA[6]_net_1\, B => PDLCFG_DT(6), S
         => \sstate[4]_net_1\, Y => \PDL_RDATA_20\);
    
    un1_sstate_27_3 : OR3
      port map(A => \sstate_i_i[0]\, B => un1_sstate_27_0_i, C
         => \sstate[2]_net_1\, Y => un1_sstate_27_3_i);
    
    AE_0_sqmuxa_126 : AO21
      port map(A => \un69_ae_2[31]\, B => \un69_ae_3[31]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_126\);
    
    \AE_7_r[6]\ : AND3FFT
      port map(A => \AE_i_m[6]_net_1\, B => \REG_i_m[159]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[6]\);
    
    un1_BITCNT_I_13 : XOR2
      port map(A => \BITCNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_13_5);
    
    \P0_m[16]\ : AND2
      port map(A => \AE_0_sqmuxa_64\, B => \P0[16]_net_1\, Y => 
        \P0_m_i[16]\);
    
    N_387_i_a2 : NOR2
      port map(A => \ISI_0_sqmuxa\, B => \sstate[6]_net_1\, Y => 
        N_389);
    
    \REG_i_m[185]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_64, Y => 
        \REG_i_m[185]_net_1\);
    
    \P0[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_39\, CLR => 
        \un1_load_res_8\, Q => \P0[9]_net_1\);
    
    \REG_i_m[190]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_69, Y => 
        \REG_i_m[190]_net_1\);
    
    un1_sstate_3_0 : OR2
      port map(A => \sstate[4]_net_1\, B => \sstate_i_i[0]\, Y
         => \un1_sstate_3_0\);
    
    \AE[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_102\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[22]\);
    
    AE_0_sqmuxa_108 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[27]\, Y => 
        \AE_0_sqmuxa_108\);
    
    un3_ae_46_1 : OR2
      port map(A => \CNT[0]_net_1\, B => \CNT[4]_net_1\, Y => 
        \un3_ae_1_i[46]\);
    
    \P[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \P_13\, CLR => 
        \un1_load_res_10\, Q => \P_PDL_c[7]\);
    
    \P0_m[1]\ : NAND2
      port map(A => \AE_0_sqmuxa_4\, B => \P0[1]_net_1\, Y => 
        \P0_m[1]_net_1\);
    
    \sstate[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[3]_net_1\, CLR => 
        \un1_load_res_11\, Q => \sstate[2]_net_1\);
    
    AE_123 : MUX2H
      port map(A => \AE_PDL_c[43]\, B => \AE_7[43]\, S => 
        \un1_sstate_14_0\, Y => \AE_123\);
    
    AE_0_sqmuxa_132 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[33]\, Y => 
        \AE_0_sqmuxa_132\);
    
    \P0_m[26]\ : AND2FT
      port map(A => \AE_0_sqmuxa_104\, B => \P0[26]_net_1\, Y => 
        \P0_m_i[26]\);
    
    \REG_i_m[199]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_78, Y => 
        \REG_i_m[199]_net_1\);
    
    un3_ae_13 : NOR3
      port map(A => \un3_ae_1[45]\, B => \un3_ae_2[15]\, C => 
        \un3_ae_1[15]\, Y => \un3_ae[13]\);
    
    \AE[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_80\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[0]\);
    
    un3_ae_43_1 : OR2FT
      port map(A => \CNT[1]_net_1\, B => \CNT[2]_net_1\, Y => 
        \un3_ae_1_i[43]\);
    
    un3_ae_1 : AND2
      port map(A => \un3_ae_1[7]\, B => \un3_ae_1[9]\, Y => 
        \un3_ae[1]\);
    
    un3_ae_35_1 : NOR2
      port map(A => \un3_ae_1_i[43]\, B => \un3_ae_1_i[47]\, Y
         => \un3_ae_2[43]\);
    
    \AE_i_m[37]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_148\, B => \AE_0_sqmuxa_150\, C
         => \AE_PDL_c[37]\, Y => \AE_i_m[37]_net_1\);
    
    \AE[30]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_110\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[30]\);
    
    AE_111 : MUX2H
      port map(A => \AE_PDL_c[31]\, B => \AE_7[31]\, S => 
        \un1_sstate_14_1\, Y => \AE_111\);
    
    AE_126 : MUX2H
      port map(A => \AE_PDL_c[46]\, B => \AE_7[46]\, S => 
        \un1_sstate_14_0\, Y => \AE_126\);
    
    un3_ae_5 : OR2
      port map(A => \un3_ae_1[5]\, B => \un3_ae_1[45]\, Y => 
        \un3_ae[5]\);
    
    \P0[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_51\, CLR => 
        \un1_load_res_6\, Q => \P0[21]_net_1\);
    
    \AE_7_r[17]\ : AND3FFT
      port map(A => \AE_i_m[17]_net_1\, B => \REG_i_m[170]_net_1\, 
        C => N_6864_2, Y => \AE_7[17]\);
    
    \AE[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_91\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[11]\);
    
    \AE[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_99\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[19]\);
    
    \P0[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_41\, CLR => 
        \un1_load_res_5\, Q => \P0[11]_net_1\);
    
    \AE_i_m[35]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_140\, B => \AE_0_sqmuxa_142\, C
         => \AE_PDL_c[35]\, Y => \AE_i_m[35]_net_1\);
    
    \P0_50_iv[6]\ : NAND3
      port map(A => \P0_m[6]_net_1\, B => 
        \PDLCFG_DT_m_44[0]_net_1\, C => \REG_m_i[129]\, Y => 
        \P0_50[6]\);
    
    \P0_50_iv[22]\ : NAND3
      port map(A => \P0_m[22]_net_1\, B => 
        \PDLCFG_DT_m_36[0]_net_1\, C => \REG_m_i_2[129]\, Y => 
        \P0_50[22]\);
    
    \AE[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_89\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[9]\);
    
    un69_ae_47_3 : AND2
      port map(A => REG_4, B => REG_6, Y => \un69_ae_3[47]\);
    
    \AE_7_r[15]\ : AND3FFT
      port map(A => \AE_i_m[15]_net_1\, B => \REG_i_m[168]_net_1\, 
        C => N_6864_2, Y => \AE_7[15]\);
    
    AE_0_sqmuxa_52 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[13]\, Y => 
        \AE_0_sqmuxa_52\);
    
    \P0[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_50\, CLR => 
        \un1_load_res_5\, Q => \P0[20]_net_1\);
    
    AE_115 : MUX2H
      port map(A => \AE_PDL_c[35]\, B => \AE_7[35]\, S => 
        \un1_sstate_14_1\, Y => \AE_115\);
    
    AE_0_sqmuxa_42 : AOI21
      port map(A => \un69_ae_1[11]\, B => \un69_ae_1[14]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_42\);
    
    \PDLCFG_DT_m_21[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[37]\, C => 
        \sstate_5[9]_net_1\, Y => \PDLCFG_DT_m_21_i[0]\);
    
    \P0[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_40\, CLR => 
        \un1_load_res_5\, Q => \P0[10]_net_1\);
    
    \REG_i_m[162]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_41, Y => 
        \REG_i_m[162]_net_1\);
    
    \PDLCFG_DT_m_41[0]\ : AND3
      port map(A => PDLCFG_DT(0), B => \un3_ae[3]\, C => 
        \sstate_8[9]_net_1\, Y => \PDLCFG_DT_m_41_i[0]\);
    
    AE_103 : MUX2H
      port map(A => \AE_PDL_c[23]\, B => \AE_7[23]\, S => 
        \un1_sstate_14_2\, Y => \AE_103\);
    
    un3_ae_37 : AND2
      port map(A => \un3_ae_1[39]\, B => un3_ae_45_0, Y => 
        \un3_ae[37]\);
    
    \SBYTE_5[7]\ : MUX2H
      port map(A => \REG[143]\, B => REG_15, S => 
        \sstate_1[6]_net_1\, Y => \SBYTE_5[7]_net_1\);
    
    un3_ae_14 : NOR2
      port map(A => \un3_ae_1[14]\, B => \un3_ae_2[7]\, Y => 
        \un3_ae[14]\);
    
    \AE_i_m[8]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_32\, B => \AE_0_sqmuxa_34\, C
         => \AE_PDL_c[8]\, Y => \AE_i_m[8]_net_1\);
    
    \REG_i_m[184]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_63, Y => 
        \REG_i_m[184]_net_1\);
    
    \REG_i_m[172]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_51, Y => 
        \REG_i_m[172]_net_1\);
    
    un3_ae_30_1 : OR2
      port map(A => \CNT[0]_net_1\, B => \CNT[5]_net_1\, Y => 
        \un3_ae_1[30]\);
    
    \REG_i_m[160]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_39, Y => 
        \REG_i_m[160]_net_1\);
    
    un3_ae_9 : OR2FT
      port map(A => \un3_ae_1[9]\, B => \un3_ae_2[15]\, Y => 
        \un3_ae[9]\);
    
    \P0_m[0]\ : AND2
      port map(A => \AE_0_sqmuxa_0\, B => \P0[0]_net_1\, Y => 
        \P0_m_i[0]\);
    
    AE_106 : MUX2H
      port map(A => \AE_PDL_c[26]\, B => \AE_7[26]\, S => 
        \un1_sstate_14_1\, Y => \AE_106\);
    
    un1_sstate_15 : NOR2
      port map(A => \sstate_i_i[0]\, B => \sstate[6]_net_1\, Y
         => \un1_sstate_15\);
    
    \REG_i_m[183]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_62, Y => 
        \REG_i_m[183]_net_1\);
    
    MODE_0_0 : DFFB
      port map(CLK => CLK_c_c, D => \MODE_0\, CLR => 
        un1_hwres_1_i, SET => \un1_reg_1_i\, Q => \MD_PDL_c_0\);
    
    AE_0_sqmuxa_136 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[34]\, Y => 
        \AE_0_sqmuxa_136\);
    
    \REG_i_m[197]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_76, Y => 
        \REG_i_m[197]_net_1\);
    
    \AE_i_m[22]\ : AOI21
      port map(A => \AE_0_sqmuxa_88\, B => \AE_0_sqmuxa_90\, C
         => \AE_PDL_c[22]\, Y => \AE_i_m[22]_net_1\);
    
    un1_sstate_27_2 : OR2
      port map(A => \sstate[3]_net_1\, B => \sstate[1]_net_1\, Y
         => un1_sstate_27_2_i);
    
    \REG_i_m[170]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_49, Y => 
        \REG_i_m[170]_net_1\);
    
    un1_cnt : NOR3
      port map(A => \un3_ae_1[41]\, B => \un3_ae_1[23]\, C => 
        \un1_cnt_0\, Y => \un1_cnt\);
    
    \REG_i_m[169]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_48, Y => 
        \REG_i_m[169]_net_1\);
    
    \PDLCFG_DT_m_25[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[11]\, Y => \PDLCFG_DT_m_25[0]_net_1\);
    
    \PDLCFG_DT_m_45[0]\ : NAND3
      port map(A => PDLCFG_DT(0), B => \un3_ae[7]\, C => 
        \sstate_8[9]_net_1\, Y => \PDLCFG_DT_m_45[0]_net_1\);
    
    VALID_29 : MUX2H
      port map(A => \REG[145]\, B => \un1_sstate_22\, S => 
        \un1_sstate_5\, Y => \VALID_29\);
    
    \AE[46]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_126\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[46]\);
    
    \AE_i_m[2]\ : AOI21
      port map(A => \AE_0_sqmuxa_8\, B => \AE_0_sqmuxa_10\, C => 
        \AE_PDL_c[2]\, Y => \AE_i_m[2]_net_1\);
    
    un1_BITCNT_I_15 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \BITCNT[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1_0[0]\);
    
    \REG_i_m[179]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_58, Y => 
        \REG_i_m[179]_net_1\);
    
    \sstate_19_0_iv[0]\ : NAND2FT
      port map(A => \sstate[4]_net_1\, B => \PDL_RACK_1_sqmuxa\, 
        Y => \sstate_19[0]\);
    
    un69_ae_47_2 : NAND2
      port map(A => REG_2, B => REG_3, Y => \un69_ae_2[47]\);
    
    un1_sstate_13_0 : OR2
      port map(A => \sstate[12]_net_1\, B => \sstate[2]_net_1\, Y
         => \un1_sstate_13_0\);
    
    P0_46 : MUX2H
      port map(A => \P0[16]_net_1\, B => \P0_50[16]\, S => 
        \un1_sstate_2_2\, Y => \P0_46\);
    
    CNT_2_I_28 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_0[0]\, B => 
        \CNT[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    P0_49 : MUX2H
      port map(A => \P0[19]_net_1\, B => \P0_50[19]\, S => 
        \un1_sstate_2_2\, Y => \P0_49\);
    
    CNT_2_I_15 : XOR2
      port map(A => \CNT[0]_net_1\, B => \sstate[9]_net_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\);
    
    \AE[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_101\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[21]\);
    
    SBYTE_131 : MUX2H
      port map(A => \SBYTE_5[2]_net_1\, B => \REG[139]\, S => 
        \un1_sstate_20\, Y => \SBYTE_131\);
    
    \AE_i_m[13]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_52\, B => \AE_0_sqmuxa_54\, C
         => \AE_PDL_c[13]\, Y => \AE_i_m[13]_net_1\);
    
    \AE[29]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_109\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[29]\);
    
    \AE_7_r[31]\ : AND3FFT
      port map(A => \AE_i_m[31]_net_1\, B => \REG_i_m[184]_net_1\, 
        C => N_6864_1, Y => \AE_7[31]\);
    
    \REG_i_m[158]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_37, Y => 
        \REG_i_m[158]_net_1\);
    
    PDLCFG_RAD_1_sqmuxa : OR2FT
      port map(A => \sstate_1[6]_net_1\, B => PDL_RREQ, Y => 
        \PDLCFG_RAD_1_sqmuxa\);
    
    P0_56 : MUX2H
      port map(A => \P0[26]_net_1\, B => \P0_50[26]\, S => 
        \un1_sstate_2_1\, Y => \P0_56\);
    
    P0_59 : MUX2H
      port map(A => \P0[29]_net_1\, B => \P0_50[29]\, S => 
        \un1_sstate_2_1\, Y => \P0_59\);
    
    \REG_m_46[129]\ : NAND2
      port map(A => \sstate_2[6]_net_1\, B => REG_8, Y => 
        \REG_m_i[129]\);
    
    un1_load_res_2 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_3, Y => 
        \un1_load_res_2\);
    
    \AE_7_r[7]\ : AND3FFT
      port map(A => \AE_i_m[7]_net_1\, B => \REG_i_m[160]_net_1\, 
        C => \AE_7_r_i[47]_net_1\, Y => \AE_7[7]\);
    
    \P0_50_iv[29]\ : NAND3
      port map(A => \PDLCFG_DT_m_13[0]_net_1\, B => 
        \P0_m[29]_net_1\, C => \REG_m_i_1[129]\, Y => \P0_50[29]\);
    
    \AE_7_r[43]\ : AND3FFT
      port map(A => \AE_i_m[43]_net_1\, B => \REG_i_m[196]_net_1\, 
        C => N_6864_0, Y => \AE_7[43]\);
    
    P0_66 : MUX2H
      port map(A => \P0[36]_net_1\, B => \P0_50[36]\, S => 
        \un1_sstate_2_1\, Y => \P0_66\);
    
    P0_69 : MUX2H
      port map(A => \P0[39]_net_1\, B => \P0_50[39]\, S => 
        \un1_sstate_2_0\, Y => \P0_69\);
    
    \AE_i_m[42]\ : AOI21
      port map(A => \AE_0_sqmuxa_168\, B => \AE_0_sqmuxa_170\, C
         => \AE_PDL_c[42]\, Y => \AE_i_m[42]_net_1\);
    
    \P[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \P_9\, CLR => 
        \un1_load_res_10\, Q => \P_PDL_c[3]\);
    
    \P0_50_iv[1]\ : NAND3FTT
      port map(A => \PDLCFG_DT_m_39_i[0]\, B => \P0_m[1]_net_1\, 
        C => \REG_m_i[129]\, Y => \P0_50[1]\);
    
    \P0[35]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_65\, CLR => 
        \un1_load_res_7\, Q => \P0[35]_net_1\);
    
    AE_0_sqmuxa_70 : AOI21
      port map(A => \un69_ae_1[23]\, B => \un69_ae_1[25]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_70\);
    
    AE_0_sqmuxa_64 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[16]\, Y => 
        \AE_0_sqmuxa_64\);
    
    \PDL_RDATA[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_17\, CLR => 
        \un1_load_res_9\, Q => \PDL_RDATA[3]_net_1\);
    
    AE_0_sqmuxa_172 : NAND2
      port map(A => \sstate_5[9]_net_1\, B => \un3_ae[43]\, Y => 
        \AE_0_sqmuxa_172\);
    
    AE_0_sqmuxa_114 : AO21
      port map(A => \un69_ae_1[28]\, B => \un69_ae_2[31]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_114\);
    
    AE_82 : MUX2H
      port map(A => \AE_PDL_c[2]\, B => \AE_7[2]\, S => 
        \un1_sstate_14\, Y => \AE_82\);
    
    \REG_i_m[167]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_46, Y => 
        \REG_i_m[167]_net_1\);
    
    un1_load_res_0_0 : OR2FT
      port map(A => LOAD_RES_0, B => HWRES_c_0, Y => 
        \un1_load_res_0_0\);
    
    un69_ae_16_1 : NOR2
      port map(A => \un69_ae_1_i[30]\, B => \un69_ae_1[41]\, Y
         => \un69_ae_1[24]\);
    
    \REG_i_m[156]\ : NOR2
      port map(A => AE_0_sqmuxa_i, B => REG_35, Y => 
        \REG_i_m[156]_net_1\);
    
    \P0[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_54\, CLR => 
        \un1_load_res_6\, Q => \P0[24]_net_1\);
    
    un69_ae_45_1 : OR2FT
      port map(A => REG_0(124), B => REG_2, Y => \un69_ae_1[45]\);
    
    un3_ae_47_1 : OR2FT
      port map(A => \CNT[0]_net_1\, B => \CNT[4]_net_1\, Y => 
        \un3_ae_1_i[47]\);
    
    AE_87 : MUX2H
      port map(A => \AE_PDL_c[7]\, B => \AE_7[7]\, S => 
        \un1_sstate_14\, Y => \AE_87\);
    
    un4_so_17_0 : MUX2H
      port map(A => SP_PDL_in(6), B => SP_PDL_in(38), S => REG_6, 
        Y => N_468);
    
    \P0_50_iv[34]\ : NAND3FFT
      port map(A => \P0_m_i[34]\, B => \PDLCFG_DT_m_18_i[0]\, C
         => \REG_m_i_1[129]\, Y => \P0_50[34]\);
    
    \P0[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_44\, CLR => 
        \un1_load_res_5\, Q => \P0[14]_net_1\);
    
    AE_112 : MUX2H
      port map(A => \AE_PDL_c[32]\, B => \AE_7[32]\, S => 
        \un1_sstate_14_1\, Y => \AE_112\);
    
    \REG_i_m[177]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_56, Y => 
        \REG_i_m[177]_net_1\);
    
    un3_ae_16_1 : NOR2
      port map(A => \un3_ae_1[30]\, B => \un3_ae_1[41]\, Y => 
        \un3_ae_1[24]\);
    
    un1_BITCNT_I_1 : AND2
      port map(A => \BITCNT[0]_net_1\, B => \un1_sstate_21\, Y
         => \DWACT_ADD_CI_0_TMP[0]\);
    
    P0_34 : MUX2H
      port map(A => \P0[4]_net_1\, B => \P0_50[4]\, S => 
        \un1_sstate_2_3\, Y => \P0_34\);
    
    \PDLCFG_DT_m_28[0]\ : NAND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[14]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_28[0]_net_1\);
    
    \AE[47]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_127\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[47]\);
    
    un4_so_10_0_i : INV
      port map(A => N_461_i_i, Y => N_461_i);
    
    \AE[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_84\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[4]\);
    
    AE_0_sqmuxa_164 : NAND2
      port map(A => \sstate_5[9]_net_1\, B => \un3_ae[41]\, Y => 
        \AE_0_sqmuxa_164\);
    
    un3_ae_3_1 : OR2FT
      port map(A => \un3_ae_1[7]\, B => \un3_ae_1[15]\, Y => 
        \un3_ae_1[5]\);
    
    AE_0_sqmuxa_10 : OAI21FTF
      port map(A => \un69_ae_1[4]\, B => \un69_ae_1[43]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_10\);
    
    \PDLCFG_DT_m_20[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[36]\, C => 
        \sstate_5[9]_net_1\, Y => \PDLCFG_DT_m_20_i[0]\);
    
    \AE_i_m[19]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_76\, B => \AE_0_sqmuxa_78\, C
         => \AE_PDL_c[19]\, Y => \AE_i_m[19]_net_1\);
    
    \PDLCFG_DT_m_40[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_2(0), C
         => \un3_ae[2]\, Y => \PDLCFG_DT_m_40[0]_net_1\);
    
    un4_so_35_0 : MUX2H
      port map(A => SP_PDL_in(3), B => SP_PDL_in(35), S => REG_6, 
        Y => N_486);
    
    P0_74 : MUX2H
      port map(A => \P0[44]_net_1\, B => \P0_50[44]\, S => 
        \un1_sstate_2_0\, Y => \P0_74\);
    
    P0_31 : MUX2H
      port map(A => \P0[1]_net_1\, B => \P0_50[1]\, S => 
        \un1_sstate_2\, Y => \P0_31\);
    
    \P0[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_33\, CLR => 
        \un1_load_res_7\, Q => \P0[3]_net_1\);
    
    P0_32 : MUX2H
      port map(A => \P0[2]_net_1\, B => \P0_50[2]\, S => 
        \un1_sstate_2\, Y => \P0_32\);
    
    AE_0_sqmuxa_180 : NAND2
      port map(A => \sstate_4[9]_net_1\, B => \un3_ae[45]\, Y => 
        \AE_0_sqmuxa_180\);
    
    un4_so_11_0 : MUX2H
      port map(A => N_456_i, B => N_461_i, S => REG_0(125), Y => 
        N_462);
    
    \P0_m[11]\ : AND2FT
      port map(A => \AE_0_sqmuxa_44\, B => \P0[11]_net_1\, Y => 
        \P0_m_i[11]\);
    
    AE_80 : MUX2H
      port map(A => \AE_PDL_c[0]\, B => \AE_7[0]\, S => 
        \un1_sstate_14\, Y => \AE_80\);
    
    AE_0_sqmuxa_152 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[38]\, Y => 
        \AE_0_sqmuxa_152\);
    
    \AE[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_87\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[7]\);
    
    \AE_i_m[10]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_40\, B => \AE_0_sqmuxa_42\, C
         => \AE_PDL_c[10]\, Y => \AE_i_m[10]_net_1\);
    
    \AE_i_m[28]\ : AOI21
      port map(A => \AE_0_sqmuxa_112\, B => \AE_0_sqmuxa_114\, C
         => \AE_PDL_c[28]\, Y => \AE_i_m[28]_net_1\);
    
    \AE[32]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_112\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[32]\);
    
    AE_0_sqmuxa_88 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[22]\, Y => 
        \AE_0_sqmuxa_88\);
    
    \PDLCFG_DT_m_27[0]\ : AND3
      port map(A => PDLCFG_DT_3(0), B => \un3_ae[13]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_27_i[0]\);
    
    \P0_50_iv[12]\ : NAND3FFT
      port map(A => \PDLCFG_DT_m_26_i[0]\, B => \P0_m_i[12]\, C
         => \REG_m_i_2[129]\, Y => \P0_50[12]\);
    
    \AE[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_86\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[6]\);
    
    \SBYTE_5[5]\ : MUX2H
      port map(A => \REG[141]\, B => REG_13, S => 
        \sstate_2[6]_net_1\, Y => \SBYTE_5[5]_net_1\);
    
    AE_0_sqmuxa_20 : NAND2
      port map(A => \sstate_8[9]_net_1\, B => \un3_ae[5]\, Y => 
        \AE_0_sqmuxa_20\);
    
    P0_71 : MUX2H
      port map(A => \P0[41]_net_1\, B => \P0_50[41]\, S => 
        \un1_sstate_2_0\, Y => \P0_71\);
    
    \P0[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_37\, CLR => 
        \un1_load_res_8\, Q => \P0[7]_net_1\);
    
    P0_72 : MUX2H
      port map(A => \P0[42]_net_1\, B => \P0_50[42]\, S => 
        \un1_sstate_2_0\, Y => \P0_72\);
    
    CNT_2_I_33 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    AE_0_sqmuxa_176 : NAND2
      port map(A => \sstate_5[9]_net_1\, B => \un3_ae[44]\, Y => 
        \AE_0_sqmuxa_176\);
    
    \P0_50_iv[31]\ : NAND3FTT
      port map(A => \P0_m_i[31]\, B => \PDLCFG_DT_m_15[0]_net_1\, 
        C => \REG_m_i_1[129]\, Y => \P0_50[31]\);
    
    un3_ae_6_1 : NOR2
      port map(A => \CNT[0]_net_1\, B => \CNT[3]_net_1\, Y => 
        \un3_ae_1[6]\);
    
    AE_84 : MUX2H
      port map(A => \AE_PDL_c[4]\, B => \AE_7[4]\, S => 
        \un1_sstate_14\, Y => \AE_84\);
    
    \AE_7_r[40]\ : AND3FFT
      port map(A => \AE_i_m[40]_net_1\, B => \REG_i_m[193]_net_1\, 
        C => N_6864_0, Y => \AE_7[40]\);
    
    un69_ae_23_1 : NOR2FT
      port map(A => REG_0(126), B => REG_0(125), Y => 
        \un69_ae_1[23]\);
    
    \P0_m[21]\ : NAND2
      port map(A => \AE_0_sqmuxa_84\, B => \P0[21]_net_1\, Y => 
        \P0_m[21]_net_1\);
    
    \P_4[1]\ : MUX2H
      port map(A => REG_9, B => PDLCFG_DT(1), S => 
        \sstate[9]_net_1\, Y => \P_4[1]_net_1\);
    
    un3_ae_36 : AND2
      port map(A => \un3_ae_1[39]\, B => \un3_ae_1[44]\, Y => 
        \un3_ae[36]\);
    
    \P0[43]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_73\, CLR => 
        \un1_load_res_8\, Q => \P0[43]_net_1\);
    
    un1_sstate_14 : OR3
      port map(A => \un1_sstate_5\, B => \sstate_0[9]_net_1\, C
         => \sstate[11]_net_1\, Y => \un1_sstate_14\);
    
    AE_88 : MUX2H
      port map(A => \AE_PDL_c[8]\, B => \AE_7[8]\, S => 
        \un1_sstate_14\, Y => \AE_88\);
    
    \AE[43]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_123\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[43]\);
    
    un3_ae_6_2 : OR2
      port map(A => \un3_ae_2[47]\, B => \un3_ae_1[15]\, Y => 
        \un3_ae_2[7]\);
    
    un69_ae_19_1 : NOR2
      port map(A => \un69_ae_1_i[31]\, B => \un69_ae_1[43]\, Y
         => \un69_ae_1[27]\);
    
    AE_121 : MUX2H
      port map(A => \AE_PDL_c[41]\, B => \AE_7[41]\, S => 
        \un1_sstate_14_0\, Y => \AE_121\);
    
    \P0_50_iv[44]\ : NAND3
      port map(A => \PDLCFG_DT_m_4[0]_net_1\, B => 
        \P0_m[44]_net_1\, C => \REG_m_i_0[129]\, Y => \P0_50[44]\);
    
    un1_load_res_6 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_3, Y => 
        \un1_load_res_6\);
    
    \BITCNT_5_r[2]\ : OA21
      port map(A => N_389, B => I_14_1, C => \sstate_0_sqmuxa\, Y
         => \BITCNT_5[2]\);
    
    \PDLCFG_RAD_6[2]\ : MUX2H
      port map(A => \CNT[2]_net_1\, B => PDL_RADDR(2), S => 
        \sstate[6]_net_1\, Y => N_503);
    
    AE_0_sqmuxa_98 : AO21
      port map(A => \un69_ae_1[24]\, B => \un69_ae_2[31]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_98\);
    
    un1_sstate_20 : OAI21
      port map(A => \sstate[3]_net_1\, B => \sstate_1[6]_net_1\, 
        C => \ISI_1_sqmuxa_1\, Y => \un1_sstate_20\);
    
    AE_0_sqmuxa_124 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[31]\, Y => 
        \AE_0_sqmuxa_124\);
    
    \PDLCFG_DT_m_24[0]\ : AND3
      port map(A => PDLCFG_DT_0_0(0), B => \un3_ae[10]\, C => 
        \sstate_7[9]_net_1\, Y => \PDLCFG_DT_m_24_i[0]\);
    
    \PDLCFG_DT_m_44[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[6]\, Y => \PDLCFG_DT_m_44[0]_net_1\);
    
    \P0_50_iv[26]\ : NAND3FTT
      port map(A => \P0_m_i[26]\, B => \PDLCFG_DT_m_10[0]_net_1\, 
        C => \REG_m_i_1[129]\, Y => \P0_50[26]\);
    
    PDLCFG_RAD_27 : MUX2H
      port map(A => \PDLCFG_RAD_6[4]_net_1\, B => 
        \PDLCFG_RAD[4]_net_1\, S => \un1_sstate_25\, Y => 
        \PDLCFG_RAD_27\);
    
    un4_so_5_0_i : INV
      port map(A => N_456_i_i, Y => N_456_i);
    
    AE_125 : MUX2H
      port map(A => \AE_PDL_c[45]\, B => \AE_7[45]\, S => 
        \un1_sstate_14_0\, Y => \AE_125\);
    
    un1_load_res_8 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_2, Y => 
        \un1_load_res_8\);
    
    \P0_m[19]\ : AND2
      port map(A => \AE_0_sqmuxa_76\, B => \P0[19]_net_1\, Y => 
        \P0_m_i[19]\);
    
    un69_ae_21_1 : NOR2
      port map(A => \un69_ae_1_i[31]\, B => \un69_ae_1[45]\, Y
         => \un69_ae_1[29]\);
    
    \P0_50_iv[8]\ : NAND3FTT
      port map(A => \PDLCFG_DT_m_46_i[0]\, B => \P0_m[8]_net_1\, 
        C => \REG_m_i[129]\, Y => \P0_50[8]\);
    
    AE_0_sqmuxa_156 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[39]\, Y => 
        \AE_0_sqmuxa_156\);
    
    \AE[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_96\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[16]\);
    
    un3_ae_19_1 : NOR2
      port map(A => \un3_ae_1_i[31]\, B => \un3_ae_1_i[43]\, Y
         => \un3_ae_1[27]\);
    
    AE_0_sqmuxa_30 : AOI21
      port map(A => \un69_ae_1[7]\, B => \un69_ae_2[7]\, C => 
        \AE_1_sqmuxa\, Y => \AE_0_sqmuxa_30\);
    
    un4_so_12_0 : MUX2H
      port map(A => SP_PDL_in(2), B => SP_PDL_in(34), S => 
        REG_0(127), Y => N_463);
    
    un3_ae_33 : AND2
      port map(A => \un3_ae_1[33]\, B => \un3_ae_1[39]\, Y => 
        \un3_ae[33]\);
    
    \P_4[7]\ : MUX2H
      port map(A => REG_15, B => PDLCFG_DT(7), S => 
        \sstate_8[9]_net_1\, Y => \P_4[7]_net_1\);
    
    un1_sstate_14_1 : OR3
      port map(A => \un1_sstate_5\, B => \sstate_0[9]_net_1\, C
         => \sstate[11]_net_1\, Y => \un1_sstate_14_1\);
    
    \P_4[3]\ : MUX2H
      port map(A => REG_11, B => PDLCFG_DT(3), S => 
        \sstate[9]_net_1\, Y => \P_4[3]_net_1\);
    
    un4_so_9_0 : MUX2H
      port map(A => N_459, B => SP_PDL_in(28), S => REG_0(126), Y
         => N_460);
    
    un3_ae_3 : NOR2
      port map(A => \un3_ae_1[5]\, B => \un3_ae_1_i[43]\, Y => 
        \un3_ae[3]\);
    
    P0_43 : MUX2H
      port map(A => \P0[13]_net_1\, B => \P0_50[13]\, S => 
        \un1_sstate_2_3\, Y => \P0_43\);
    
    AE_101 : MUX2H
      port map(A => \AE_PDL_c[21]\, B => \AE_7[21]\, S => 
        \un1_sstate_14_2\, Y => \AE_101\);
    
    \P0_m[29]\ : NAND2FT
      port map(A => \AE_0_sqmuxa_116\, B => \P0[29]_net_1\, Y => 
        \P0_m[29]_net_1\);
    
    un4_so_33_0_i : INV
      port map(A => N_484_i_i, Y => N_484_i);
    
    \PDLCFG_DT_m_5[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[45]\, Y => \PDLCFG_DT_m_5[0]_net_1\);
    
    \AE_7_r_i_1[47]\ : NOR2
      port map(A => \sstate[12]_net_1\, B => \sstate[11]_net_1\, 
        Y => N_6864_1);
    
    P0_53 : MUX2H
      port map(A => \P0[23]_net_1\, B => \P0_50[23]\, S => 
        \un1_sstate_2_2\, Y => \P0_53\);
    
    \P0_m[42]\ : AND2FT
      port map(A => \AE_0_sqmuxa_168\, B => \P0[42]_net_1\, Y => 
        \P0_m_i[42]\);
    
    \P0_50_iv[19]\ : NAND3FFT
      port map(A => \P0_m_i[19]\, B => \PDLCFG_DT_m_33_i[0]\, C
         => \REG_m_i_2[129]\, Y => \P0_50[19]\);
    
    AE_0_sqmuxa_142 : AOI21
      port map(A => \un69_ae_1[39]\, B => \un69_ae_2[43]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_142\);
    
    \P0_50_iv[41]\ : NAND3FTT
      port map(A => \P0_m_i[41]\, B => \PDLCFG_DT_m_1[0]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[41]\);
    
    un4_so_10_0 : MUX2H
      port map(A => N_455, B => N_460, S => REG_0(124), Y => 
        N_461_i_i);
    
    \P0_50_iv[9]\ : NAND3FTT
      port map(A => \P0_m_i[9]\, B => \PDLCFG_DT_m_23[0]_net_1\, 
        C => \REG_m_i[129]\, Y => \P0_50[9]\);
    
    \P0[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_56\, CLR => 
        \un1_load_res_6\, Q => \P0[26]_net_1\);
    
    \AE_i_m[16]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_64\, B => \AE_0_sqmuxa_66\, C
         => \AE_PDL_c[16]\, Y => \AE_i_m[16]_net_1\);
    
    AE_105 : MUX2H
      port map(A => \AE_PDL_c[25]\, B => \AE_7[25]\, S => 
        \un1_sstate_14_1\, Y => \AE_105\);
    
    P0_63 : MUX2H
      port map(A => \P0[33]_net_1\, B => \P0_50[33]\, S => 
        \un1_sstate_2_1\, Y => \P0_63\);
    
    un4_so_33_0 : MUX2H
      port map(A => N_478, B => N_483, S => REG_5, Y => N_484_i_i);
    
    \P0[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_46\, CLR => 
        \un1_load_res_5\, Q => \P0[16]_net_1\);
    
    \AE_7_r[22]\ : AND3FFT
      port map(A => \AE_i_m[22]_net_1\, B => \REG_i_m[175]_net_1\, 
        C => N_6864_2, Y => \AE_7[22]\);
    
    \REG_m_46_1[129]\ : NAND2
      port map(A => \sstate_0[6]_net_1\, B => REG_8, Y => 
        \REG_m_i_1[129]\);
    
    \PDLCFG_RAD_6_r[3]\ : AND2
      port map(A => N_504, B => \PDLCFG_RAD_1_sqmuxa\, Y => 
        \PDLCFG_RAD_6[3]_net_1\);
    
    \P[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \P_10\, CLR => 
        \un1_load_res_10\, Q => \P_PDL_c[4]\);
    
    \P0_50_iv[38]\ : NAND3FFT
      port map(A => \P0_m_i[38]\, B => \PDLCFG_DT_m_22_i[0]\, C
         => \REG_m_i_0[129]\, Y => \P0_50[38]\);
    
    \AE[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_88\, CLR => 
        \un1_load_res_3\, Q => \AE_PDL_c[8]\);
    
    un1_load_res_9 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_2, Y => 
        \un1_load_res_9\);
    
    \AE_7_r[46]\ : AND3FFT
      port map(A => \AE_i_m[46]_net_1\, B => \REG_i_m[199]_net_1\, 
        C => N_6864_0, Y => \AE_7[46]\);
    
    \AE[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_111\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[31]\);
    
    un3_ae_34 : AND2
      port map(A => \un3_ae_1[39]\, B => \un3_ae_1[42]\, Y => 
        \un3_ae[34]\);
    
    \AE[39]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_119\, CLR => 
        \un1_load_res_2\, Q => \AE_PDL_c[39]\);
    
    \PDL_RDATA[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_21\, CLR => 
        \un1_load_res_10\, Q => \PDL_RDATA[7]_net_1\);
    
    un4_so_18_0 : MUX2H
      port map(A => N_468, B => SP_PDL_in(22), S => REG_5, Y => 
        N_469);
    
    un1_reg_1 : MUX2H
      port map(A => LOAD_RES, B => REG_i_0(121), S => HWRES_c_2, 
        Y => un1_reg_1_i_i);
    
    PDLCFG_RAD_1_sqmuxa_1 : NOR2FT
      port map(A => \sstate[11]_net_1\, B => \un1_cnt\, Y => 
        \sstate_19_1[10]\);
    
    \P0_m[34]\ : AND2
      port map(A => \AE_0_sqmuxa_136\, B => \P0[34]_net_1\, Y => 
        \P0_m_i[34]\);
    
    un3_ae_17_1 : NOR2
      port map(A => \un3_ae_1_i[31]\, B => \un3_ae_1[41]\, Y => 
        \un3_ae_1[25]\);
    
    CNT_2_I_26 : XOR2
      port map(A => \CNT[5]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => \CNT_2[5]\);
    
    \SBYTE_5[6]\ : MUX2H
      port map(A => \REG[142]\, B => REG_14, S => 
        \sstate_2[6]_net_1\, Y => \SBYTE_5[6]_net_1\);
    
    un3_ae_12 : NOR3
      port map(A => \un3_ae_1[45]\, B => \un3_ae_1[14]\, C => 
        \un3_ae_1[15]\, Y => \un3_ae[12]\);
    
    \AE[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_97\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[17]\);
    
    \REG_m[136]\ : AND2
      port map(A => \sstate_2[6]_net_1\, B => REG_15, Y => 
        \REG_m_i[136]\);
    
    \P0_50_iv[33]\ : NAND3FFT
      port map(A => \P0_m_i[33]\, B => \PDLCFG_DT_m_17_i[0]\, C
         => \REG_m_i_1[129]\, Y => \P0_50[33]\);
    
    \AE_i_m[7]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_28\, B => \AE_0_sqmuxa_30\, C
         => \AE_PDL_c[7]\, Y => \AE_i_m[7]_net_1\);
    
    AE_0_sqmuxa_134 : AOI21
      port map(A => \un69_ae_1[33]\, B => \un69_ae_1[39]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_134\);
    
    AE_0_sqmuxa_118 : AO21
      port map(A => \un69_ae_1[29]\, B => \un69_ae_2[31]\, C => 
        \AE_1_sqmuxa_2\, Y => \AE_0_sqmuxa_118\);
    
    \AE[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_106\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[26]\);
    
    un4_so_14_0 : MUX2H
      port map(A => SP_PDL_in(10), B => SP_PDL_in(42), S => REG_6, 
        Y => N_465);
    
    \AE_i_m[24]\ : AOI21
      port map(A => \AE_0_sqmuxa_96\, B => \AE_0_sqmuxa_98\, C
         => \AE_PDL_c[24]\, Y => \AE_i_m[24]_net_1\);
    
    \PDLCFG_DT_m_1[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[41]\, Y => \PDLCFG_DT_m_1[0]_net_1\);
    
    un4_so_8_0 : MUX2H
      port map(A => SP_PDL_in(12), B => SP_PDL_in(44), S => 
        REG_0(127), Y => N_459);
    
    \P0_m[46]\ : AND2FT
      port map(A => \AE_0_sqmuxa_184\, B => \P0[46]_net_1\, Y => 
        \P0_m_i[46]\);
    
    \AE_7_r[33]\ : AND3FFT
      port map(A => \AE_i_m[33]_net_1\, B => \REG_i_m[186]_net_1\, 
        C => N_6864_1, Y => \AE_7[33]\);
    
    \CNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_2[1]\, CLR => 
        \un1_load_res_4\, Q => \CNT[1]_net_1\);
    
    un69_ae_20_1 : NOR2
      port map(A => \un69_ae_1_i[30]\, B => \un69_ae_1[45]\, Y
         => \un69_ae_1[28]\);
    
    CNT_2_I_1 : AND2
      port map(A => \CNT[0]_net_1\, B => \sstate[9]_net_1\, Y => 
        \DWACT_ADD_CI_0_TMP_0[0]\);
    
    \P0_m[8]\ : NAND2
      port map(A => \AE_0_sqmuxa_32\, B => \P0[8]_net_1\, Y => 
        \P0_m[8]_net_1\);
    
    \SBYTE_5[2]\ : MUX2H
      port map(A => \REG[138]\, B => REG_10, S => 
        \sstate_2[6]_net_1\, Y => \SBYTE_5[2]_net_1\);
    
    AE_0_sqmuxa_146 : AOI21
      port map(A => \un69_ae_1[39]\, B => \un69_ae_1[44]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_146\);
    
    un69_ae_18_1 : NOR2
      port map(A => \un69_ae_1_i[30]\, B => \un69_ae_1[43]\, Y
         => \un69_ae_1[26]\);
    
    un3_ae_10 : NOR2FT
      port map(A => \un3_ae_1[11]\, B => \un3_ae_1[14]\, Y => 
        \un3_ae[10]\);
    
    \P0_50_iv[0]\ : NAND3FFT
      port map(A => \PDLCFG_DT_m_38_i[0]\, B => \P0_m_i[0]\, C
         => \REG_m_i[129]\, Y => \P0_50[0]\);
    
    un4_so_39_0 : MUX2H
      port map(A => N_487, B => N_492, S => REG_3, Y => N_490_i_i);
    
    AE_0_sqmuxa_168 : NAND2
      port map(A => \sstate_5[9]_net_1\, B => \un3_ae[42]\, Y => 
        \AE_0_sqmuxa_168\);
    
    un69_ae_35_1 : NOR2
      port map(A => \un69_ae_1[43]\, B => \un69_ae_1_i[47]\, Y
         => \un69_ae_2[43]\);
    
    un4_so_27_0 : MUX2H
      port map(A => N_477, B => N_482, S => REG_3, Y => N_478);
    
    AE_122 : MUX2H
      port map(A => \AE_PDL_c[42]\, B => \AE_7[42]\, S => 
        \un1_sstate_14_0\, Y => \AE_122\);
    
    \P0[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_57\, CLR => 
        \un1_load_res_6\, Q => \P0[27]_net_1\);
    
    un4_so_36_0 : MUX2H
      port map(A => N_486, B => SP_PDL_in(19), S => REG_5, Y => 
        N_487);
    
    \P0[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_47\, CLR => 
        \un1_load_res_5\, Q => \P0[17]_net_1\);
    
    ISI_0_sqmuxa : NAND2
      port map(A => \sstate[1]_net_1\, B => \un5_bitcnt\, Y => 
        \ISI_0_sqmuxa\);
    
    AE_0_sqmuxa_1 : NAND2
      port map(A => \sstate_1[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        AE_0_sqmuxa_i_1);
    
    P_10 : MUX2H
      port map(A => \P_PDL_c[4]\, B => \P_4[4]_net_1\, S => 
        \un1_sstate_2\, Y => \P_10\);
    
    \P0_50_iv[35]\ : NAND3FFT
      port map(A => \P0_m_i[35]\, B => \PDLCFG_DT_m_19_i[0]\, C
         => \REG_m_i_1[129]\, Y => \P0_50[35]\);
    
    ISI_78 : MUX2H
      port map(A => ISI_5, B => \SI_PDL_c\, S => \un1_sstate_18\, 
        Y => \ISI_78\);
    
    MODE_0 : MUX2H
      port map(A => \MD_PDL_c_0\, B => \MODE_2\, S => 
        \un1_sstate_5\, Y => \MODE_0\);
    
    un3_ae_47_2 : NAND2
      port map(A => \CNT[1]_net_1\, B => \CNT[2]_net_1\, Y => 
        \un3_ae_2[47]\);
    
    \P0_m[33]\ : AND2
      port map(A => \AE_0_sqmuxa_132\, B => \P0[33]_net_1\, Y => 
        \P0_m_i[33]\);
    
    \AE[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_93\, CLR => 
        \un1_load_res_0\, Q => \AE_PDL_c[13]\);
    
    \AE_i_m[44]\ : AOI21
      port map(A => \AE_0_sqmuxa_176\, B => \AE_0_sqmuxa_178\, C
         => \AE_PDL_c[44]\, Y => \AE_i_m[44]_net_1\);
    
    un4_so_21_0 : MUX2H
      port map(A => N_466, B => N_471, S => REG_0(124), Y => 
        N_472_i_i);
    
    un3_ae_18_1 : NOR2
      port map(A => \un3_ae_1[30]\, B => \un3_ae_1_i[43]\, Y => 
        \un3_ae_1[26]\);
    
    un1_sstate_18 : OAI21
      port map(A => \sstate[12]_net_1\, B => \un1_sstate_1\, C
         => \ISI_0_sqmuxa\, Y => \un1_sstate_18\);
    
    AE_0_sqmuxa_2 : OA21FTF
      port map(A => \un69_ae_0_0\, B => \un69_ae_1[15]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_2\);
    
    \SBYTE[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_129\, CLR => 
        \un1_load_res_10\, Q => \REG[137]\);
    
    \P0_m[15]\ : NAND2
      port map(A => \AE_0_sqmuxa_60\, B => \P0[15]_net_1\, Y => 
        \P0_m[15]_net_1\);
    
    \P0_50_iv[16]\ : NAND3FFT
      port map(A => \PDLCFG_DT_m_30_i[0]\, B => \P0_m_i[16]\, C
         => \REG_m_i_2[129]\, Y => \P0_50[16]\);
    
    AE_96 : MUX2H
      port map(A => \AE_PDL_c[16]\, B => \AE_7[16]\, S => 
        \un1_sstate_14_2\, Y => \AE_96\);
    
    AE_99 : MUX2H
      port map(A => \AE_PDL_c[19]\, B => \AE_7[19]\, S => 
        \un1_sstate_14_2\, Y => \AE_99\);
    
    AE_102 : MUX2H
      port map(A => \AE_PDL_c[22]\, B => \AE_7[22]\, S => 
        \un1_sstate_14_2\, Y => \AE_102\);
    
    P_12 : MUX2H
      port map(A => \P_PDL_c[6]\, B => \P_4[6]_net_1\, S => 
        \un1_sstate_2\, Y => \P_12\);
    
    AE_0_sqmuxa_2_0 : NAND2
      port map(A => \sstate_0[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        AE_0_sqmuxa_i_2);
    
    un69_ae_6_0_1 : NOR2
      port map(A => REG_1, B => REG_4, Y => \un69_ae_1[6]\);
    
    \AE[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_107\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[27]\);
    
    un1_load_res_4 : OR2FT
      port map(A => LOAD_RES_3, B => HWRES_c_0_3, Y => 
        \un1_load_res_4\);
    
    \P0_50_iv[43]\ : NAND3FTT
      port map(A => \P0_m_i[43]\, B => \PDLCFG_DT_m_3[0]_net_1\, 
        C => \REG_m_i_0[129]\, Y => \P0_50[43]\);
    
    \AE_i_m[17]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_68\, B => \AE_0_sqmuxa_70\, C
         => \AE_PDL_c[17]\, Y => \AE_i_m[17]_net_1\);
    
    \P0_m[30]\ : AND2FT
      port map(A => \AE_0_sqmuxa_120\, B => \P0[30]_net_1\, Y => 
        \P0_m_i[30]\);
    
    \AE_7_r[39]\ : AND3FFT
      port map(A => \AE_i_m[39]_net_1\, B => \REG_i_m[192]_net_1\, 
        C => N_6864_0, Y => \AE_7[39]\);
    
    AE_0_sqmuxa_54 : OA21FTF
      port map(A => \un69_ae_13_0\, B => \un69_ae_1[15]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_54\);
    
    AE_0_sqmuxa_44 : NAND2
      port map(A => \sstate_7[9]_net_1\, B => \un3_ae[11]\, Y => 
        \AE_0_sqmuxa_44\);
    
    \CNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_2[2]\, CLR => 
        \un1_load_res_4\, Q => \CNT[2]_net_1\);
    
    un3_ae_27 : NAND2
      port map(A => \un3_ae_1[27]\, B => \un3_ae_2[31]\, Y => 
        \un3_ae[27]\);
    
    CNT_2_I_34 : AND2
      port map(A => \CNT[2]_net_1\, B => \CNT[3]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    AE_0_sqmuxa : NAND2
      port map(A => \sstate_2[6]_net_1\, B => \MD_PDL_c_0\, Y => 
        AE_0_sqmuxa_i);
    
    \REG_i_m[198]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_77, Y => 
        \REG_i_m[198]_net_1\);
    
    \P0[42]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_72\, CLR => 
        \un1_load_res_7\, Q => \P0[42]_net_1\);
    
    \AE_7_r[28]\ : AND3FFT
      port map(A => \AE_i_m[28]_net_1\, B => \REG_i_m[181]_net_1\, 
        C => N_6864_1, Y => \AE_7[28]\);
    
    \AE_i_m[15]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_60\, B => \AE_0_sqmuxa_62\, C
         => \AE_PDL_c[15]\, Y => \AE_i_m[15]_net_1\);
    
    un3_ae_47 : NAND2
      port map(A => \un3_ae_3[47]\, B => \un3_ae_4[47]\, Y => 
        \un3_ae[47]\);
    
    \AE_7_r[47]\ : AND3FFT
      port map(A => \AE_i_m[47]_net_1\, B => \REG_i_m[200]_net_1\, 
        C => N_6864_0, Y => \AE_7[47]\);
    
    un3_ae_11 : OR2FT
      port map(A => \un3_ae_1[11]\, B => \un3_ae_2[15]\, Y => 
        \un3_ae[11]\);
    
    \sstate[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_19_1[10]\, CLR => 
        \un1_load_res_11\, Q => \sstate[10]_net_1\);
    
    \P0_m[25]\ : AND2FT
      port map(A => \AE_0_sqmuxa_100\, B => \P0[25]_net_1\, Y => 
        \P0_m_i[25]\);
    
    \AE_7_r[30]\ : AND3FFT
      port map(A => \AE_i_m[30]_net_1\, B => \REG_i_m[183]_net_1\, 
        C => N_6864_1, Y => \AE_7[30]\);
    
    AE_0_sqmuxa_128 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[32]\, Y => 
        \AE_0_sqmuxa_128\);
    
    un1_sstate_27 : OR3
      port map(A => \PDLCFG_RAD_0_sqmuxa_1\, B => 
        un1_sstate_27_2_i, C => un1_sstate_27_3_i, Y => 
        \un1_sstate_27\);
    
    \P0_m[4]\ : NAND2
      port map(A => \AE_0_sqmuxa_16\, B => \P0[4]_net_1\, Y => 
        \P0_m[4]_net_1\);
    
    un1_sstate_2 : OR2
      port map(A => \sstate_0[9]_net_1\, B => \sstate_1[6]_net_1\, 
        Y => \un1_sstate_2\);
    
    \AE_7_r[45]\ : AND3FFT
      port map(A => \AE_i_m[45]_net_1\, B => \REG_i_m[198]_net_1\, 
        C => N_6864_0, Y => \AE_7[45]\);
    
    \REG_i_m[181]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_60, Y => 
        \REG_i_m[181]_net_1\);
    
    un3_ae_8 : NOR2FT
      port map(A => \un3_ae_1[9]\, B => \un3_ae_1[14]\, Y => 
        \un3_ae[8]\);
    
    un3_ae_15 : NOR2
      port map(A => \un3_ae_2[7]\, B => \un3_ae_2[15]\, Y => 
        \un3_ae[15]\);
    
    \PDLCFG_DT_m_23[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_1(0), C
         => \un3_ae[9]\, Y => \PDLCFG_DT_m_23[0]_net_1\);
    
    \PDLCFG_DT_m_43[0]\ : OR3FFT
      port map(A => \sstate_4[9]_net_1\, B => PDLCFG_DT_2(0), C
         => \un3_ae[5]\, Y => \PDLCFG_DT_m_43[0]_net_1\);
    
    \PDLCFG_DT_m_4[0]\ : OR3FFT
      port map(A => \sstate_3[9]_net_1\, B => PDLCFG_DT_0(0), C
         => \un3_ae[44]\, Y => \PDLCFG_DT_m_4[0]_net_1\);
    
    \P0[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_31\, CLR => 
        \un1_load_res_5\, Q => \P0[1]_net_1\);
    
    \P0_50_iv[45]\ : NAND3
      port map(A => \PDLCFG_DT_m_5[0]_net_1\, B => 
        \P0_m[45]_net_1\, C => \REG_m_i_0[129]\, Y => \P0_50[45]\);
    
    un3_ae_23_1 : OR2FT
      port map(A => \CNT[4]_net_1\, B => \CNT[3]_net_1\, Y => 
        \un3_ae_1[23]\);
    
    \SBYTE[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_130\, CLR => 
        \un1_load_res_10\, Q => \REG[138]\);
    
    PDLCFG_RAD_0_sqmuxa_1 : AND2
      port map(A => \sstate[11]_net_1\, B => \un1_cnt\, Y => 
        \PDLCFG_RAD_0_sqmuxa_1\);
    
    \REG_i_m[196]\ : NOR2
      port map(A => AE_0_sqmuxa_i_0, B => REG_75, Y => 
        \REG_i_m[196]_net_1\);
    
    un4_so_4_0 : MUX2H
      port map(A => N_454, B => SP_PDL_in(24), S => REG_0(126), Y
         => N_455);
    
    \AE_i_m[6]\ : AOI21
      port map(A => \AE_0_sqmuxa_24\, B => \AE_0_sqmuxa_26\, C
         => \AE_PDL_c[6]\, Y => \AE_i_m[6]_net_1\);
    
    \AE[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \AE_103\, CLR => 
        \un1_load_res_1\, Q => \AE_PDL_c[23]\);
    
    AE_0_sqmuxa_174 : AO21
      port map(A => \un69_ae_2[43]\, B => \un69_ae_3[47]\, C => 
        \AE_1_sqmuxa_0\, Y => \AE_0_sqmuxa_174\);
    
    un4_so_22_0 : MUX2H
      port map(A => N_467_i, B => N_472_i, S => REG_4, Y => N_473);
    
    \P0[33]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_63\, CLR => 
        \un1_load_res_7\, Q => \P0[33]_net_1\);
    
    AE_0_sqmuxa_68 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[17]\, Y => 
        \AE_0_sqmuxa_68\);
    
    \AE_i_m[32]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_128\, B => \AE_0_sqmuxa_130\, C
         => \AE_PDL_c[32]\, Y => \AE_i_m[32]_net_1\);
    
    AE_0_sqmuxa_100 : NAND2
      port map(A => \sstate_6[9]_net_1\, B => \un3_ae[25]\, Y => 
        \AE_0_sqmuxa_100\);
    
    \AE_7_r[12]\ : AND3FFT
      port map(A => \AE_i_m[12]_net_1\, B => \REG_i_m[165]_net_1\, 
        C => N_6864_2, Y => \AE_7[12]\);
    
    un3_ae_31_1 : OR2FT
      port map(A => \CNT[0]_net_1\, B => \CNT[5]_net_1\, Y => 
        \un3_ae_1_i[31]\);
    
    \SBYTE[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_132\, CLR => 
        \un1_load_res_11\, Q => \REG[140]\);
    
    AE_0_sqmuxa_80 : NOR2FT
      port map(A => \sstate_2[9]_net_1\, B => \un3_ae[20]\, Y => 
        \AE_0_sqmuxa_80\);
    
    un4_so_47_0 : MUX2H
      port map(A => N_474, B => N_497, S => REG_1, Y => un4_so);
    
    \P0[38]\ : DFFC
      port map(CLK => CLK_c_c, D => \P0_68\, CLR => 
        \un1_load_res_7\, Q => \P0[38]_net_1\);
    
    un4_so_20_0 : MUX2H
      port map(A => N_470, B => SP_PDL_in(30), S => REG_5, Y => 
        N_471);
    
    \P_4[2]\ : MUX2H
      port map(A => REG_10, B => PDLCFG_DT(2), S => 
        \sstate[9]_net_1\, Y => \P_4[2]_net_1\);
    
    P0_48 : MUX2H
      port map(A => \P0[18]_net_1\, B => \P0_50[18]\, S => 
        \un1_sstate_2_2\, Y => \P0_48\);
    
    \sstate[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_19[5]\, CLR => 
        \un1_load_res\, Q => \sstate[5]_net_1\);
    
    \REG_i_m[168]\ : NOR2
      port map(A => AE_0_sqmuxa_i_2, B => REG_47, Y => 
        \REG_i_m[168]_net_1\);
    
    un69_ae_10_1 : NOR2
      port map(A => \un69_ae_1[15]\, B => \un69_ae_1[43]\, Y => 
        \un69_ae_1[11]\);
    
    \PDL_RDATA[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RDATA_14\, CLR => 
        \un1_load_res_9\, Q => \PDL_RDATA[0]_net_1\);
    
    \BITCNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_5[0]\, CLR => 
        \un1_load_res_4\, Q => \BITCNT[0]_net_1\);
    
    AE_0_sqmuxa_76 : NOR2FT
      port map(A => \sstate_1[9]_net_1\, B => \un3_ae[19]\, Y => 
        \AE_0_sqmuxa_76\);
    
    P0_58 : MUX2H
      port map(A => \P0[28]_net_1\, B => \P0_50[28]\, S => 
        \un1_sstate_2_1\, Y => \P0_58\);
    
    \PDLCFG_RAD_6[4]\ : MUX2H
      port map(A => \CNT[4]_net_1\, B => PDL_RADDR(4), S => 
        \sstate[6]_net_1\, Y => N_505);
    
    \REG_i_m[178]\ : NOR2
      port map(A => AE_0_sqmuxa_i_1, B => REG_57, Y => 
        \REG_i_m[178]_net_1\);
    
    \P0_m[37]\ : NAND2
      port map(A => \AE_0_sqmuxa_148\, B => \P0[37]_net_1\, Y => 
        \P0_m[37]_net_1\);
    
    \BITCNT_5_r[1]\ : OA21
      port map(A => N_389, B => I_13_5, C => \sstate_0_sqmuxa\, Y
         => \BITCNT_5[1]\);
    
    \AE_i_m[21]\ : OA21TTF
      port map(A => \AE_0_sqmuxa_84\, B => \AE_0_sqmuxa_86\, C
         => \AE_PDL_c[21]\, Y => \AE_i_m[21]_net_1\);
    
    P0_68 : MUX2H
      port map(A => \P0[38]_net_1\, B => \P0_50[38]\, S => 
        \un1_sstate_2_0\, Y => \P0_68\);
    
    AE_0_sqmuxa_154 : AOI21
      port map(A => \un69_ae_1[38]\, B => \un69_ae_1[39]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_154\);
    
    un4_so_28_0 : MUX2H
      port map(A => N_476, B => N_481, S => REG_3, Y => N_479_i_i);
    
    un4_so_41_0 : MUX2H
      port map(A => N_491, B => SP_PDL_in(23), S => REG_5, Y => 
        N_492);
    
    un3_ae_7_1 : NOR2FT
      port map(A => \CNT[0]_net_1\, B => \CNT[3]_net_1\, Y => 
        \un3_ae_1[7]\);
    
    \PDLCFG_DT_m_22[0]\ : AND3
      port map(A => PDLCFG_DT_2(0), B => \un3_ae[38]\, C => 
        \sstate_5[9]_net_1\, Y => \PDLCFG_DT_m_22_i[0]\);
    
    AE_0_sqmuxa_138 : AOI21
      port map(A => \un69_ae_1[39]\, B => \un69_ae_1[42]\, C => 
        \AE_1_sqmuxa_1\, Y => \AE_0_sqmuxa_138\);
    
    \PDLCFG_RAD[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDLCFG_RAD_23\, CLR => 
        \un1_load_res_8\, Q => \PDLCFG_RAD[0]_net_1\);
    
    \PDLCFG_DT_m_42[0]\ : AND3
      port map(A => PDLCFG_DT(0), B => \un3_ae[4]\, C => 
        \sstate_8[9]_net_1\, Y => \PDLCFG_DT_m_42_i[0]\);
    
    \AE_7_r[36]\ : AND3FFT
      port map(A => \AE_i_m[36]_net_1\, B => \REG_i_m[189]_net_1\, 
        C => N_6864_0, Y => \AE_7[36]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity PDLCFG is

    port( CROMWDT       : in    std_logic_vector(7 downto 0);
          PDLCFG_RAD    : in    std_logic_vector(5 downto 0);
          CROMWAD       : in    std_logic_vector(5 downto 0);
          PDLCFG_DT_0   : out   std_logic_vector(0 to 0);
          PDLCFG_DT_1   : out   std_logic_vector(0 to 0);
          PDLCFG_DT_2   : out   std_logic_vector(0 to 0);
          PDLCFG_DT_3   : out   std_logic_vector(0 to 0);
          PDLCFG_DT     : out   std_logic_vector(7 downto 0);
          PDLCFG_DT_0_0 : out   std_logic_vector(0 to 0);
          PDLCFG_nRD    : in    std_logic;
          PDLCFG_nWR    : in    std_logic;
          CLK_c_c       : in    std_logic
        );

end PDLCFG;

architecture DEF_ARCH of PDLCFG is 

  component BFR
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component RAM256x9SSTP
    generic (MEMORYFILE:string := "");

    port( DO8    : out   std_logic;
          DO7    : out   std_logic;
          DO6    : out   std_logic;
          DO5    : out   std_logic;
          DO4    : out   std_logic;
          DO3    : out   std_logic;
          DO2    : out   std_logic;
          DO1    : out   std_logic;
          DO0    : out   std_logic;
          DOS    : out   std_logic;
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          DI8    : in    std_logic := 'U';
          DI7    : in    std_logic := 'U';
          DI6    : in    std_logic := 'U';
          DI5    : in    std_logic := 'U';
          DI4    : in    std_logic := 'U';
          DI3    : in    std_logic := 'U';
          DI2    : in    std_logic := 'U';
          DI1    : in    std_logic := 'U';
          DI0    : in    std_logic := 'U';
          WRB    : in    std_logic := 'U';
          RDB    : in    std_logic := 'U';
          WBLKB  : in    std_logic := 'U';
          RBLKB  : in    std_logic := 'U';
          PARODD : in    std_logic := 'U';
          WCLKS  : in    std_logic := 'U';
          RCLKS  : in    std_logic := 'U';
          DIS    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \PDLCFG_DT_0_0[0]\, M0_DO8, \PDLCFG_DT[0]\, net00011, 
        \GND\, \VCC\ : std_logic;

begin 

    PDLCFG_DT(0) <= \PDLCFG_DT[0]\;
    PDLCFG_DT_0_0(0) <= \PDLCFG_DT_0_0[0]\;

    M0_2 : BFR
      port map(A => \PDLCFG_DT_0_0[0]\, Y => PDLCFG_DT_2(0));
    
    M0_1 : BFR
      port map(A => \PDLCFG_DT_0_0[0]\, Y => PDLCFG_DT_1(0));
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    M0 : RAM256x9SSTP
      generic map(MEMORYFILE => "PDLCFG_M0.mem")

      port map(DO8 => M0_DO8, DO7 => PDLCFG_DT(7), DO6 => 
        PDLCFG_DT(6), DO5 => PDLCFG_DT(5), DO4 => PDLCFG_DT(4), 
        DO3 => PDLCFG_DT(3), DO2 => PDLCFG_DT(2), DO1 => 
        PDLCFG_DT(1), DO0 => \PDLCFG_DT[0]\, DOS => net00011, 
        WADDR7 => \GND\, WADDR6 => \GND\, WADDR5 => CROMWAD(5), 
        WADDR4 => CROMWAD(4), WADDR3 => CROMWAD(3), WADDR2 => 
        CROMWAD(2), WADDR1 => CROMWAD(1), WADDR0 => CROMWAD(0), 
        RADDR7 => \GND\, RADDR6 => \GND\, RADDR5 => PDLCFG_RAD(5), 
        RADDR4 => PDLCFG_RAD(4), RADDR3 => PDLCFG_RAD(3), RADDR2
         => PDLCFG_RAD(2), RADDR1 => PDLCFG_RAD(1), RADDR0 => 
        PDLCFG_RAD(0), DI8 => \GND\, DI7 => CROMWDT(7), DI6 => 
        CROMWDT(6), DI5 => CROMWDT(5), DI4 => CROMWDT(4), DI3 => 
        CROMWDT(3), DI2 => CROMWDT(2), DI1 => CROMWDT(1), DI0 => 
        CROMWDT(0), WRB => PDLCFG_nWR, RDB => PDLCFG_nRD, WBLKB
         => \GND\, RBLKB => \GND\, PARODD => \GND\, WCLKS => 
        CLK_c_c, RCLKS => CLK_c_c, DIS => \GND\);
    
    M0_0 : BFR
      port map(A => \PDLCFG_DT_0_0[0]\, Y => PDLCFG_DT_0(0));
    
    M0_0_0 : BFR
      port map(A => \PDLCFG_DT[0]\, Y => \PDLCFG_DT_0_0[0]\);
    
    M0_3 : BFR
      port map(A => \PDLCFG_DT_0_0[0]\, Y => PDLCFG_DT_3(0));
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity VINTERF is

    port( TICK            : in    std_logic_vector(2 to 2);
          RAMDT           : in    std_logic_vector(7 downto 0);
          VADm            : out   std_logic_vector(31 downto 0);
          RAMAD_VME       : out   std_logic_vector(8 downto 0);
          AMB_c           : in    std_logic_vector(5 downto 0);
          LB_in           : in    std_logic_vector(31 downto 0);
          OR_RDATA        : out   std_logic_vector(9 downto 0);
          PULSE_0         : out   std_logic;
          PULSE_1         : out   std_logic;
          PULSE_2         : out   std_logic;
          PULSE_3         : out   std_logic;
          PULSE_6         : out   std_logic;
          PULSE_7         : out   std_logic;
          PULSE_8         : out   std_logic;
          PULSE_9         : out   std_logic;
          PULSE_10        : out   std_logic;
          OR_RADDR        : in    std_logic_vector(5 downto 0);
          VDB_in_0        : in    std_logic_vector(15 downto 0);
          VDB_in          : in    std_logic_vector(31 downto 0);
          LB_i            : out   std_logic_vector(31 downto 0);
          DPR             : in    std_logic_vector(31 downto 0);
          FBOUT           : in    std_logic_vector(7 downto 0);
          LBSP_c          : in    std_logic_vector(2 to 2);
          REGMAP_35       : out   std_logic;
          REGMAP_31       : out   std_logic;
          REG_c_21        : in    std_logic;
          REG_c_22        : in    std_logic;
          REG_c_23        : in    std_logic;
          REG_c_0         : out   std_logic;
          LBSP_in_0       : in    std_logic;
          LBSP_in_1       : in    std_logic;
          LBSP_in_15      : in    std_logic;
          LBSP_in_16      : in    std_logic;
          LBSP_in_17      : in    std_logic;
          LBSP_in_18      : in    std_logic;
          LBSP_in_19      : in    std_logic;
          LBSP_in_20      : in    std_logic;
          LBSP_in_21      : in    std_logic;
          LBSP_in_22      : in    std_logic;
          LBSP_in_23      : in    std_logic;
          LBSP_in_24      : in    std_logic;
          LBSP_in_25      : in    std_logic;
          LBSP_in_26      : in    std_logic;
          LBSP_in_27      : in    std_logic;
          LBSP_in_28      : in    std_logic;
          LBSP_in_29      : in    std_logic;
          LBSP_in_30      : in    std_logic;
          LBSP_in_31      : in    std_logic;
          VAD_in_0        : in    std_logic;
          VAD_in_1        : in    std_logic;
          VAD_in_2        : in    std_logic;
          VAD_in_3        : in    std_logic;
          VAD_in_4        : in    std_logic;
          VAD_in_5        : in    std_logic;
          VAD_in_6        : in    std_logic;
          VAD_in_7        : in    std_logic;
          VAD_in_8        : in    std_logic;
          VAD_in_9        : in    std_logic;
          VAD_in_10       : in    std_logic;
          VAD_in_11       : in    std_logic;
          VAD_in_12       : in    std_logic;
          VAD_in_13       : in    std_logic;
          VAD_in_14       : in    std_logic;
          VAD_in_27       : in    std_logic;
          VAD_in_28       : in    std_logic;
          VAD_in_29       : in    std_logic;
          VAD_in_30       : in    std_logic;
          GA_c            : in    std_logic_vector(3 downto 0);
          VDBm_0          : out   std_logic;
          VDBm_1          : out   std_logic;
          VDBm_2          : out   std_logic;
          VDBm_3          : out   std_logic;
          VDBm_4          : out   std_logic;
          VDBm_5          : out   std_logic;
          VDBm_6          : out   std_logic;
          VDBm_7          : out   std_logic;
          VDBm_8          : out   std_logic;
          VDBm_9          : out   std_logic;
          VDBm_10         : out   std_logic;
          VDBm_12         : out   std_logic;
          VDBm_13         : out   std_logic;
          VDBm_14         : out   std_logic;
          VDBm_15         : out   std_logic;
          VDBm_16         : out   std_logic;
          VDBm_17         : out   std_logic;
          VDBm_18         : out   std_logic;
          VDBm_19         : out   std_logic;
          VDBm_20         : out   std_logic;
          VDBm_22         : out   std_logic;
          VDBm_23         : out   std_logic;
          VDBm_24         : out   std_logic;
          VDBm_25         : out   std_logic;
          VDBm_26         : out   std_logic;
          VDBm_27         : out   std_logic;
          VDBm_28         : out   std_logic;
          VDBm_29         : out   std_logic;
          VDBm_30         : out   std_logic;
          VDBm_31         : out   std_logic;
          VDBm_i_m2       : out   std_logic_vector(11 to 11);
          REG_126         : out   std_logic;
          REG_125         : out   std_logic;
          REG_124         : out   std_logic;
          REG_123         : out   std_logic;
          REG_344         : out   std_logic;
          REG_345         : out   std_logic;
          REG_359         : out   std_logic;
          REG_360         : out   std_logic;
          REG_361         : out   std_logic;
          REG_362         : out   std_logic;
          REG_363         : out   std_logic;
          REG_364         : out   std_logic;
          REG_365         : out   std_logic;
          REG_366         : out   std_logic;
          REG_367         : out   std_logic;
          REG_368         : out   std_logic;
          REG_369         : out   std_logic;
          REG_370         : out   std_logic;
          REG_371         : out   std_logic;
          REG_372         : out   std_logic;
          REG_373         : out   std_logic;
          REG_374         : out   std_logic;
          REG_375         : out   std_logic;
          REG_408         : out   std_logic;
          REG_480         : out   std_logic;
          REG_80          : out   std_logic;
          REG_81          : out   std_logic;
          REG_82          : out   std_logic;
          REG_83          : out   std_logic;
          REG_84          : out   std_logic;
          REG_85          : out   std_logic;
          REG_86          : out   std_logic;
          REG_87          : out   std_logic;
          REG_88          : out   std_logic;
          REG_89          : out   std_logic;
          REG_90          : out   std_logic;
          REG_96          : out   std_logic;
          REG_97          : out   std_logic;
          REG_98          : out   std_logic;
          REG_99          : out   std_logic;
          REG_100         : out   std_logic;
          REG_101         : out   std_logic;
          REG_102         : out   std_logic;
          REG_103         : out   std_logic;
          REG_376         : out   std_logic;
          REG_120         : out   std_logic;
          REG_152         : out   std_logic;
          REG_232         : out   std_logic;
          REG_248         : out   std_logic;
          REG_168         : out   std_logic;
          REG_184         : out   std_logic;
          REG_104         : in    std_logic;
          REG_136         : in    std_logic;
          REG_31          : in    std_logic;
          REG_47          : out   std_logic;
          REG_440         : out   std_logic;
          REG_456         : in    std_logic;
          REG_441         : out   std_logic;
          REG_457         : in    std_logic;
          REG_473         : in    std_logic;
          REG_121         : out   std_logic;
          REG_153         : out   std_logic;
          REG_233         : out   std_logic;
          REG_249         : out   std_logic;
          REG_169         : out   std_logic;
          REG_185         : out   std_logic;
          REG_105         : in    std_logic;
          REG_137         : in    std_logic;
          REG_32          : in    std_logic;
          REG_16          : in    std_logic;
          REG_48          : out   std_logic;
          REG_377         : out   std_logic;
          REG_409         : out   std_logic;
          REG_442         : out   std_logic;
          REG_458         : in    std_logic;
          REG_474         : in    std_logic;
          REG_378         : out   std_logic;
          REG_410         : out   std_logic;
          REG_154         : out   std_logic;
          REG_170         : out   std_logic;
          REG_122         : out   std_logic;
          REG_250         : out   std_logic;
          REG_138         : in    std_logic;
          REG_186         : out   std_logic;
          REG_234         : out   std_logic;
          REG_33          : in    std_logic;
          REG_49          : out   std_logic;
          REG_34          : in    std_logic;
          REG_50          : out   std_logic;
          REG_155         : out   std_logic;
          REG_171         : out   std_logic;
          REG_251         : out   std_logic;
          REG_139         : in    std_logic;
          REG_187         : out   std_logic;
          REG_235         : out   std_logic;
          REG_443         : out   std_logic;
          REG_459         : in    std_logic;
          REG_379         : out   std_logic;
          REG_411         : out   std_logic;
          REG_475         : in    std_logic;
          REG_51          : out   std_logic;
          REG_35          : in    std_logic;
          REG_19          : in    std_logic;
          REG_156         : out   std_logic;
          REG_172         : out   std_logic;
          REG_252         : out   std_logic;
          REG_140         : in    std_logic;
          REG_188         : out   std_logic;
          REG_236         : out   std_logic;
          REG_332         : in    std_logic;
          REG_444         : out   std_logic;
          REG_460         : in    std_logic;
          REG_380         : out   std_logic;
          REG_412         : out   std_logic;
          REG_476         : in    std_logic;
          REG_445         : out   std_logic;
          REG_461         : in    std_logic;
          REG_413         : out   std_logic;
          REG_381         : out   std_logic;
          REG_52          : out   std_logic;
          REG_36          : in    std_logic;
          REG_157         : out   std_logic;
          REG_173         : out   std_logic;
          REG_253         : out   std_logic;
          REG_141         : in    std_logic;
          REG_189         : out   std_logic;
          REG_237         : out   std_logic;
          REG_333         : in    std_logic;
          REG_477         : in    std_logic;
          REG_462         : in    std_logic;
          REG_478         : in    std_logic;
          REG_382         : out   std_logic;
          REG_414         : out   std_logic;
          REG_37          : in    std_logic;
          REG_5           : out   std_logic;
          REG_53          : out   std_logic;
          REG_158         : out   std_logic;
          REG_174         : out   std_logic;
          REG_254         : out   std_logic;
          REG_142         : in    std_logic;
          REG_190         : out   std_logic;
          REG_238         : out   std_logic;
          REG_334         : in    std_logic;
          REG_463         : in    std_logic;
          REG_383         : out   std_logic;
          REG_415         : out   std_logic;
          REG_54          : out   std_logic;
          REG_38          : in    std_logic;
          REG_159         : out   std_logic;
          REG_175         : out   std_logic;
          REG_255         : out   std_logic;
          REG_143         : in    std_logic;
          REG_191         : out   std_logic;
          REG_239         : out   std_logic;
          REG_479         : in    std_logic;
          REG_464         : in    std_logic;
          REG_416         : out   std_logic;
          REG_39          : in    std_logic;
          REG_7           : out   std_logic;
          REG_55          : out   std_logic;
          REG_128         : out   std_logic;
          REG_160         : out   std_logic;
          REG_240         : out   std_logic;
          REG_256         : out   std_logic;
          REG_176         : out   std_logic;
          REG_192         : out   std_logic;
          REG_112         : in    std_logic;
          REG_144         : in    std_logic;
          REG_465         : in    std_logic;
          REG_56          : out   std_logic;
          REG_40          : in    std_logic;
          REG_161         : out   std_logic;
          REG_177         : out   std_logic;
          REG_129         : out   std_logic;
          REG_257         : out   std_logic;
          REG_113         : in    std_logic;
          REG_193         : out   std_logic;
          REG_241         : out   std_logic;
          REG_417         : out   std_logic;
          REG_466         : in    std_logic;
          REG_57          : out   std_logic;
          REG_41          : in    std_logic;
          REG_162         : out   std_logic;
          REG_178         : out   std_logic;
          REG_130         : out   std_logic;
          REG_258         : out   std_logic;
          REG_114         : in    std_logic;
          REG_194         : out   std_logic;
          REG_242         : out   std_logic;
          REG_418         : out   std_logic;
          REG_467         : in    std_logic;
          REG_42          : in    std_logic;
          REG_58          : out   std_logic;
          REG_163         : out   std_logic;
          REG_179         : out   std_logic;
          REG_131         : out   std_logic;
          REG_259         : out   std_logic;
          REG_115         : in    std_logic;
          REG_195         : out   std_logic;
          REG_243         : out   std_logic;
          REG_419         : out   std_logic;
          REG_468         : in    std_logic;
          REG_43          : in    std_logic;
          REG_59          : out   std_logic;
          REG_164         : out   std_logic;
          REG_180         : out   std_logic;
          REG_132         : out   std_logic;
          REG_260         : out   std_logic;
          REG_116         : in    std_logic;
          REG_196         : out   std_logic;
          REG_244         : out   std_logic;
          REG_420         : out   std_logic;
          REG_469         : in    std_logic;
          REG_60          : out   std_logic;
          REG_44          : in    std_logic;
          REG_165         : out   std_logic;
          REG_181         : out   std_logic;
          REG_133         : out   std_logic;
          REG_261         : out   std_logic;
          REG_117         : in    std_logic;
          REG_197         : out   std_logic;
          REG_245         : out   std_logic;
          REG_421         : out   std_logic;
          REG_470         : in    std_logic;
          REG_61          : out   std_logic;
          REG_45          : in    std_logic;
          REG_166         : out   std_logic;
          REG_182         : out   std_logic;
          REG_134         : out   std_logic;
          REG_262         : out   std_logic;
          REG_118         : in    std_logic;
          REG_198         : out   std_logic;
          REG_246         : out   std_logic;
          REG_422         : out   std_logic;
          REG_455         : out   std_logic;
          REG_471         : in    std_logic;
          REG_423         : out   std_logic;
          REG_46          : in    std_logic;
          REG_62          : out   std_logic;
          REG_167         : out   std_logic;
          REG_183         : out   std_logic;
          REG_135         : out   std_logic;
          REG_263         : out   std_logic;
          REG_119         : in    std_logic;
          REG_199         : out   std_logic;
          REG_247         : out   std_logic;
          REG_63          : out   std_logic;
          REG_424         : out   std_logic;
          REG_64          : out   std_logic;
          REG_425         : out   std_logic;
          REG_65          : out   std_logic;
          REG_426         : out   std_logic;
          REG_66          : out   std_logic;
          REG_427         : out   std_logic;
          REG_67          : out   std_logic;
          REG_428         : out   std_logic;
          REG_68          : out   std_logic;
          REG_429         : out   std_logic;
          REG_69          : out   std_logic;
          REG_430         : out   std_logic;
          REG_70          : out   std_logic;
          REG_431         : out   std_logic;
          REG_71          : out   std_logic;
          REG_432         : out   std_logic;
          REG_72          : out   std_logic;
          REG_433         : out   std_logic;
          REG_73          : out   std_logic;
          REG_434         : out   std_logic;
          REG_74          : out   std_logic;
          REG_435         : out   std_logic;
          REG_75          : out   std_logic;
          REG_436         : out   std_logic;
          REG_76          : out   std_logic;
          REG_437         : out   std_logic;
          REG_77          : out   std_logic;
          REG_438         : out   std_logic;
          REG_78          : out   std_logic;
          REG_439         : out   std_logic;
          REG_4           : out   std_logic;
          REG_79          : out   std_logic;
          TST_c_c         : out   std_logic_vector(3 to 3);
          TST_c_4         : out   std_logic;
          TST_c_0         : out   std_logic;
          TST_c_5         : out   std_logic;
          TST_c_2         : out   std_logic;
          TST_c_1         : out   std_logic;
          REG_i_0_116     : out   std_logic;
          REG_i_0_0       : out   std_logic;
          REG_i_0_75      : out   std_logic;
          REG_i_0_260     : out   std_logic;
          REG_i_0_261     : out   std_logic;
          REG_i_0_275     : out   std_logic;
          REG_i_0_276     : out   std_logic;
          REG_i_0_277     : out   std_logic;
          REG_i_0_278     : out   std_logic;
          REG_i_0_279     : out   std_logic;
          REG_i_0_280     : out   std_logic;
          REG_i_0_281     : out   std_logic;
          REG_i_0_282     : out   std_logic;
          REG_i_0_283     : out   std_logic;
          REG_i_0_284     : out   std_logic;
          REG_i_0_285     : out   std_logic;
          REG_i_0_286     : out   std_logic;
          REG_i_0_287     : out   std_logic;
          REG_i_0_288     : out   std_logic;
          REG_i_0_289     : out   std_logic;
          REG_i_0_290     : out   std_logic;
          REG_i_0_291     : out   std_logic;
          REG_i_0_393     : out   std_logic;
          REG_i_0_391     : out   std_logic;
          REG_i_0_395     : out   std_logic;
          REG_i_0_388     : out   std_logic;
          REG_i_0_389     : out   std_logic;
          REG_i_0_390     : out   std_logic;
          REG_i_0_392     : out   std_logic;
          REG_i_0_394     : out   std_logic;
          REG_0           : out   std_logic_vector(127 downto 124);
          HWRES_c_16      : in    std_logic;
          HWRES_c_15      : in    std_logic;
          CLEAR_22        : in    std_logic;
          CLEAR_21        : in    std_logic;
          CLEAR_25        : in    std_logic;
          CLEAR_24        : in    std_logic;
          CLEAR_23        : in    std_logic;
          CLEAR_27        : in    std_logic;
          CLEAR_26        : in    std_logic;
          HWRES_c_18      : in    std_logic;
          HWRES_c_22      : in    std_logic;
          CLEAR_28        : in    std_logic;
          CLEAR           : in    std_logic;
          HWRES_c_17      : in    std_logic;
          HWRES_c_21      : in    std_logic;
          HWRES_c_12      : in    std_logic;
          HWRES_c_23      : in    std_logic;
          RAMRD           : out   std_logic;
          HWRES_c_19      : in    std_logic;
          OR_RACK         : out   std_logic;
          HWRES_c_14      : in    std_logic;
          OR_RREQ         : in    std_logic;
          HWRES_c_20      : in    std_logic;
          EF              : in    std_logic;
          CLEAR_20        : in    std_logic;
          ASB_c           : in    std_logic;
          un5_noe16ri_0_0 : out   std_logic;
          un7_noe32ri_0_0 : out   std_logic;
          WRITEB_c        : in    std_logic;
          nLBAS_c         : out   std_logic;
          LB_nOE          : out   std_logic;
          LWORDB_in       : in    std_logic;
          MYBERR_c        : out   std_logic;
          IACKB_c         : in    std_logic;
          nLBRDY_c        : in    std_logic;
          FWIMG2LOAD      : out   std_logic;
          NLBLAST_c       : out   std_logic;
          NLBRD_c         : out   std_logic;
          NLBCLR_c        : in    std_logic;
          EVREAD          : out   std_logic;
          NRDMEB          : out   std_logic;
          DTEST_FIFO      : in    std_logic;
          RUN_c           : out   std_logic;
          N_2052          : out   std_logic;
          d_m7            : in    std_logic;
          EV_RES_c        : in    std_logic;
          L0_c_c          : in    std_logic;
          L1A_c_c         : in    std_logic;
          L1R_c_c         : in    std_logic;
          L2A_c_c         : in    std_logic;
          L2R_c_c         : in    std_logic;
          LOS_c_c         : in    std_logic;
          N_441           : out   std_logic;
          SPULSE0_c_c     : in    std_logic;
          SPULSE1_c_c     : in    std_logic;
          SPULSE2_c_c     : in    std_logic;
          DS1B_c          : in    std_logic;
          DS0B_c          : in    std_logic;
          N_500           : out   std_logic;
          NDTKIN_c        : out   std_logic;
          NOE16W_c        : out   std_logic;
          NOE32W_c        : out   std_logic;
          NOEAD_c         : out   std_logic;
          NSELCLK_c       : out   std_logic;
          NSELCLK_c_i_0   : out   std_logic;
          CLEAR_0         : in    std_logic;
          EVRDY_c         : in    std_logic;
          HWRES_c_1       : in    std_logic;
          NOEAD_c_i_0     : out   std_logic;
          N_2613_0        : out   std_logic;
          RUN_c_0         : out   std_logic;
          HWRES_c_0       : in    std_logic;
          NOEAD_c_0       : out   std_logic;
          NOEAD_c_1       : out   std_logic;
          HWRES_c_22_0    : in    std_logic;
          ALICLK_c        : in    std_logic;
          un7_noe32ri_0   : out   std_logic;
          un5_noe16ri_0   : out   std_logic;
          WDOGTO          : out   std_logic;
          HWRES_c_0_6     : in    std_logic;
          HWRES_c_0_5     : in    std_logic;
          HWRES_c_0_4     : in    std_logic;
          HWRES_c_0_3     : in    std_logic;
          HWRES_c_23_0    : in    std_logic;
          HWRES_c_21_0    : in    std_logic;
          HWRES_c_13_0    : in    std_logic;
          HWRES_c_0_0     : in    std_logic;
          NOEAD_c_0_0     : out   std_logic;
          HWRES_c_13      : in    std_logic;
          CLK_c_c         : in    std_logic;
          RUN_c_0_0       : out   std_logic;
          HWRES_c_0_6_0   : in    std_logic
        );

end VINTERF;

architecture DEF_ARCH of VINTERF is 

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFF
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OAI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component LD
    port( EN : in    std_logic := 'U';
          D  : in    std_logic := 'U';
          Q  : out   std_logic
        );
  end component;

  component AOI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \un10_hwres_6_0\, WDOGTO_2, \REG3_514_180\, 
        un15_hwres_i, \un12_wdog_0_a3\, WDOGTO_1, WDOGTO_0, 
        \STATE1_0[1]_net_1\, \un10_hwres_32\, \STATE1_ns[9]\, 
        \TST_c_0[0]\, \ASBSF1\, \MBLTCYC\, \ADACKCYC\, 
        \un10_hwres_7_0\, \un10_hwres_8_0\, \un10_hwres_32_0\, 
        \REG_1_132\, \REG_1_133\, \REG_1_134\, \REG_1_135\, 
        \BLTCYC_2\, \BLTCYC_77\, \BLTCYC_1\, \BLTCYC_0\, 
        \SINGCYC_2\, \SINGCYC_147\, \SINGCYC_1\, \SINGCYC_0\, 
        \WRITES_1\, \WRITES_2\, \WRITES_0\, \REGMAP_0[2]_net_1\, 
        \un13_reg_ads_0_a2_0_a2\, \REGMAP_0[7]_net_1\, 
        \un33_reg_ads_0_a2_0_a2\, \REGMAP_0[16]_net_1\, 
        \un54_reg_ads_0_a3_0_a2\, \REGMAP_0[18]_net_1\, 
        \un61_reg_ads_0_a3_0_a2\, \REGMAP_0[19]_net_1\, 
        \un64_reg_ads_0_a3_0_a2\, \REGMAP_0[20]_net_1\, 
        \un67_reg_ads_0_a3_0_a2\, \REGMAP_0[24]_net_1\, 
        \un81_reg_ads_0_a3_0_a2\, \REGMAP_0[29]_net_1\, 
        \un105_reg_ads_0_a3_0_a2\, \STATE1_0[9]_net_1\, 
        \STATE1_ns[1]\, \STATE1_0[8]_net_1\, \STATE1_ns[2]\, 
        \STATE1_0[7]_net_1\, \STATE1_ns[3]\, \STATE1_1[2]_net_1\, 
        \STATE1_ns[8]\, \STATE1_0[2]_net_1\, \un10_hwres_35\, 
        \un10_hwres_34\, \un10_hwres_33\, \un10_hwres_31\, 
        \un10_hwres_30\, \un10_hwres_29\, \un10_hwres_28\, 
        \un10_hwres_27\, \un10_hwres_26\, \un10_hwres_25\, 
        \un10_hwres_24\, \un10_hwres_23\, \un10_hwres_22\, 
        \un10_hwres_21\, \un10_hwres_20\, \un10_hwres_19\, 
        \un10_hwres_18\, \un10_hwres_17\, \un10_hwres_16\, 
        \un10_hwres_15\, \un10_hwres_14\, \un10_hwres_13\, 
        \un10_hwres_12\, \un10_hwres_11\, \un10_hwres_10\, 
        \un10_hwres_9\, \un10_hwres_8\, \un10_hwres_7\, 
        \un10_hwres_6\, \un10_hwres_5\, \un10_hwres_4\, \WDOGTO\, 
        \un10_hwres_3\, \un10_hwres_2\, \un10_hwres_1\, 
        \un10_hwres_0\, \REGMAP_1[31]_net_1\, 
        \un111_reg_ads_0_a3_0_a2\, \REGMAP_0[31]_net_1\, 
        \REGMAP_1[28]_net_1\, \un102_reg_ads_0_a3_0_a2\, 
        \REGMAP_0[28]_net_1\, \REGMAP_0[26]_net_1\, 
        \un94_reg_ads_0_a3_0_a2\, \REGMAP_1[13]_net_1\, 
        \un84_reg_ads_0_a3_0_a2\, \REGMAP_0[13]_net_1\, N_566_1, 
        N_436, \NOEAD_c_0_0\, \un7_noe32ri_0_0_a2_0\, \LWORDS\, 
        \STATE5_3[0]_net_1\, \STATE5_ns[0]\, \STATE5_2[0]_net_1\, 
        \STATE5_1[0]_net_1\, \STATE5_0[0]_net_1\, 
        \STATE5_0[2]_net_1\, \STATE5_ns_i_0[2]_net_1\, N_83_0, 
        N_2524, N_2523_0, \REGMAP[15]_net_1\, N_1898, N_66_0, 
        \STATE5[1]_net_1\, \TST_c_0[1]\, N_2403, \TST_c_0[2]\, 
        \DSSF1\, \TST_c_1[5]\, \un37_reg_ads_0_a2_4_a2\, 
        \TST_c_0[5]\, N_85_4, \EVREAD_DS\, \STATE2[1]_net_1\, 
        N_85_3, N_85_2, N_85_1, N_85_0, N_7_i_1, N_425, N_7_i_0, 
        N_1996_4, N_426, \STATE2_i_0[3]\, N_1996_3, N_1996_2, 
        N_1996_1, N_1996_0, STATE5_0_sqmuxa_1, N_2608, N_2606_i_i, 
        STATE5_0_sqmuxa_0, LB_i_6_sn_N_2_1, LB_i_6_sn_N_2_0, 
        N_2572_3, N_2572_2, N_2572_1, N_2572_0, N_2511_0, 
        \REGMAP[6]_net_1\, un1_STATE1_34_1, N_2535, 
        \un1_STATE1_34_0_0\, \un1_STATE1_34_0\, 
        PULSE_0_sqmuxa_1_2, PULSE_0_sqmuxa_1_1, 
        PULSE_0_sqmuxa_1_0, un1_STATE2_13_4_1, \STATE2[2]_net_1\, 
        N_472_i_0, un1_STATE2_12_0_0_1_i, un1_STATE2_13_4_0, 
        un1_STATE2_16_1, un1_STATE2_16_0_0_0_i, N_79, N_580, 
        un1_STATE2_16_0, N_441_0, \REGMAP_i_i[33]\, 
        \REGMAP[34]_net_1\, N_2613_1, N_479, LB_DOUT_0_sqmuxa_1, 
        \REGMAP[36]_net_1\, LB_DOUT_0_sqmuxa_0, N_2033_0, 
        \REGMAP[30]_net_1\, N_2512_0, \VDBi_16_1_a2_3_0[1]_net_1\, 
        REG_0_sqmuxa_0, REG1_0_sqmuxa_0, \REGMAP[1]_net_1\, 
        N_2507_1, N_2507_0, \VDBi_9_sqmuxa_0\, \un776_regmap_23\, 
        \VDBi_9_sqmuxa_1\, \VDBi_9_sqmuxa_i_1\, N_616_1, N_428, 
        N_616_0, N_2570_1, \LB_WRITE_sync\, N_2603, N_2570_0, 
        N_2816_i_0_0, \REGMAP_i_i_0[23]\, 
        \un78_reg_ads_0_a3_0_a2\, N_457_i_0_1, \REGMAP[0]_net_1\, 
        N_457_i_0_0, N_3008_i_0, \REGMAP_i_i_0[33]\, 
        \un114_reg_ads_0_a3_0_a2\, N_2880_i_0, \REGMAP[25]_net_1\, 
        N_3234_i_1, N_2409, un1_STATE1_15, N_3234_i_0, N_3170_i_1, 
        N_3170_i_0, N_3104_i_0, N_3072_i_1, N_3072_i_0, 
        N_2976_i_0, N_2944_i_0, N_2784_i_0, N_2752_i_0, 
        N_2720_i_0, N_2688_i_0, \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \WDOG[1]_net_1\, \DWACT_ADD_CI_0_g_array_12_1[0]\, 
        \WDOG_i_0_i[4]\, \DWACT_ADD_CI_0_g_array_12[0]\, 
        \WDOG[2]_net_1\, \WDOGRES_i\, \WDOGRES\, 
        \STATE2_i[4]_net_1\, \STATE2[4]_net_1\, \NOEAD_c_0\, 
        WDOGRES1_i, N_2371_i_0, \REG[399]\, \REG[397]\, 
        \REG[395]\, \REG[394]\, \REG[393]\, \STATE2_ns_i[5]\, 
        N_1756, \STATE2[5]_net_1\, \REG[400]\, \REG[396]\, 
        \REG[398]\, \REG[296]\, \REG[295]\, \REG[294]\, 
        \REG[293]\, \REG[292]\, \REG[291]\, \REG[290]\, 
        \REG[289]\, \REG[288]\, \REG[287]\, \REG[286]\, 
        \REG[285]\, \REG[284]\, \REG[283]\, \REG[282]\, 
        \REG[281]\, \REG[280]\, \REG[266]\, \REG[265]\, 
        \NOE16W_c\, \CLOSEDTK\, N_488, \VDBi[21]_net_1\, 
        \PIPEB[21]_net_1\, \PIPEA[21]_net_1\, 
        \OR_RACK_1_sqmuxa_i_i_a2\, N_2597_1, \STATE5[2]_net_1\, 
        N_2540, \VDBi[11]_net_1\, \PIPEB[11]_net_1\, 
        \PIPEA[11]_net_1\, \TCNT_0_sqmuxa_i_s\, N_43, N_2532, 
        N_2561, \STATE1_tr27_i_0\, \STATE1_tr27_i_a2_0_0\, N_2533, 
        \DS_i_a2\, N_83, N_2327, \VDBi[31]_net_1\, 
        \PIPEB[31]_net_1\, \PIPEA[31]_net_1\, N_2326, 
        \VDBi[30]_net_1\, \PIPEB[30]_net_1\, \PIPEA[30]_net_1\, 
        N_2325, \VDBi[29]_net_1\, \PIPEB[29]_net_1\, 
        \PIPEA[29]_net_1\, N_2324, \VDBi[28]_net_1\, 
        \PIPEB_i_i[28]\, \PIPEA_i_0_i[28]\, N_2323, 
        \VDBi[27]_net_1\, \PIPEB[27]_net_1\, \PIPEA[27]_net_1\, 
        N_2322, \VDBi[26]_net_1\, \PIPEB[26]_net_1\, 
        \PIPEA[26]_net_1\, N_2321, \VDBi[25]_net_1\, 
        \PIPEB[25]_net_1\, \PIPEA[25]_net_1\, N_2320, 
        \VDBi[24]_net_1\, \PIPEB[24]_net_1\, \PIPEA[24]_net_1\, 
        N_2319, \VDBi[23]_net_1\, \PIPEB[23]_net_1\, 
        \PIPEA[23]_net_1\, N_2318, \VDBi[22]_net_1\, 
        \PIPEB[22]_net_1\, \PIPEA[22]_net_1\, N_2316, 
        \VDBi[20]_net_1\, \PIPEB[20]_net_1\, \PIPEA[20]_net_1\, 
        N_2315, \VDBi[19]_net_1\, \PIPEB[19]_net_1\, 
        \PIPEA[19]_net_1\, N_2314, \VDBi[18]_net_1\, 
        \PIPEB[18]_net_1\, \PIPEA[18]_net_1\, N_2313, 
        \VDBi[17]_net_1\, \PIPEB[17]_net_1\, \PIPEA[17]_net_1\, 
        N_2312, \VDBi[16]_net_1\, \PIPEB[16]_net_1\, 
        \PIPEA[16]_net_1\, N_2311, \VDBi[15]_net_1\, 
        \PIPEB[15]_net_1\, \PIPEA[15]_net_1\, N_2310, 
        \VDBi[14]_net_1\, \PIPEB[14]_net_1\, \PIPEA[14]_net_1\, 
        N_2309, \VDBi[13]_net_1\, \PIPEB[13]_net_1\, 
        \PIPEA[13]_net_1\, N_2308, \VDBi[12]_net_1\, 
        \PIPEB[12]_net_1\, \PIPEA[12]_net_1\, N_2306, 
        \VDBi[10]_net_1\, \PIPEB[10]_net_1\, \PIPEA[10]_net_1\, 
        N_2305, \VDBi[9]_net_1\, \PIPEB[9]_net_1\, 
        \PIPEA[9]_net_1\, N_2304, \VDBi[8]_net_1\, 
        \PIPEB[8]_net_1\, \PIPEA[8]_net_1\, N_2303, 
        \VDBi[7]_net_1\, \PIPEB[7]_net_1\, \PIPEA[7]_net_1\, 
        \BLTCYC\, N_2302, \VDBi[6]_net_1\, \PIPEB[6]_net_1\, 
        \PIPEA[6]_net_1\, N_2301, \VDBi[5]_net_1\, \SINGCYC\, 
        \PIPEB[5]_net_1\, \PIPEA[5]_net_1\, N_2300, 
        \VDBi[4]_net_1\, \PIPEB[4]_net_1\, \PIPEA[4]_net_1\, 
        N_2299, \VDBi[3]_net_1\, \PIPEB[3]_net_1\, 
        \PIPEA[3]_net_1\, N_2298, \VDBi[2]_net_1\, 
        \PIPEB[2]_net_1\, \PIPEA[2]_net_1\, N_2297, 
        \VDBi[1]_net_1\, \PIPEB[1]_net_1\, \PIPEA[1]_net_1\, 
        N_2296, \VDBi[0]_net_1\, \PIPEB[0]_net_1\, 
        \PIPEA[0]_net_1\, \un4_asb_NE\, \un4_asb_0\, \un4_asb_1\, 
        \un4_asb_NE_0\, \un4_asb_2\, \un4_asb_3\, \STATE1_ns[0]\, 
        \STATE1[10]_net_1\, \STATE1_ns_0_0[0]_net_1\, N_2410, 
        N_2429, N_2599_1, \LB_REQ_sync\, \STATE5_ns_i_0_0_i[2]\, 
        N_1861, N_2593_i, \OR_RREQ_sync\, \STATE5_ns[1]\, 
        \STATE5_ns_0_0_0_i[1]\, N_2595, N_2596, N_2607, N_2597, 
        \REQUESTER\, \STATE5_ns_0_0_0_i[0]\, N_2600, 
        \REQUESTER_1_i_0\, N_2589, \LB_ACK_1_sqmuxa_i_0\, 
        \STATE5_i_0[2]\, \STATE2_ns[4]\, N_725, \STATE2_ns[3]\, 
        \STATE2_ns_0_0_0[3]_net_1\, N_449, \STATE2_ns[0]\, N_1762, 
        N_1756_1, N_2552_1, \STATE1_ns_0_iv_0_a2_0_1[9]_net_1\, 
        N_2551_i, N_486, N_2531, N_2550, N_2550_1, \un776_regmap\, 
        \STATE1_ns[7]\, N_2430, N_2547, \STATE1[3]_net_1\, 
        \STATE1_ns[6]\, \STATE1[4]_net_1\, N_2612, \STATE1_ns[5]\, 
        \STATE1_ns_1_iv_0_0_a2_0_0[5]_net_1\, N_572_i, N_573_1, 
        N_462, N_480, \STATE1_ns[4]\, N_2413, N_570_i, 
        \STATE1[9]_net_1\, \STATE1[6]_net_1\, N_2565, 
        \STATE1_ns_1_iv_0_1[3]_net_1\, N_2544, N_2545, N_2542, 
        \REGMAP[10]_net_1\, \LB_ACK_sync\, \STATE1[0]_net_1\, 
        \STATE1_ns_0_iv_0_0_0_i[1]\, N_627, N_2431, N_629, 
        N_2455_1, \VDBi_652\, \VDBi_92[31]\, 
        \VDBi_92_0_iv_0_4_i[31]\, \VDBi_92_0_iv_0_2_i[31]\, 
        \VDBi_92_0_iv_0_1_i[31]\, N_615, \LB_s[31]_net_1\, N_792, 
        \VDBi_92_0_iv_0_0[31]_net_1\, N_610, N_723, N_790, N_612, 
        N_793, \REG[513]\, \VDBi_651\, \VDBi_92[30]\, 
        \VDBi_71[30]_net_1\, N_2613, \VDBi_92_0_iv_1[30]_net_1\, 
        \VDBi_60[30]_net_1\, \VDBi_55[30]_net_1\, 
        \VDBi_23[30]_net_1\, \VDBi_18[30]_net_1\, 
        \REG_i[512]_net_1\, \REG[512]\, \LB_s[30]_net_1\, 
        \VDBi_92_0_iv_0[30]_net_1\, \PIPEA_m[30]_net_1\, 
        \VDBi_650\, \VDBi_92[29]\, \VDBi_71[29]_net_1\, 
        \VDBi_92_0_iv_1[29]_net_1\, \VDBi_60[29]_net_1\, 
        \VDBi_55[29]_net_1\, \VDBi_23[29]_net_1\, 
        \VDBi_18[29]_net_1\, \REG_i[511]_net_1\, \REG[511]\, 
        \LB_s[29]_net_1\, \VDBi_92_0_iv_0[29]_net_1\, 
        \PIPEA_m[29]_net_1\, \VDBi_649\, \VDBi_92[28]\, 
        \VDBi_71[28]_net_1\, \VDBi_92_0_iv_1[28]_net_1\, 
        \VDBi_60[28]_net_1\, \VDBi_55[28]_net_1\, 
        \VDBi_23[28]_net_1\, \VDBi_18[28]_net_1\, 
        \REG_i[510]_net_1\, \REG[510]\, \LB_s[28]_net_1\, 
        \VDBi_92_0_iv_0[28]_net_1\, \PIPEA_m[28]_net_1\, 
        \VDBi_648\, \VDBi_92[27]\, \VDBi_71[27]_net_1\, 
        \VDBi_92_0_iv_1[27]_net_1\, \VDBi_60[27]_net_1\, 
        \VDBi_55[27]_net_1\, \VDBi_23[27]_net_1\, 
        \VDBi_18[27]_net_1\, \REG_i[509]_net_1\, \REG[509]\, 
        \LB_s[27]_net_1\, \VDBi_92_0_iv_0[27]_net_1\, 
        \PIPEA_m[27]_net_1\, \VDBi_647\, \VDBi_92[26]\, 
        \VDBi_71[26]_net_1\, \VDBi_92_0_iv_1[26]_net_1\, 
        \VDBi_60[26]_net_1\, \VDBi_55[26]_net_1\, 
        \VDBi_23[26]_net_1\, \VDBi_18[26]_net_1\, 
        \REG_i[508]_net_1\, \REG[508]\, \LB_s[26]_net_1\, 
        \VDBi_92_0_iv_0[26]_net_1\, \PIPEA_m[26]_net_1\, 
        \VDBi_646\, \VDBi_92[25]\, \VDBi_92_0_iv_0_4_i[25]\, 
        \VDBi_92_0_iv_0_2_i[25]\, \VDBi_92_0_iv_0_1_i[25]\, N_608, 
        \LB_s[25]_net_1\, \VDBi_92_0_iv_0_0[25]_net_1\, N_603, 
        N_605, \REG[507]\, \VDBi_645\, \VDBi_92[24]\, 
        \VDBi_71[24]_net_1\, \VDBi_92_0_iv_1[24]_net_1\, 
        \VDBi_60[24]_net_1\, \VDBi_55[24]_net_1\, 
        \VDBi_23[24]_net_1\, \VDBi_18[24]_net_1\, 
        \REG_i[506]_net_1\, \REG[506]\, \LB_s[24]_net_1\, 
        \VDBi_92_0_iv_0[24]_net_1\, \PIPEA_m[24]_net_1\, 
        \VDBi_644\, \VDBi_92[23]\, \VDBi_71[23]_net_1\, 
        \VDBi_92_0_iv_1[23]_net_1\, \VDBi_60[23]_net_1\, 
        \VDBi_55[23]_net_1\, \VDBi_23[23]_net_1\, 
        \VDBi_18[23]_net_1\, \REG_i[505]_net_1\, \REG[505]\, 
        \LB_s[23]_net_1\, \VDBi_92_0_iv_0[23]_net_1\, 
        \PIPEA_m[23]_net_1\, \VDBi_643\, \VDBi_92[22]\, 
        \VDBi_71[22]_net_1\, \VDBi_92_0_iv_1[22]_net_1\, 
        \VDBi_60[22]_net_1\, \VDBi_55[22]_net_1\, 
        \VDBi_23[22]_net_1\, \VDBi_18[22]_net_1\, 
        \REG_i[504]_net_1\, \REG[504]\, \LB_s[22]_net_1\, 
        \VDBi_92_0_iv_0[22]_net_1\, \PIPEA_m[22]_net_1\, 
        \VDBi_642\, \VDBi_92[21]\, \VDBi_92_0_iv_0_0_4_i[21]\, 
        \VDBi_92_0_iv_0_0_2_i[21]\, \VDBi_92_0_iv_0_0_1_i[21]\, 
        N_592, \LB_s[21]_net_1\, \VDBi_92_0_iv_0_0_0[21]_net_1\, 
        N_669, N_587, \N_2613_0\, N_589, N_680, \REG[503]\, 
        \VDBi_641\, \VDBi_92[20]\, \VDBi_71[20]_net_1\, 
        \VDBi_92_0_iv_1[20]_net_1\, \VDBi_60[20]_net_1\, 
        \VDBi_55[20]_net_1\, \REGMAP[26]_net_1\, 
        \VDBi_23[20]_net_1\, \VDBi_18[20]_net_1\, 
        \REG_i[502]_net_1\, \REG[502]\, \LB_s[20]_net_1\, 
        \VDBi_92_0_iv_0[20]_net_1\, \PIPEA_m[20]_net_1\, 
        \VDBi_640\, \VDBi_92[19]\, \VDBi_71[19]_net_1\, 
        \VDBi_92_0_iv_1[19]_net_1\, \VDBi_60[19]_net_1\, 
        \VDBi_55[19]_net_1\, \VDBi_23[19]_net_1\, 
        \VDBi_18[19]_net_1\, \REG[501]\, \LB_s[19]_net_1\, 
        \VDBi_92_0_iv_0[19]_net_1\, \PIPEA_m[19]_net_1\, 
        \VDBi_639\, \VDBi_92[18]\, \VDBi_71[18]_net_1\, 
        \VDBi_92_0_iv_1[18]_net_1\, \VDBi_60[18]_net_1\, 
        \VDBi_55[18]_net_1\, \VDBi_23[18]_net_1\, 
        \VDBi_18[18]_net_1\, \REG[500]\, \LB_s[18]_net_1\, 
        \VDBi_92_0_iv_0[18]_net_1\, \PIPEA_m[18]_net_1\, 
        \VDBi_638\, \VDBi_92[17]\, \VDBi_71[17]_net_1\, 
        \VDBi_92_0_iv_1[17]_net_1\, \VDBi_60[17]_net_1\, 
        \VDBi_55[17]_net_1\, \VDBi_23[17]_net_1\, 
        \VDBi_18[17]_net_1\, \REG_i[499]_net_1\, \REG[499]\, 
        \LB_s[17]_net_1\, \VDBi_92_0_iv_0[17]_net_1\, 
        \PIPEA_m[17]_net_1\, \VDBi_637\, \VDBi_92[16]\, 
        \VDBi_71[16]_net_1\, \VDBi_92_0_iv_1[16]_net_1\, 
        \VDBi_60[16]_net_1\, \VDBi_55[16]_net_1\, 
        \VDBi_23[16]_net_1\, \VDBi_18[16]_net_1\, 
        \REG_i[498]_net_1\, \REG[498]\, \LB_s[16]_net_1\, 
        \VDBi_92_0_iv_0[16]_net_1\, \PIPEA_m[16]_net_1\, 
        \VDBi_636\, \VDBi_92[15]\, \VDBi_77[15]_net_1\, 
        \VDBi_92_0_iv_1[15]_net_1\, \VDBi_66[15]_net_1\, 
        \VDBi_77_d[15]_net_1\, \VDBi_77_s[8]_net_1\, 
        \VDBi_60[15]_net_1\, N_2032, \VDBi_58[15]_net_1\, 
        \VDBi_53_0_iv_5_i[15]\, \VDBi_23_m_i[15]\, \VDBi_58_0[9]\, 
        \VDBi_53_0_iv_3_i[15]\, \VDBi_53_0_iv_0_i[15]\, 
        \VDBi_53_0_iv_1_i[15]\, \REGMAP_i_i[23]\, 
        \REG_1_m[200]_net_1\, \REGMAP[12]_net_1\, 
        \REG_1_m[264]_net_1\, \VDBi_53_0_iv_2[15]_net_1\, 
        \REG_1_m[168]_net_1\, \VDBi_23[15]_net_1\, 
        \VDBi_18[15]_net_1\, \REG[497]\, \VDBi_16[15]\, N_2497_i, 
        N_2496_i, \REGMAP[7]_net_1\, \REG[15]\, \REG[408]\, 
        \REG[392]\, N_2067, \LB_s[15]_net_1\, 
        \VDBi_92_0_iv_0[15]_net_1\, \PIPEA_m[15]_net_1\, 
        \VDBi_635\, \VDBi_92[14]\, \VDBi_77[14]_net_1\, 
        \VDBi_92_0_iv_1[14]_net_1\, \VDBi_71[14]_net_1\, N_2066, 
        \VDBi_66[14]_net_1\, \VDBi_60[14]_net_1\, N_2031, 
        \VDBi_58[14]_net_1\, \VDBi_53_0_iv_5_i[14]\, 
        \VDBi_23_m_i[14]\, \VDBi_53_0_iv_3_i[14]\, 
        \VDBi_53_0_iv_0_i[14]\, \VDBi_53_0_iv_1_i[14]\, 
        \REG_1_m[199]_net_1\, \REG_1_m[263]_net_1\, 
        \VDBi_53_0_iv_2[14]_net_1\, \REG_1_m[167]_net_1\, 
        \VDBi_23[14]_net_1\, \VDBi_16[14]\, \VDBi_23_d[14]_net_1\, 
        \VDBi_23_s[7]_net_1\, N_2495_i, N_2494_i, \REG[14]\, 
        \REG[496]\, \REG[407]\, \REG[391]\, \REG[455]\, 
        \LB_s[14]_net_1\, \VDBi_92_0_iv_0[14]_net_1\, 
        \PIPEA_m[14]_net_1\, \VDBi_634\, \VDBi_92[13]\, 
        \VDBi_77[13]_net_1\, \VDBi_92_0_iv_1[13]_net_1\, 
        \VDBi_71[13]_net_1\, N_2065, \VDBi_66[13]_net_1\, 
        \VDBi_60[13]_net_1\, N_2030, \VDBi_58[13]_net_1\, 
        \VDBi_53_0_iv_5_i[13]\, \VDBi_23_m_i[13]\, 
        \VDBi_53_0_iv_3_i[13]\, \VDBi_53_0_iv_0_i[13]\, 
        \VDBi_53_0_iv_1_i[13]\, \REG_1_m[198]_net_1\, 
        \REG_1_m[262]_net_1\, \VDBi_53_0_iv_2[13]_net_1\, 
        \REG_1_m[166]_net_1\, \VDBi_23[13]_net_1\, \VDBi_16[13]\, 
        \VDBi_23_d[13]_net_1\, N_2493_i, N_2492_i, \REG[13]\, 
        \REG[495]\, \REG[406]\, \REG[390]\, \REG[454]\, 
        \LB_s[13]_net_1\, \VDBi_92_0_iv_0[13]_net_1\, 
        \PIPEA_m[13]_net_1\, \VDBi_633\, \VDBi_92[12]\, N_502, 
        \VDBi_92_0_iv_0_1[12]_net_1\, N_495, N_496, 
        \VDBi_66[12]_net_1\, \REGMAP[31]_net_1\, 
        \VDBi_66_d[12]_net_1\, \VDBi_58[12]_net_1\, 
        \VDBi_66_s[1]_net_1\, N_2029, \REG[405]\, \REG[389]\, 
        \VDBi_53_0_iv_5_i[12]\, N_412_i, \VDBi_53_0_iv_3_i[12]\, 
        \VDBi_53_0_iv_0_i[12]\, \VDBi_53_0_iv_1_i[12]\, 
        \REG_1_m[197]_net_1\, \REG_1_m[261]_net_1\, 
        \VDBi_53_0_iv_2[12]_net_1\, \REG_1_m[165]_net_1\, N_494, 
        N_497, \REG[494]\, \VDBi_16[12]\, N_2491_i, N_2490_i, 
        \REG[12]\, \REG[453]\, \LB_s[12]_net_1\, 
        \VDBi_92_0_iv_0_0[12]_net_1\, N_599, \VDBi_632\, 
        \VDBi_92[11]\, \VDBi_77[11]_net_1\, 
        \VDBi_92_0_iv_1[11]_net_1\, \VDBi_71[11]_net_1\, N_2063, 
        \VDBi_66[11]_net_1\, \VDBi_66_d[11]_net_1\, 
        \VDBi_58[11]_net_1\, N_2028, \REG[404]\, \REG[388]\, 
        \VDBi_53_0_iv_5_i[11]\, \VDBi_23_m_i[11]\, 
        \VDBi_53_0_iv_3_i[11]\, \VDBi_53_0_iv_0_i[11]\, 
        \VDBi_53_0_iv_1_i[11]\, \REG_1_m[196]_net_1\, 
        \REG_1_m[260]_net_1\, \VDBi_53_0_iv_2[11]_net_1\, 
        \REG_1_m[164]_net_1\, \VDBi_23[11]_net_1\, 
        \VDBi_18[11]_net_1\, \REG[493]\, \REGMAP[13]_net_1\, 
        \VDBi_16[11]\, \TST_c[5]\, N_2489_i, N_2488_i, \REG[11]\, 
        \REG[452]\, \LB_s[11]_net_1\, \VDBi_92_0_iv_0[11]_net_1\, 
        \PIPEA_m[11]_net_1\, \VDBi_631\, \VDBi_92[10]\, N_503, 
        \VDBi_92_0_iv_0_0_1[10]_net_1\, N_490, N_2062, 
        \VDBi_66[10]_net_1\, \VDBi_60[10]_net_1\, N_2027, 
        \VDBi_58[10]_net_1\, \REGMAP[28]_net_1\, 
        \VDBi_53_0_iv_5_i[10]\, \VDBi_23_m_i[10]\, 
        \VDBi_53_0_iv_3_i[10]\, \VDBi_53_0_iv_0_i[10]\, 
        \VDBi_53_0_iv_1_i[10]\, \REG_1_m[195]_net_1\, 
        \REG_1_m[259]_net_1\, \VDBi_53_0_iv_2[10]_net_1\, 
        \REG_1_m[163]_net_1\, \VDBi_23[10]_net_1\, \VDBi_16[10]\, 
        \VDBi_23_d[10]_net_1\, N_2487_i, N_2486_i, \REG[10]\, 
        \REG[492]\, \REG[403]\, \REG[387]\, \REG[451]\, 
        \LB_s[10]_net_1\, \VDBi_92_0_iv_0_0_0[10]_net_1\, N_624, 
        \VDBi_630\, \VDBi_92[9]\, un1_STATE1_34, 
        \VDBi_77[9]_net_1\, \VDBi_92_0_iv_1[9]_net_1\, 
        \VDBi_71[9]_net_1\, N_2061, \N_441\, \VDBi_66[9]_net_1\, 
        \VDBi_60[9]_net_1\, N_2026, N_2033, \VDBi_58[9]_net_1\, 
        \RUN_c_0_0\, \VDBi_53_0_iv_5_i[9]\, \VDBi_23_m_i[9]\, 
        \VDBi_53_0_iv_3_i[9]\, \VDBi_53_0_iv_0_i[9]\, 
        \VDBi_53_0_iv_1_i[9]\, \REG_1_m[194]_net_1\, 
        \REG_1_m[258]_net_1\, \REGMAP[16]_net_1\, 
        \VDBi_53_0_iv_2[9]_net_1\, \REG_1_m[162]_net_1\, 
        \VDBi_23[9]_net_1\, \VDBi_16[9]\, \VDBi_23_d[9]_net_1\, 
        N_2485_i, N_2484_i, \REG[9]\, \REG[491]\, \REG[402]\, 
        \REG[386]\, \REGMAP[29]_net_1\, \REG[450]\, 
        \LB_s[9]_net_1\, N_7_i, \VDBi_92_0_iv_0[9]_net_1\, 
        \PIPEA_m[9]_net_1\, N_457_i_0, \VDBi_629\, \VDBi_92[8]\, 
        \VDBi_77[8]_net_1\, \VDBi_92_0_iv_1[8]_net_1\, 
        \VDBi_66[8]_net_1\, \VDBi_77_d[8]_net_1\, 
        \VDBi_60[8]_net_1\, N_2025, \VDBi_60_d[8]_net_1\, 
        \VDBi_55[8]_net_1\, \VDBi_60_s[5]_net_1\, 
        \VDBi_23_m_i[8]\, \VDBi_53_0_iv_6_i[8]\, 
        \VDBi_53_0_iv_5_i[8]\, \VDBi_53_0_iv_2_i[8]\, 
        \VDBi_53_0_iv_0_i[8]\, \REGMAP_i_i[17]\, 
        \REG_m[113]_net_1\, \REG_1_m[177]_net_1\, 
        \VDBi_53_0_iv_3_i[8]\, \REG_1_m_i[241]\, \REG_1_m_i[257]\, 
        \REG_1_m[129]_net_1\, \VDBi_23[8]_net_1\, 
        \VDBi_18[8]_net_1\, \REG[490]\, \VDBi_16[8]\, 
        \VDBi_16_1_0_i[8]\, N_2482_i, \REG[24]\, N_2483, N_2512, 
        \REG[401]\, \NSELCLK_c\, N_2060, \REG[449]\, 
        \LB_s[8]_net_1\, \VDBi_92_0_iv_0[8]_net_1\, 
        \STATE1[2]_net_1\, \PIPEA_m[8]_net_1\, \VDBi_628\, 
        \VDBi_92[7]\, N_508, \VDBi_92_iv_0_2[7]_net_1\, N_476, 
        N_492, N_493, \VDBi_60[7]_net_1\, 
        \VDBi_71_i_m2_d[7]_net_1\, \VDBi_71_s[4]_net_1\, 
        \VDBi_58[7]_net_1\, \VDBi_53_0_iv_5_i[7]\, 
        \VDBi_23_m_i[7]\, \VDBi_53_0_iv_3_i[7]\, 
        \VDBi_53_0_iv_0_i[7]\, \VDBi_53_0_iv_1_i[7]\, 
        \REG_1_m[192]_net_1\, \REGMAP[20]_net_1\, 
        \REG_1_m[256]_net_1\, \REGMAP[24]_net_1\, \REG[128]\, 
        \VDBi_53_0_iv_2[7]_net_1\, \REGMAP[19]_net_1\, 
        \REG_1_m[160]_net_1\, \REGMAP[18]_net_1\, \VDBi_9_sqmuxa\, 
        \VDBi_23[7]_net_1\, \VDBi_16[7]\, \VDBi_23_d[7]_net_1\, 
        \VDBi_16_1_0_i[7]\, N_2479_i, \REGMAP[2]_net_1\, N_2480, 
        \REG[7]\, N_2511, \REG[489]\, N_2024, \REG[448]\, 
        \LB_s[7]_net_1\, \VDBi_92_iv_0_1[7]_net_1\, 
        \VDBi_92_iv_0_0[7]_net_1\, \RAMDTS[7]_net_1\, N_596, 
        \VDBi_627\, \VDBi_92[6]\, \VDBi_80[6]_net_1\, 
        \VDBi_92_iv_2[6]_net_1\, \VDBi_71[6]_net_1\, 
        \VDBi_80_d[6]_net_1\, \VDBi_80_s[2]_net_1\, 
        \VDBi_58[6]_net_1\, \VDBi_71_d[6]_net_1\, 
        \VDBi_71_s[1]_net_1\, \VDBi_55[6]_net_1\, 
        \REGMAP[27]_net_1\, \VDBi_23_m_i[6]\, 
        \VDBi_53_0_iv_5_i[6]\, \VDBi_53_0_iv_3_i[6]\, 
        \VDBi_53_0_iv_0_i[6]\, \VDBi_53_0_iv_1_i[6]\, 
        \REG_1_m[191]_net_1\, \REG_1_m[255]_net_1\, \REG_0[127]\, 
        \VDBi_53_0_iv_2[6]_net_1\, \REG_1_m[159]_net_1\, 
        \VDBi_23[6]_net_1\, N_491, \REG[488]\, \VDBi_16[6]\, 
        \VDBi_16_1_0_i[6]\, N_2476_i, N_2477, 
        \VDBi_66_d[6]_net_1\, N_2023, N_2058, \REGMAP[35]_net_1\, 
        \REG[447]\, \LB_s[6]_net_1\, \VDBi_92_iv_1[6]_net_1\, 
        \VDBi_92_iv_0[6]_net_1\, \RAMDTS[6]_net_1\, 
        \FBOUT_m[6]_net_1\, \VDBi_626\, \VDBi_92[5]\, 
        \VDBi_80[5]_net_1\, \VDBi_92_iv_2[5]_net_1\, 
        \VDBi_77[5]_net_1\, \VDBi_66[5]_net_1\, 
        \VDBi_77_d[5]_net_1\, \VDBi_60[5]_net_1\, N_2022, 
        \VDBi_60_d[5]_net_1\, \VDBi_55[5]_net_1\, 
        \VDBi_23_m_i[5]\, \VDBi_53_0_iv_5_i[5]\, 
        \VDBi_53_0_iv_3_i[5]\, \VDBi_53_0_iv_0_i[5]\, 
        \VDBi_53_0_iv_1_i[5]\, \REG_1_m[190]_net_1\, 
        \REG_1_m[254]_net_1\, \REG_0[126]\, 
        \VDBi_53_0_iv_2[5]_net_1\, \REG_1_m[158]_net_1\, 
        \VDBi_23[5]_net_1\, \VDBi_16[5]\, \VDBi_23_d[5]_net_1\, 
        \VDBi_16_1_0_i[5]\, N_2473_i, N_2474, \REG[5]\, 
        \REG[487]\, N_2057, \LB_s[5]_net_1\, 
        \VDBi_92_iv_1[5]_net_1\, \VDBi_92_iv_0[5]_net_1\, 
        \RAMDTS[5]_net_1\, \STATE1[1]_net_1\, \FBOUT_m[5]_net_1\, 
        \VDBi_625\, \VDBi_92[4]\, \VDBi_80[4]_net_1\, 
        \VDBi_92_iv_2[4]_net_1\, \VDBi_77[4]_net_1\, 
        \VDBi_77_d[4]_net_1\, \VDBi_60[4]_net_1\, 
        \VDBi_77_s[3]_net_1\, \VDBi_71_d[4]_net_1\, N_2056, 
        N_2021, \VDBi_58[4]_net_1\, \VDBi_55[4]_net_1\, 
        \VDBi_23_m_i[4]\, \VDBi_53_0_iv_5_i[4]\, 
        \VDBi_53_0_iv_3_i[4]\, \VDBi_53_0_iv_0_i[4]\, 
        \VDBi_53_0_iv_1_i[4]\, \REG_1_m[189]_net_1\, 
        \REG_1_m[253]_net_1\, \REG_0[125]\, 
        \VDBi_53_0_iv_2[4]_net_1\, \REG_1_m[157]_net_1\, 
        \VDBi_23[4]_net_1\, \VDBi_16[4]\, \VDBi_23_d[4]_net_1\, 
        \VDBi_16_1_0_i[4]\, N_2470_i, N_2471, \REG[4]\, 
        \REG[486]\, \LB_s[4]_net_1\, \VDBi_92_iv_1[4]_net_1\, 
        \VDBi_92_iv_0[4]_net_1\, \RAMDTS[4]_net_1\, 
        \FBOUT_m[4]_net_1\, \VDBi_624\, \VDBi_92[3]\, 
        \VDBi_80[3]_net_1\, \VDBi_92_iv_2[3]_net_1\, 
        \VDBi_80_d[3]_net_1\, \VDBi_60[3]_net_1\, 
        \VDBi_80_s[3]_net_1\, \VDBi_77_d[3]_net_1\, 
        \VDBi_71_d[3]_net_1\, N_2055, N_2020, \VDBi_58[3]_net_1\, 
        \VDBi_55[3]_net_1\, \VDBi_23_m_i[3]\, 
        \VDBi_53_0_iv_5_i[3]\, \VDBi_53_0_iv_3_i[3]\, 
        \VDBi_53_0_iv_0_i[3]\, \VDBi_53_0_iv_1_i[3]\, 
        \REG_1_m[188]_net_1\, \REG_1_m[252]_net_1\, \REG_0[124]\, 
        \VDBi_53_0_iv_2[3]_net_1\, \REG_1_m[156]_net_1\, 
        \VDBi_23[3]_net_1\, \VDBi_18[3]_net_1\, \REG[485]\, 
        \VDBi_16[3]\, \VDBi_16_1_0_i[3]\, N_2467_i, \REG[19]\, 
        N_2468, \REG[3]\, \LB_s[3]_net_1\, 
        \VDBi_92_iv_1[3]_net_1\, \VDBi_92_iv_0[3]_net_1\, 
        \RAMDTS[3]_net_1\, \FBOUT_m[3]_net_1\, \VDBi_623\, 
        \VDBi_92[2]\, \VDBi_80[2]_net_1\, \VDBi_92_iv_2[2]_net_1\, 
        \VDBi_71[2]_net_1\, \VDBi_80_d[2]_net_1\, 
        \VDBi_60[2]_net_1\, \VDBi_71_d[2]_net_1\, 
        \VDBi_60_d[2]_net_1\, \VDBi_55[2]_net_1\, \VDBi_53[2]\, 
        \VDBi_23[2]_net_1\, \VDBi_53_0_iv_5[2]_net_1\, 
        \VDBi_18[2]_net_1\, \REG[484]\, \VDBi_16[2]\, N_2464_i, 
        \VDBi_16_1_0_i[2]\, N_2465, \REG[2]\, 
        \VDBi_53_0_iv_3_i[2]\, \VDBi_53_0_iv_0_i[2]\, 
        \VDBi_53_0_iv_1_i[2]\, \REG_1_m[187]_net_1\, 
        \REG_1_m[251]_net_1\, \VDBi_53_0_iv_2[2]_net_1\, 
        \REG_1_m[155]_net_1\, N_2019, N_2054, \LB_s[2]_net_1\, 
        \VDBi_92_iv_1[2]_net_1\, \VDBi_92_iv_0[2]_net_1\, 
        \RAMDTS[2]_net_1\, \FBOUT_m[2]_net_1\, \VDBi_622\, 
        \VDBi_92[1]\, \VDBi_80[1]_net_1\, \VDBi_92_iv_2[1]_net_1\, 
        \VDBi_71[1]_net_1\, \VDBi_80_d[1]_net_1\, 
        \VDBi_71_d_0[1]_net_1\, \VDBi_55[1]_net_1\, 
        \VDBi_71_s_0[1]_net_1\, \VDBi_71_d[1]_net_1\, 
        \VDBi_66_d[1]_net_1\, N_2018, \VDBi_53[1]\, 
        \VDBi_23[1]_net_1\, \VDBi_53_0_iv_6[1]_net_1\, 
        \VDBi_18[1]_net_1\, \REG[483]\, \VDBi_16[1]\, N_2461_i, 
        \VDBi_16_1_0_i[1]\, N_2462, \REG[1]\, 
        \VDBi_53_0_iv_5_i[1]\, \VDBi_53_0_iv_2_i[1]\, 
        \VDBi_53_0_iv_0_i[1]\, \REG_m[106]_net_1\, 
        \REG_1_m[170]_net_1\, \VDBi_53_0_iv_3_i[1]\, 
        \REG_1_m_i[234]\, \REG_1_m_i[250]\, \REG_1_m[122]_net_1\, 
        N_2053, \LB_s[1]_net_1\, \VDBi_92_iv_1[1]_net_1\, 
        \VDBi_92_iv_0[1]_net_1\, \RAMDTS[1]_net_1\, 
        \FBOUT_m[1]_net_1\, \VDBi_621\, \VDBi_92[0]\, 
        un1_STATE1_34_0_a2_1_1_i, \VDBi_80_m_i_i[0]\, 
        \VDBi_92_iv_1_i[0]\, \LB_s_m_i[0]\, \LB_s[0]_net_1\, 
        \VDBi_92_iv_0[0]_net_1\, \RAMDTS[0]_net_1\, 
        \FBOUT_m[0]_net_1\, \VDBi_66[0]_net_1\, 
        \VDBi_80_m_0_m4_0_a2\, VDBi_80_m_0_m4_0_a2_1_i, 
        \REGMAP[32]_net_1\, \VDBi_60[0]_net_1\, N_2017, 
        \VDBi_60_d[0]_net_1\, \VDBi_53[0]\, \VDBi_60_s[0]_net_1\, 
        \VDBi_58_d[0]_net_1\, \VDBi_23[0]_net_1\, 
        \VDBi_53_0_iv_6[0]_net_1\, \VDBi_21[0]_net_1\, \REG[482]\, 
        \VDBi_18[0]_net_1\, \REG[80]\, \REGMAP[9]_net_1\, 
        \VDBi_16[0]\, \VDBi_16_1_1_i[0]\, N_2377_i, N_2380_1, 
        \VDBi_16_1_a3_1_0[0]_net_1\, \VDBi_16_1_0[0]_net_1\, 
        \REGMAP[14]_net_1\, N_2380, \VDBi_16_1_a3_2_0[0]_net_1\, 
        \REG_c[0]\, \REGMAP_i_0[12]\, \VDBi_9_sqmuxa_i_0\, 
        \VDBi_53_0_iv_5_i[0]\, \VDBi_53_0_iv_2_i[0]\, 
        \VDBi_53_0_iv_0_i[0]\, \REG_m[105]_net_1\, 
        \REG_1_m[169]_net_1\, \VDBi_53_0_iv_3_i[0]\, 
        \REG_1_m_i[233]\, \REG_1_m_i[249]\, \REG_1_m[121]_net_1\, 
        \PIPEA_620\, \PIPEA_7[31]\, N_366, \PIPEA1[31]_net_1\, 
        \PIPEA_619\, \PIPEA_7[30]\, N_539, \PIPEA1[30]_net_1\, 
        \PIPEA_618\, \PIPEA_7[29]\, N_538, \PIPEA1[29]_net_1\, 
        \PIPEA_617\, \PIPEA_7[28]\, N_537, \PIPEA1[28]_net_1\, 
        \PIPEA_616\, \PIPEA_7[27]\, N_536, \PIPEA1[27]_net_1\, 
        \PIPEA_615\, \PIPEA_7[26]\, N_535, \PIPEA1[26]_net_1\, 
        \PIPEA_614\, \PIPEA_7[25]\, N_534, \PIPEA1[25]_net_1\, 
        \PIPEA_613\, \PIPEA_7[24]\, N_533, \PIPEA1[24]_net_1\, 
        \PIPEA_612\, \PIPEA_7[23]\, N_532, \PIPEA1[23]_net_1\, 
        \PIPEA_611\, \PIPEA_7[22]\, N_531, \PIPEA1[22]_net_1\, 
        \PIPEA_610\, \PIPEA_7[21]\, N_530, \PIPEA1[21]_net_1\, 
        \PIPEA_609\, \PIPEA_7[20]\, N_529, \PIPEA1[20]_net_1\, 
        \PIPEA_608\, \PIPEA_7[19]\, N_528, \PIPEA1[19]_net_1\, 
        \PIPEA_607\, \PIPEA_7[18]\, N_527, \PIPEA1[18]_net_1\, 
        \PIPEA_606\, \PIPEA_7[17]\, N_526, \PIPEA1[17]_net_1\, 
        \PIPEA_605\, \PIPEA_7[16]\, N_525, \PIPEA1[16]_net_1\, 
        \PIPEA_604\, \PIPEA_7[15]\, N_524, \PIPEA1[15]_net_1\, 
        \PIPEA_603\, \PIPEA_7[14]\, N_523, \PIPEA1[14]_net_1\, 
        \PIPEA_602\, \PIPEA_7[13]\, N_522, \PIPEA1[13]_net_1\, 
        \PIPEA_601\, \PIPEA_7[12]\, N_521, \PIPEA1[12]_net_1\, 
        \PIPEA_600\, \PIPEA_7[11]\, N_520, \PIPEA1[11]_net_1\, 
        \PIPEA_599\, \PIPEA_7[10]\, N_519, \PIPEA1[10]_net_1\, 
        \PIPEA_598\, \PIPEA_7[9]\, un1_STATE2_16, N_518, 
        \PIPEA1[9]_net_1\, \PIPEA_597\, \PIPEA_7[8]\, N_517, 
        \PIPEA1[8]_net_1\, \PIPEA_596\, \PIPEA_7[7]\, N_516, 
        \PIPEA1[7]_net_1\, \PIPEA_595\, \PIPEA_7[6]\, N_515, 
        \PIPEA1[6]_net_1\, \PIPEA_594\, \PIPEA_7[5]\, N_514, 
        \PIPEA1[5]_net_1\, \PIPEA_593\, \PIPEA_7[4]\, N_513, 
        \PIPEA1[4]_net_1\, \PIPEA_592\, \PIPEA_7[3]\, N_512, 
        \PIPEA1[3]_net_1\, \PIPEA_591\, \PIPEA_7[2]\, N_511, 
        \PIPEA1[2]_net_1\, \PIPEA_590\, \PIPEA_7[1]\, N_510, 
        \PIPEA1[1]_net_1\, \PIPEA_589\, \PIPEA_7[0]\, N_509, 
        \PIPEA1[0]_net_1\, \NRDMEBi_588\, N_42_i_0, 
        \un1_NRDMEBi_2_sqmuxa_1_i_a3_i\, N_584, \EFS\, N_622, 
        N_7139_i, N_2499_i, un1_NRDMEBi_2_sqmuxa_2_i_1_i, N_2500, 
        \STATE2[0]_net_1\, N_583, \PIPEA1_587\, N_296, 
        \PIPEA1_586\, \PIPEA1_9[30]\, \PIPEA1_585\, 
        \PIPEA1_9[29]\, \PIPEA1_584\, \PIPEA1_9[28]\, 
        \PIPEA1_583\, N_294, \PIPEA1_582\, N_292, \PIPEA1_581\, 
        N_290, \PIPEA1_580\, N_288, \PIPEA1_579\, N_286, 
        \PIPEA1_578\, N_284, \PIPEA1_577\, N_282, \PIPEA1_576\, 
        N_280, \PIPEA1_575\, N_278, \PIPEA1_574\, N_276, 
        \PIPEA1_573\, N_274, \PIPEA1_572\, N_272, \PIPEA1_571\, 
        N_270, \PIPEA1_570\, N_268, \PIPEA1_569\, N_266, 
        \PIPEA1_568\, N_264, \PIPEA1_567\, N_262, \PIPEA1_566\, 
        N_260, \PIPEA1_565\, N_258, un1_STATE2_13_4, \PIPEA1_564\, 
        N_256, N_85, \PIPEA1_563\, N_254, \PIPEA1_562\, N_252, 
        \PIPEA1_561\, N_250, \PIPEA1_560\, N_248, \PIPEA1_559\, 
        N_246, \PIPEA1_558\, N_244, \PIPEA1_557\, N_242, 
        \PIPEA1_556\, N_238, N_620_i_i, N_485, \END_PK\, 
        \END_PK_555\, N_44, \un1_STATE2_13_i_0_a2_0_0\, N_581, 
        N_582_1, N_459, N_450_i, N_676, N_440, N_77_i_i_o2_1_i, 
        N_652, \un1_STATE2_13_i_0_a2_1_0_0\, \LB_ADDR_554\, 
        \LB_ADDR[11]_net_1\, \VAS[11]_net_1\, LB_ADDR_0_sqmuxa_2, 
        \LB_ADDR_553\, \LB_ADDR[10]_net_1\, \VAS[10]_net_1\, 
        \LB_ADDR_552\, \LB_ADDR[9]_net_1\, \VAS[9]_net_1\, 
        \LB_ADDR_551\, \LB_ADDR[8]_net_1\, \VAS[8]_net_1\, 
        \LB_ADDR_550\, \LB_ADDR[7]_net_1\, \VAS[7]_net_1\, 
        \LB_ADDR_549\, \LB_ADDR[6]_net_1\, \VAS[6]_net_1\, 
        \LB_ADDR_548\, \LB_ADDR[5]_net_1\, \VAS[5]_net_1\, 
        \LB_ADDR_547\, \LB_ADDR[4]_net_1\, \VAS[4]_net_1\, 
        \LB_ADDR_546\, \LB_ADDR[3]_net_1\, \VAS[3]_net_1\, 
        \LB_ADDR_545\, \LB_ADDR[2]_net_1\, \VAS[2]_net_1\, 
        \LB_ADDR_544\, \LB_ADDR[1]_net_1\, \VAS[1]_net_1\, 
        \LB_ADDR_0_sqmuxa_1\, \LB_i_543\, \LB_i_6[31]\, N_2213, 
        \LB_DOUT[31]_net_1\, \LB_i_542\, \LB_i_6[30]\, N_2212, 
        \LB_DOUT[30]_net_1\, \LB_i_541\, \LB_i_6[29]\, N_2211, 
        \LB_DOUT[29]_net_1\, \LB_i_540\, \LB_i_6[28]\, N_2210, 
        \LB_DOUT[28]_net_1\, \LB_i_539\, \LB_i_6[27]\, N_2209, 
        \LB_DOUT[27]_net_1\, \LB_i_538\, \LB_i_6[26]\, N_2208, 
        \LB_DOUT[26]_net_1\, \LB_i_537\, \LB_i_6[25]\, N_2207, 
        \LB_DOUT[25]_net_1\, \LB_i_536\, \LB_i_6[24]\, N_2206, 
        \LB_DOUT[24]_net_1\, \LB_i_535\, \LB_i_6[23]\, N_2205, 
        \LB_DOUT[23]_net_1\, \LB_i_534\, \LB_i_6[22]\, N_2204, 
        \LB_DOUT[22]_net_1\, \LB_i_533\, \LB_i_6[21]\, N_2203, 
        \LB_DOUT[21]_net_1\, \LB_i_532\, \LB_i_6[20]\, N_2202, 
        \LB_DOUT[20]_net_1\, \LB_i_531\, \LB_i_6[19]\, N_2201, 
        \LB_DOUT[19]_net_1\, \LB_i_530\, \LB_i_6[18]\, N_2200, 
        \LB_DOUT[18]_net_1\, \LB_i_529\, \LB_i_6[17]\, N_2199, 
        \LB_DOUT[17]_net_1\, \LB_i_528\, \LB_i_6[16]\, N_2198, 
        \LB_DOUT[16]_net_1\, \LB_i_527\, \LB_i_6[15]\, N_2197, 
        \LB_DOUT[15]_net_1\, \LB_i_526\, \LB_i_6[14]\, N_2196, 
        \LB_DOUT[14]_net_1\, \LB_i_525\, \LB_i_6[13]\, N_2195, 
        \LB_DOUT[13]_net_1\, \LB_i_524\, \LB_i_6[12]\, N_2194, 
        \LB_DOUT[12]_net_1\, \LB_i_523\, \LB_i_6[11]_net_1\, 
        N_2227, N_2181, N_2193, \LB_DOUT[11]_net_1\, \LB_i_522\, 
        \LB_i_6[10]_net_1\, N_2226, N_2180, N_2192, 
        \LB_DOUT[10]_net_1\, \LB_i_521\, \LB_i_6[9]_net_1\, 
        N_2570, N_2225, N_2179, N_2191, LB_i_6_sn_N_2, 
        \LB_DOUT[9]_net_1\, \LB_i_520\, \LB_i_6[8]_net_1\, N_2224, 
        N_2178, N_2190, \LB_DOUT[8]_net_1\, \LB_i_519\, 
        \LB_i_6[7]_net_1\, N_2223, N_2177, N_2189, 
        \LB_DOUT[7]_net_1\, \LB_i_518\, \LB_i_6[6]_net_1\, N_2222, 
        N_2176, N_2188, \LB_DOUT[6]_net_1\, \LB_i_517\, 
        \LB_i_6[5]_net_1\, N_2221, N_2175, N_2187, 
        \LB_DOUT[5]_net_1\, \LB_i_516\, \LB_i_6[4]_net_1\, N_2220, 
        N_2174, N_2186, \LB_DOUT[4]_net_1\, \LB_i_515\, 
        \LB_i_6[3]_net_1\, N_2219, N_2173, N_2185, 
        \STATE5[0]_net_1\, \LB_DOUT[3]_net_1\, \LB_i_514\, 
        \LB_i_6[2]_net_1\, N_2218, N_2172, N_2184, 
        \LB_DOUT[2]_net_1\, \LB_i_513\, \LB_i_6[1]_net_1\, N_2217, 
        N_2171, N_2183, \LB_DOUT[1]_net_1\, \LB_i_512\, 
        \LB_i_6[0]\, N_66, N_2573, N_2182, \LB_DOUT[0]_net_1\, 
        \REG_1_511\, N_2416_i, \REG_1_510\, \REG_1_509\, 
        \REG_1_508\, \REG_1_507\, \REG_1_506\, \REG_1_505\, 
        \REG_1_504\, \REG_1_498\, \REG_1_497\, \REG_1_496\, 
        \REG_1_495\, \REG_88[88]_net_1\, N_2159, N_2566, 
        \REG[88]\, N_20, \REG_1_494\, \REG_88[87]_net_1\, N_2158, 
        \REG[87]\, \REG_1_493\, \REG_88[86]_net_1\, N_2157, 
        \REG[86]\, \REG_1_492\, \REG_88[85]_net_1\, N_2156, 
        \REG[85]\, \REG_1_491\, \REG_88[84]_net_1\, N_2155, 
        \REG[84]\, \REG_1_490\, \REG_88[83]_net_1\, N_2154, 
        \REG[83]\, \REG_1_489\, \REG_88[82]_net_1\, N_2153, 
        \REG[82]\, \REG_1_488\, \REG_88[81]_net_1\, N_2152, 
        \REG[81]\, \STATE1[8]_net_1\, \REG_1_487\, N_3236_i, 
        \REG_1_486\, \REG[79]\, \REG_1_485\, \REG[78]\, 
        \REG_1_484\, \REG[77]\, \REG_1_483\, \REG[76]\, 
        \REG_1_482\, \REG[75]\, \REG_1_481\, \REG[74]\, 
        \REG_1_480\, \REG[73]\, \REG_1_479\, \REG[72]\, 
        \REG_1_478\, \REG[71]\, \REG_1_477\, \REG[70]\, 
        \REG_1_476\, \REG[69]\, \REG_1_475\, \REG[68]\, 
        \REG_1_474\, \REG[67]\, \REG_1_473\, \REG[66]\, 
        \REG_1_472\, \REG[65]\, \REG_1_471\, \REG[64]\, 
        \REG_1_470\, \REG[63]\, \REG_1_469\, \REG[62]\, 
        \REG_1_468\, \REG[61]\, \REG_1_467\, \REG[60]\, 
        \REG_1_466\, \REG[59]\, \REG_1_465\, \REG[58]\, 
        \REG_1_464\, \REG[57]\, N_3234_i, \REG_1_463\, \REG[56]\, 
        \REG_1_462\, \REG[55]\, \REG_1_461\, \REG[54]\, 
        \REG_1_460\, \REG[53]\, \REG_1_459\, \REG[52]\, 
        \REG_1_458\, \REG[51]\, \REG_1_457\, \REG[50]\, 
        \REG_1_456\, \REG[49]\, \REG_1_455\, \REG[48]\, N_231, 
        N_446, \REG_1_454\, \REG_1_453\, \REG_1_452\, \REG_1_451\, 
        \REG_1_450\, \REG_1_449\, \REG_1_448\, \REG_1_447\, 
        \REG_1_446\, \REG_1_445\, \REG_1_444\, \REG_1_443\, 
        \REG_1_442\, \REG_1_441\, \REG_1_440\, \REG_1_439\, 
        \REG_1_438\, \REG_1_437\, \REG_1_436\, \REG_1_435\, 
        \REG_1_434\, \REG_1_433\, \REG_1_432\, N_3170_i, 
        \REG_1_431\, \REG_1_430\, \REG_1_429\, \REG_1_428\, 
        \REG_1_427\, \REG_1_426\, \REG_1_425\, \REG_1_424\, 
        \REG_1_423\, PULSE_0_sqmuxa_1, \REG_1_422\, 
        FWIMG2LOAD_0_sqmuxa, \REG_1_421\, \REG[456]\, \REG_1_420\, 
        \REG_1_419\, \REG_1_418\, \REG_1_417\, \REG_1_416\, 
        \REG_1_415\, \REG_1_414\, \REG_1_413\, N_3104_i, 
        \REG_1_412\, \REG_1_411\, \REG[446]\, \REG_1_410\, 
        \REG[445]\, \REG_1_409\, \REG[444]\, \REG_1_408\, 
        \REG[443]\, \REG_1_407\, \REG[442]\, \REG_1_406\, 
        \REG[441]\, \REG_1_405\, \REG[440]\, \REG_1_404\, 
        \REG[439]\, \REG_1_403\, \REG[438]\, \REG_1_402\, 
        \REG[437]\, \REG_1_401\, \REG[436]\, \REG_1_400\, 
        \REG[435]\, \REG_1_399\, \REG[434]\, \REG_1_398\, 
        \REG[433]\, \REG_1_397\, \REG[432]\, \REG_1_396\, 
        \REG[431]\, \REG_1_395\, \REG[430]\, \REG_1_394\, 
        \REG[429]\, \REG_1_393\, \REG[428]\, \REG_1_392\, 
        \REG[427]\, \REG_1_391\, \REG[426]\, \REG_1_390\, 
        \REG[425]\, \REG_1_389\, \REG[424]\, \REG_1_388\, 
        \REG[423]\, \REG_1_387\, \REG[422]\, \REG_1_386\, 
        \REG[421]\, \REG_1_385\, \REG[420]\, \REG_1_384\, 
        \REG[419]\, \REG_1_383\, \REG[418]\, N_3072_i, 
        \REG_1_382\, \REG[417]\, \REG_1_381\, \REG[416]\, 
        \REG_1_380\, \REG[415]\, \REG_1_379\, \REG[414]\, 
        \REG_1_378\, \REG[413]\, \REG_1_377\, \REG[412]\, 
        \REG_1_376\, \REG[411]\, \REG_1_375\, \REG[410]\, 
        \REG_1_374\, \REG_1_373\, \REG_1_372\, \REG_1_371\, 
        \REG_1_370\, \REG_1_369\, \REG_1_368\, \REG_1_367\, 
        \REG_1_366\, \REG_1_365\, N_3008_i, \REG_1_364\, 
        \REG_1_363\, \REG_1_362\, \REG_1_361\, \REG_1_360\, 
        \REG_1_359\, \REG_1_358\, \REG_1_357\, \REG_1_356\, 
        \REG_1_355\, \REG_1_354\, \REG_1_353\, \REG_1_352\, 
        \REG_1_351\, \REG_1_350\, \REG_1_349\, \REG[384]\, 
        N_2976_i, \REG_1_348\, \REG[383]\, \REG_1_347\, 
        \REG[382]\, \REG_1_346\, \REG[381]\, \REG_1_345\, 
        \REG[380]\, \REG_1_344\, \REG[379]\, \REG_1_343\, 
        \REG[378]\, \REG_1_342\, \REG[377]\, \REG_1_341\, 
        \REG_1_340\, \REG_1_339\, \REG_1_338\, \REG_1_337\, 
        \REG_1_336\, \REG_1_335\, \REG_1_334\, \REG_1_333\, 
        \REG_1_332\, \REG_1_331\, N_2944_i, \REG_1_330\, 
        \REG_1_329\, \REG_1_328\, \REG_1_327\, \REG_1_326\, 
        \REG_1_325\, \REG_1_311\, \REG_1_310\, \REG_1_309\, 
        \REG_1_308\, \REG_1_307\, \REG_1_306\, \REG_1_305\, 
        \REG_1_304\, \REG_1_303\, \REG_1_302\, \REG_1_301\, 
        \REG_1_300\, \REG_1_299\, N_2880_i, \REG_1_298\, 
        \REG_1_297\, \REG_1_296\, \REG_1_295\, \REG_1_294\, 
        \REG_1_293\, \REG_1_279\, \REG_1_278\, \REG_1_277\, 
        \REG[264]\, \REG_1_276\, \REG[263]\, \REG_1_275\, 
        \REG[262]\, \REG_1_274\, \REG[261]\, \REG_1_273\, 
        \REG[260]\, \REG_1_272\, \REG[259]\, \REG_1_271\, 
        \REG[258]\, \REG_1_270\, \REG[257]\, \REG_1_269\, 
        \REG[256]\, N_2816_i_0, \REG_1_268\, \REG[255]\, 
        \REG_1_267\, \REG[254]\, \REG_1_266\, \REG[253]\, 
        \REG_1_265\, \REG[252]\, \REG_1_264\, \REG[251]\, 
        \REG_1_263\, \REG[250]\, \REG_1_262\, \REG[249]\, 
        \REG_1_261\, \REG[248]\, \REG_1_260\, \REG[247]\, 
        \REG_1_259\, \REG[246]\, \REG_1_258\, \REG[245]\, 
        \REG_1_257\, \REG[244]\, \REG_1_256\, \REG[243]\, 
        \REG_1_255\, \REG[242]\, \REG_1_254\, \REG[241]\, 
        \REG_1_253\, \REG[240]\, N_2784_i, \REG_1_252\, 
        \REG[239]\, \REG_1_251\, \REG[238]\, \REG_1_250\, 
        \REG[237]\, \REG_1_249\, \REG[236]\, \REG_1_248\, 
        \REG[235]\, \REG_1_247\, \REG[234]\, \REG_1_246\, 
        \REG[233]\, \PULSE_1_245\, \PULSE_42[10]\, un1_STATE1_17, 
        \PULSE[10]\, \STATE1[7]_net_1\, \PULSE_1_244\, N_2387, 
        \PULSE[9]\, \PULSE_1_243\, N_2386, \PULSE[8]\, 
        \PULSE_1_242\, N_2388, \PULSE[7]\, \REGMAP_i_0_i[11]\, 
        \PULSE_1_241\, \PULSE_42[6]\, \un1_STATE1_17_0_1\, 
        \PULSE_42_tz[6]\, \PULSE[6]\, \WRITES\, \REG_1_240\, 
        \REG[200]\, \REG_1_239\, \REG[199]\, \REG_1_238\, 
        \REG[198]\, \REG_1_237\, \REG[197]\, \REG_1_236\, 
        \REG[196]\, \REG_1_235\, \REG[195]\, \REG_1_234\, 
        \REG[194]\, \REG_1_233\, \REG[193]\, \REG_1_232\, 
        \REG[192]\, N_2752_i, \REG_1_231\, \REG[191]\, 
        \REG_1_230\, \REG[190]\, \REG_1_229\, \REG[189]\, 
        \REG_1_228\, \REG[188]\, \REG_1_227\, \REG[187]\, 
        \REG_1_226\, \REG[186]\, \REG_1_225\, \REG[185]\, 
        \REG_1_224\, \REG[184]\, \REG_1_223\, \REG[183]\, 
        \REG_1_222\, \REG[182]\, \REG_1_221\, \REG[181]\, 
        \REG_1_220\, \REG[180]\, \REG_1_219\, \REG[179]\, 
        \REG_1_218\, \REG[178]\, \REG_1_217\, \REG[177]\, 
        \REG_1_216\, \REG[176]\, N_2720_i, \REG_1_215\, 
        \REG[175]\, \REG_1_214\, \REG[174]\, \REG_1_213\, 
        \REG[173]\, \REG_1_212\, \REG[172]\, \REG_1_211\, 
        \REG[171]\, \REG_1_210\, \REG[170]\, \REG_1_209\, 
        \REG[169]\, \REG_1_208\, \REG[168]\, \REG_1_207\, 
        \REG[167]\, \REG_1_206\, \REG[166]\, \REG_1_205\, 
        \REG[165]\, \REG_1_204\, \REG[164]\, \REG_1_203\, 
        \REG[163]\, \REG_1_202\, \REG[162]\, \REG_1_201\, 
        \REG[161]\, \REG_1_200\, \REG[160]\, N_2688_i, 
        \REG_1_199\, \REG[159]\, \REG_1_198\, \REG[158]\, 
        \REG_1_197\, \REG[157]\, \REG_1_196\, \REG[156]\, 
        \REG_1_195\, \REG[155]\, \REG_1_194\, \REG[154]\, 
        \REG_1_193\, \REG[153]\, \NOEDTKi_192\, NOEDTKi_10, 
        \TST_c_c[3]\, un1_STATE1_32, \un1_STATE1_32_0_3\, 
        \un1_STATE1_32_0_2\, STATE1_tr12_7_0_o2_4_i, 
        STATE1_tr12_7_0_o2_0_i, STATE1_tr12_7_0_o2_1_i, 
        \TCNT_i_i[4]\, \TCNT[5]_net_1\, \TCNT_i_i[6]\, 
        \TCNT[7]_net_1\, STATE1_tr12_7_0_o2_2_i, \TCNT_i_i[0]\, 
        \TCNT[1]_net_1\, \TCNT_i_i[2]\, \TCNT[3]_net_1\, 
        \un1_STATE1_32_0_1\, N_2408, N_2451, \PURGED\, \TST_c[2]\, 
        un1_LB_DOUT_0_sqmuxa, un1_LB_DOUT_0_sqmuxa_0_1_i, 
        \STATE1[5]_net_1\, \OR_RDATA_191\, N_33, N_1832, 
        \OR_RDATA_190\, N_31, N_2572, \OR_RDATA_189\, N_29, 
        \OR_RDATA_188\, N_2568, \OR_RDATA_187\, N_25, 
        \OR_RDATA_186\, N_2567, \OR_RDATA_185\, N_21, 
        \OR_RDATA_184\, N_19, \OR_RDATA_183\, N_17, 
        \OR_RDATA_182\, N_13, N_1837, \EVREADi_181\, N_16, N_86, 
        \REG1_15[514]_net_1\, \RUN_c\, \REG1_1_sqmuxa\, 
        REG1_0_sqmuxa_1, \LB_DOUT_179\, \LB_DOUT_178\, 
        \LB_DOUT_177\, \LB_DOUT_176\, \LB_DOUT_175\, 
        \LB_DOUT_174\, \LB_DOUT_173\, \LB_DOUT_172\, 
        \LB_DOUT_171\, \LB_DOUT_170\, \LB_DOUT_169\, 
        \LB_DOUT_168\, \LB_DOUT_167\, \LB_DOUT_166\, 
        \LB_DOUT_165\, \LB_DOUT_164\, \LB_DOUT_163\, 
        \LB_DOUT_162\, \LB_DOUT_161\, \LB_DOUT_160\, 
        \LB_DOUT_159\, LB_DOUT_0_sqmuxa, \LB_DOUT_158\, 
        \LB_DOUT_157\, \LB_DOUT_156\, \LB_DOUT_155\, 
        \LB_DOUT_154\, \LB_DOUT_153\, \LB_DOUT_152\, 
        \LB_DOUT_151\, \LB_DOUT_150\, \LB_DOUT_149\, 
        \LB_DOUT_148\, N_2436_i, N_222_i, N_232, N_2434_1, 
        \nLBRD_146\, N_2569, N_2601_i, N_2602_i, N_2592, 
        \EVREAD_DS_145\, \TST_c_i_0[2]\, un1_EVREAD_DS_1_sqmuxa_1, 
        N_665, un1_STATE2_12_0_o2_2_i_a2_0_i, \N_77_i_i_o2_1_0\, 
        \REG_1_144\, \REG[136]\, \REG_1_143\, \REG[135]\, 
        \REG_1_142\, \REG[134]\, \REG_1_141\, \REG[133]\, 
        \REG_1_140\, \REG[132]\, \REG_1_139\, \REG[131]\, 
        \REG_1_138\, \REG[130]\, \REG_1_137\, \REG[129]\, 
        \REG_1_136\, REG_0_sqmuxa, \REG_1_131\, \REG[123]\, 
        \REG_1_130\, \REG[122]\, \REG_1_129\, \REG[121]\, 
        \REG3_128\, \REG3_127\, \REG3_126\, \REG3_125\, 
        \REG3_124\, \REG3_123\, \REG3_122\, \REG3_121\, \REG[8]\, 
        \REG3_120\, REG1_0_sqmuxa, \REG3_119\, \REG[6]\, 
        \REG3_118\, \REG3_117\, \REG3_116\, \REG3_115\, 
        \REG3_114\, \REG3_113\, \nLBLAST_112\, \STATE5_i_0[0]\, 
        N_1828, N_65, \FWIMG2LOAD_111\, \LB_s_110\, \LB_s_109\, 
        \LB_s_108\, \LB_s_107\, \LB_s_106\, \LB_s_105\, 
        \LB_s_104\, \LB_s_103\, \LB_s_102\, \LB_s_101\, 
        \LB_s_100\, \LB_s_99\, \LB_s_98\, \LB_s_97\, \LB_s_96\, 
        \LB_s_95\, \LB_s_94\, \LB_s_93\, \LB_s_92\, \LB_s_91\, 
        \LB_s_90\, \LB_s_89\, STATE5_0_sqmuxa, \LB_s_88\, 
        \LB_s_87\, \LB_s_86\, \LB_s_85\, \LB_s_84\, \LB_s_83\, 
        \LB_s_82\, \LB_s_81\, \LB_s_80\, \LB_s_79\, 
        un2_nlbrdy_i_0, \MBLTCYC_78\, \TST_c_i_0[0]\, N_2385, 
        N_2434_i, N_228, N_237, \ADACKCYC_76\, N_59, 
        \un2_vsel_1_i_a2_0\, un2_vsel_1_i_a2_1_0_i, 
        un2_vsel_1_i_a2_1_1_i, \CYCS\, \CYCS1\, \PULSE_1_75\, 
        N_2391, N_2454, \PULSE[3]\, \PULSE_1_74\, N_2390, N_2418, 
        \PULSE[2]\, \REGMAP[5]_net_1\, \PULSE_1_73\, N_2389, 
        N_2417, \PULSE[1]\, \REGMAP_i_0_i[4]\, \PULSE_1_72\, 
        N_2392, \un1_STATE1_20_i_a2_0_a2_2\, N_1698, 
        \STATE1_i_0[5]\, N_2419, \PULSE[0]\, \REGMAP_i_0_i[3]\, 
        \WDOGRES_71\, un1_WDOGRES_0_sqmuxa, 
        un1_WDOGRES_0_sqmuxa_0_a2_0_2_i, 
        un1_WDOGRES_0_sqmuxa_0_a2_0_3_i, \WDOG[5]_net_1\, 
        \un1_WDOGRES_0_sqmuxa_0_a2_0_i\, \WDOG[0]_net_1\, 
        \WDOG[3]_net_1\, \REG_1_19_70\, N_11, N_2577_i, N_2576_i, 
        un2_nlbrdy_0_a2_2_i, \LBUSTMO_i_0_i[3]\, 
        \LBUSTMO[4]_net_1\, \LBUSTMO_i_0_i[0]\, 
        \LBUSTMO_i_0_i[1]\, \LBUSTMO[2]_net_1\, \WDOGCLEAR_69\, 
        \WDOGCLEAR\, un1_STATE1_29, N_2420, \LB_WRITE_68\, 
        \LB_WRITE\, N_2384, \LB_REQ_67\, \LB_REQ\, LB_REQ_8, 
        \un1_STATE1_28_i_0\, N_2428_i, \STATE1_i_0[8]\, 
        \un1_STATE1_28_i_a2_1_0\, \VAS_66\, \VAS[15]_net_1\, 
        \VAS_65\, \VAS[14]_net_1\, \VAS_64\, \VAS[13]_net_1\, 
        \VAS_63\, \VAS[12]_net_1\, \VAS_62\, \VAS_61\, \VAS_60\, 
        \VAS_59\, \VAS_58\, \VAS_57\, \TST_c[1]\, \VAS_56\, 
        \VAS_55\, \VAS_54\, \VAS_53\, \VAS_52\, \PIPEB_51\, N_236, 
        \PIPEB_50\, \PIPEB_4[30]\, \PIPEB_49\, \PIPEB_4[29]\, 
        \PIPEB_48\, \PIPEB_4[28]\, \PIPEB_47\, N_2637, \PIPEB_46\, 
        N_2636, \PIPEB_45\, N_229, \PIPEB_44\, N_2635, \PIPEB_43\, 
        N_225, \PIPEB_42\, N_2634, \PIPEB_41\, N_2633, \PIPEB_40\, 
        N_2632, \PIPEB_39\, N_2631, \PIPEB_38\, N_199, \PIPEB_37\, 
        N_2630, \PIPEB_36\, N_186, \PIPEB_35\, N_2629, \PIPEB_34\, 
        N_2628, \PIPEB_33\, N_2627, \PIPEB_32\, N_2626, 
        \PIPEB_31\, N_2625, \PIPEB_30\, N_2624, \PIPEB_29\, 
        N_2623, N_616, \PIPEB_28\, N_2622, N_1996, \PIPEB_27\, 
        N_2621, \PIPEB_26\, N_2620, \PIPEB_25\, N_2619, 
        \PIPEB_24\, N_2618, \PIPEB_23\, N_2617, \PIPEB_22\, 
        N_2616, \PIPEB_21\, N_2615, \PIPEB_20\, N_2614, 
        \MYBERRi_19\, un1_MYBERRi_1_sqmuxa, N_2424, \TST_c[0]\, 
        \LWORDS_18\, \CYCSF1_17\, \CYCSF1\, N_2423, N_230, 
        \REG_1_24_16\, \LB_nOE_15\, un1_STATE5_8, 
        \un1_STATE5_8_0_a2_0\, \PURGED_14\, \EVREAD\, un22_bltcyc, 
        \DSSF1_13\, DSSF1_2, N_2421, \RAMAD_VME_12\, 
        \RAMAD_VME_11\, \RAMAD_VME_10\, \RAMAD_VME_9\, 
        \RAMAD_VME_8\, \RAMAD_VME_7\, \RAMAD_VME_6\, 
        \RAMAD_VME_5\, \RAMAD_VME_4\, \nLBASi_3\, \TCNT_10[7]\, 
        \N_1897\, I_34_1, \TCNT_10[6]\, N_2397, I_27, 
        \TCNT_10[5]\, I_33_1, \TCNT_10[4]\, I_28, \TCNT_10[3]\, 
        I_30_2, \TCNT_10[2]\, I_32_1, \N_1897_1\, \N_1897_0\, 
        \TCNT_10[1]\, I_31_1, \TCNT_10[0]\, 
        \DWACT_ADD_CI_0_partial_sum[0]\, \TCNT_10_0_o2_0_i[6]\, 
        N_2455, un776_regmap_25_i, un776_regmap_26_i, 
        \un776_regmap_23_0\, \REGMAP[21]_net_1\, 
        \REGMAP[22]_net_1\, un776_regmap_23_2_i, 
        un776_regmap_21_i, un776_regmap_20_i, \un776_regmap_17\, 
        \un776_regmap_13\, un776_regmap_9_i, \un776_regmap_4\, 
        un776_regmap_6_i, un776_regmap_0_i, \un776_regmap_14\, 
        \un776_regmap_19\, un776_regmap_7_i, un776_regmap_8_0_i, 
        \un7_ronly_0_a3_0_a2\, un7_ronly_0_a3_0_a2_1_i, N_658, 
        N_2369, \LBUSTMO_3[4]\, I_22_1, \LBUSTMO_3[3]\, I_21_1, 
        \LBUSTMO_3[2]\, I_20_3, \LBUSTMO_3[1]\, I_19_0, 
        \LBUSTMO_3[0]\, \DWACT_ADD_CI_0_partial_sum_0[0]\, 
        \un8_d32_0_a3_0_a2\, N_656, \un123_reg_ads_0_a2_3_a2\, 
        N_672, un84_reg_ads_1, \un120_reg_ads_0_a3_0_a2\, 
        un120_reg_ads_1, \un117_reg_ads_0_a3_0_a2\, N_684_i, 
        un98_reg_ads_1, N_690, N_674, N_716, un111_reg_ads_1, 
        \un108_reg_ads_0_a3_0_a2\, un105_reg_ads_1_0, N_683_i, 
        N_671, N_688, N_666, \un98_reg_ads_0_a3_0_a2\, N_682, 
        N_660, N_685, \un90_reg_ads_0_a3_0_a2\, 
        un90_reg_ads_0_a3_0_a2_0_i, N_673, 
        \un87_reg_ads_0_a3_0_a2\, N_675, un13_reg_ads_1, N_724, 
        N_689_i, un43_reg_ads_1, \un74_reg_ads_0_a3\, N_198, 
        \un74_reg_ads_0_a3_1\, N_463, \VAS_i_0[2]\, 
        \un70_reg_ads_0_a3_0_a2\, N_791, \un57_reg_ads_0_a3_0_a2\, 
        N_678, \un50_reg_ads_0_a2_3_a2\, \un46_reg_ads_0_a3_0_a2\, 
        N_694, N_662, \un43_reg_ads_0_a3_0_a2\, N_681_i, 
        \un40_reg_ads_0_a3_0_a2\, un33_reg_ads_1, N_667, 
        \un29_reg_ads_0_a2_0_a2\, \un25_reg_ads_0_a3_0_a2\, 
        un17_reg_ads_1, \un21_reg_ads_0_a3_0_a2\, N_664, 
        \un17_reg_ads_0_a3_0_a2\, \un10_reg_ads_0_a2_1_a2\, N_659, 
        \un2_reg_ads_0_a3_0_a2\, \un29_reg_ads_0_a2_0_a2_2_0\, 
        \un7_ronly_0_a3_0_a2_0_0\, N_2507, un12_wdog_0_a3_0_i, 
        un12_wdog_0_a3_1_i, \un10_hwres\, \un7_cycs_0_a2\, 
        \LB_ACK\, \TST_c[4]\, \NRDMEB\, \NLBRD_c\, \NLBLAST_c\, 
        FWIMG2LOAD_net_1, \MYBERR_c\, LB_nOE_net_1, \nLBAS_c\, 
        \RAMAD_VME[0]_net_1\, \RAMAD_VME[1]_net_1\, 
        \RAMAD_VME[2]_net_1\, \RAMAD_VME[3]_net_1\, 
        \RAMAD_VME[4]_net_1\, \RAMAD_VME[5]_net_1\, 
        \RAMAD_VME[6]_net_1\, \RAMAD_VME[7]_net_1\, 
        \RAMAD_VME[8]_net_1\, \REG[481]\, \REG[345]\, \REG[346]\, 
        \REG[360]\, \REG[361]\, \REG[362]\, \REG[363]\, 
        \REG[364]\, \REG[365]\, \REG[366]\, \REG[367]\, 
        \REG[368]\, \REG[369]\, \REG[370]\, \REG[371]\, 
        \REG[372]\, \REG[373]\, \REG[374]\, \REG[375]\, 
        \REG[376]\, \REG[409]\, \OR_RDATA[0]_net_1\, 
        \OR_RDATA[1]_net_1\, \OR_RDATA[2]_net_1\, 
        \OR_RDATA[3]_net_1\, \OR_RDATA[4]_net_1\, 
        \OR_RDATA[5]_net_1\, \OR_RDATA[6]_net_1\, 
        \OR_RDATA[7]_net_1\, \OR_RDATA[8]_net_1\, 
        \OR_RDATA[9]_net_1\, \LB_i[0]_net_1\, \LB_i[1]_net_1\, 
        \LB_i[2]_net_1\, \LB_i[3]_net_1\, \LB_i[4]_net_1\, 
        \LB_i[5]_net_1\, \LB_i[6]_net_1\, \LB_i[7]_net_1\, 
        \LB_i[8]_net_1\, \LB_i[9]_net_1\, \LB_i[10]_net_1\, 
        \LB_i[11]_net_1\, \LB_i[12]_net_1\, \LB_i[13]_net_1\, 
        \LB_i[14]_net_1\, \LB_i[15]_net_1\, \LB_i[16]_net_1\, 
        \LB_i[17]_net_1\, \LB_i[18]_net_1\, \LB_i[19]_net_1\, 
        \LB_i[20]_net_1\, \LB_i[21]_net_1\, \LB_i[22]_net_1\, 
        \LB_i[23]_net_1\, \LB_i[24]_net_1\, \LB_i[25]_net_1\, 
        \LB_i[26]_net_1\, \LB_i[27]_net_1\, \LB_i[28]_net_1\, 
        \LB_i[29]_net_1\, \LB_i[30]_net_1\, \LB_i[31]_net_1\, 
        \REG[89]\, \REG[90]\, \REG[91]\, \REG[97]\, \REG[98]\, 
        \REG[99]\, \REG[100]\, \REG[101]\, \REG[102]\, \REG[103]\, 
        \REG[104]\, \DWACT_ADD_CI_0_partial_sum_1[0]\, 
        \WDOG_3[1]\, \WDOG_3[2]\, \WDOG_3[3]\, \WDOG_3[4]\, 
        \WDOG_3[5]\, \DWACT_ADD_CI_0_pog_array_1_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\, 
        \DWACT_ADD_CI_0_g_array_2_0[0]\, 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_0[0]\, 
        \DWACT_ADD_CI_0_TMP_0[0]\, 
        \DWACT_ADD_CI_0_g_array_0_1[0]\, 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, 
        \DWACT_ADD_CI_0_g_array_0_3[0]\, 
        \DWACT_ADD_CI_0_partial_sum[4]\, 
        \DWACT_ADD_CI_0_partial_sum[3]\, 
        \DWACT_ADD_CI_0_partial_sum[2]\, 
        \DWACT_ADD_CI_0_partial_sum[1]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_3[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_4[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_1_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_2_0[0]\, 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_5[0]\, 
        \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_g_array_0_6[0]\, 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, 
        \DWACT_ADD_CI_0_g_array_0_2_0[0]\, 
        \DWACT_ADD_CI_0_g_array_12_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, 
        \DWACT_ADD_CI_0_g_array_0_4[0]\, 
        \DWACT_ADD_CI_0_g_array_1_2_0[0]\, 
        \DWACT_ADD_CI_0_g_array_0_5[0]\, 
        \DWACT_ADD_CI_0_g_array_1_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_0_3_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_0[0]\, 
        \DWACT_ADD_CI_0_TMP_1[0]\, 
        \DWACT_ADD_CI_0_g_array_0_1_0[0]\, 
        \DWACT_ADD_CI_0_partial_sum[7]\, 
        \DWACT_ADD_CI_0_partial_sum[5]\, 
        \DWACT_ADD_CI_0_partial_sum_0[2]\, 
        \DWACT_ADD_CI_0_partial_sum_0[1]\, 
        \DWACT_ADD_CI_0_partial_sum_0[3]\, 
        \DWACT_ADD_CI_0_partial_sum_0[4]\, 
        \DWACT_ADD_CI_0_partial_sum[6]\, \VCC\, \GND\
         : std_logic;

begin 

    RAMAD_VME(8) <= \RAMAD_VME[8]_net_1\;
    RAMAD_VME(7) <= \RAMAD_VME[7]_net_1\;
    RAMAD_VME(6) <= \RAMAD_VME[6]_net_1\;
    RAMAD_VME(5) <= \RAMAD_VME[5]_net_1\;
    RAMAD_VME(4) <= \RAMAD_VME[4]_net_1\;
    RAMAD_VME(3) <= \RAMAD_VME[3]_net_1\;
    RAMAD_VME(2) <= \RAMAD_VME[2]_net_1\;
    RAMAD_VME(1) <= \RAMAD_VME[1]_net_1\;
    RAMAD_VME(0) <= \RAMAD_VME[0]_net_1\;
    OR_RDATA(9) <= \OR_RDATA[9]_net_1\;
    OR_RDATA(8) <= \OR_RDATA[8]_net_1\;
    OR_RDATA(7) <= \OR_RDATA[7]_net_1\;
    OR_RDATA(6) <= \OR_RDATA[6]_net_1\;
    OR_RDATA(5) <= \OR_RDATA[5]_net_1\;
    OR_RDATA(4) <= \OR_RDATA[4]_net_1\;
    OR_RDATA(3) <= \OR_RDATA[3]_net_1\;
    OR_RDATA(2) <= \OR_RDATA[2]_net_1\;
    OR_RDATA(1) <= \OR_RDATA[1]_net_1\;
    OR_RDATA(0) <= \OR_RDATA[0]_net_1\;
    PULSE_0 <= \PULSE[0]\;
    PULSE_1 <= \PULSE[1]\;
    PULSE_2 <= \PULSE[2]\;
    PULSE_3 <= \PULSE[3]\;
    PULSE_6 <= \PULSE[6]\;
    PULSE_7 <= \PULSE[7]\;
    PULSE_8 <= \PULSE[8]\;
    PULSE_9 <= \PULSE[9]\;
    PULSE_10 <= \PULSE[10]\;
    LB_i(31) <= \LB_i[31]_net_1\;
    LB_i(30) <= \LB_i[30]_net_1\;
    LB_i(29) <= \LB_i[29]_net_1\;
    LB_i(28) <= \LB_i[28]_net_1\;
    LB_i(27) <= \LB_i[27]_net_1\;
    LB_i(26) <= \LB_i[26]_net_1\;
    LB_i(25) <= \LB_i[25]_net_1\;
    LB_i(24) <= \LB_i[24]_net_1\;
    LB_i(23) <= \LB_i[23]_net_1\;
    LB_i(22) <= \LB_i[22]_net_1\;
    LB_i(21) <= \LB_i[21]_net_1\;
    LB_i(20) <= \LB_i[20]_net_1\;
    LB_i(19) <= \LB_i[19]_net_1\;
    LB_i(18) <= \LB_i[18]_net_1\;
    LB_i(17) <= \LB_i[17]_net_1\;
    LB_i(16) <= \LB_i[16]_net_1\;
    LB_i(15) <= \LB_i[15]_net_1\;
    LB_i(14) <= \LB_i[14]_net_1\;
    LB_i(13) <= \LB_i[13]_net_1\;
    LB_i(12) <= \LB_i[12]_net_1\;
    LB_i(11) <= \LB_i[11]_net_1\;
    LB_i(10) <= \LB_i[10]_net_1\;
    LB_i(9) <= \LB_i[9]_net_1\;
    LB_i(8) <= \LB_i[8]_net_1\;
    LB_i(7) <= \LB_i[7]_net_1\;
    LB_i(6) <= \LB_i[6]_net_1\;
    LB_i(5) <= \LB_i[5]_net_1\;
    LB_i(4) <= \LB_i[4]_net_1\;
    LB_i(3) <= \LB_i[3]_net_1\;
    LB_i(2) <= \LB_i[2]_net_1\;
    LB_i(1) <= \LB_i[1]_net_1\;
    LB_i(0) <= \LB_i[0]_net_1\;
    REGMAP_35 <= \REGMAP[35]_net_1\;
    REGMAP_31 <= \REGMAP[31]_net_1\;
    REG_c_0 <= \REG_c[0]\;
    REG_344 <= \REG[345]\;
    REG_345 <= \REG[346]\;
    REG_359 <= \REG[360]\;
    REG_360 <= \REG[361]\;
    REG_361 <= \REG[362]\;
    REG_362 <= \REG[363]\;
    REG_363 <= \REG[364]\;
    REG_364 <= \REG[365]\;
    REG_365 <= \REG[366]\;
    REG_366 <= \REG[367]\;
    REG_367 <= \REG[368]\;
    REG_368 <= \REG[369]\;
    REG_369 <= \REG[370]\;
    REG_370 <= \REG[371]\;
    REG_371 <= \REG[372]\;
    REG_372 <= \REG[373]\;
    REG_373 <= \REG[374]\;
    REG_374 <= \REG[375]\;
    REG_375 <= \REG[376]\;
    REG_408 <= \REG[409]\;
    REG_480 <= \REG[481]\;
    REG_80 <= \REG[81]\;
    REG_81 <= \REG[82]\;
    REG_82 <= \REG[83]\;
    REG_83 <= \REG[84]\;
    REG_84 <= \REG[85]\;
    REG_85 <= \REG[86]\;
    REG_86 <= \REG[87]\;
    REG_87 <= \REG[88]\;
    REG_88 <= \REG[89]\;
    REG_89 <= \REG[90]\;
    REG_90 <= \REG[91]\;
    REG_96 <= \REG[97]\;
    REG_97 <= \REG[98]\;
    REG_98 <= \REG[99]\;
    REG_99 <= \REG[100]\;
    REG_100 <= \REG[101]\;
    REG_101 <= \REG[102]\;
    REG_102 <= \REG[103]\;
    REG_103 <= \REG[104]\;
    REG_376 <= \REG[377]\;
    REG_120 <= \REG[121]\;
    REG_152 <= \REG[153]\;
    REG_232 <= \REG[233]\;
    REG_248 <= \REG[249]\;
    REG_168 <= \REG[169]\;
    REG_184 <= \REG[185]\;
    REG_47 <= \REG[48]\;
    REG_440 <= \REG[441]\;
    REG_441 <= \REG[442]\;
    REG_121 <= \REG[122]\;
    REG_153 <= \REG[154]\;
    REG_233 <= \REG[234]\;
    REG_249 <= \REG[250]\;
    REG_169 <= \REG[170]\;
    REG_185 <= \REG[186]\;
    REG_48 <= \REG[49]\;
    REG_377 <= \REG[378]\;
    REG_409 <= \REG[410]\;
    REG_442 <= \REG[443]\;
    REG_378 <= \REG[379]\;
    REG_410 <= \REG[411]\;
    REG_154 <= \REG[155]\;
    REG_170 <= \REG[171]\;
    REG_122 <= \REG[123]\;
    REG_250 <= \REG[251]\;
    REG_186 <= \REG[187]\;
    REG_234 <= \REG[235]\;
    REG_49 <= \REG[50]\;
    REG_50 <= \REG[51]\;
    REG_155 <= \REG[156]\;
    REG_171 <= \REG[172]\;
    REG_251 <= \REG[252]\;
    REG_187 <= \REG[188]\;
    REG_235 <= \REG[236]\;
    REG_443 <= \REG[444]\;
    REG_379 <= \REG[380]\;
    REG_411 <= \REG[412]\;
    REG_51 <= \REG[52]\;
    REG_156 <= \REG[157]\;
    REG_172 <= \REG[173]\;
    REG_252 <= \REG[253]\;
    REG_188 <= \REG[189]\;
    REG_236 <= \REG[237]\;
    REG_444 <= \REG[445]\;
    REG_380 <= \REG[381]\;
    REG_412 <= \REG[413]\;
    REG_445 <= \REG[446]\;
    REG_413 <= \REG[414]\;
    REG_381 <= \REG[382]\;
    REG_52 <= \REG[53]\;
    REG_157 <= \REG[158]\;
    REG_173 <= \REG[174]\;
    REG_253 <= \REG[254]\;
    REG_189 <= \REG[190]\;
    REG_237 <= \REG[238]\;
    REG_382 <= \REG[383]\;
    REG_414 <= \REG[415]\;
    REG_5 <= \REG[6]\;
    REG_53 <= \REG[54]\;
    REG_158 <= \REG[159]\;
    REG_174 <= \REG[175]\;
    REG_254 <= \REG[255]\;
    REG_190 <= \REG[191]\;
    REG_238 <= \REG[239]\;
    REG_383 <= \REG[384]\;
    REG_415 <= \REG[416]\;
    REG_54 <= \REG[55]\;
    REG_159 <= \REG[160]\;
    REG_175 <= \REG[176]\;
    REG_255 <= \REG[256]\;
    REG_191 <= \REG[192]\;
    REG_239 <= \REG[240]\;
    REG_416 <= \REG[417]\;
    REG_7 <= \REG[8]\;
    REG_55 <= \REG[56]\;
    REG_128 <= \REG[129]\;
    REG_160 <= \REG[161]\;
    REG_240 <= \REG[241]\;
    REG_256 <= \REG[257]\;
    REG_176 <= \REG[177]\;
    REG_192 <= \REG[193]\;
    REG_56 <= \REG[57]\;
    REG_161 <= \REG[162]\;
    REG_177 <= \REG[178]\;
    REG_129 <= \REG[130]\;
    REG_257 <= \REG[258]\;
    REG_193 <= \REG[194]\;
    REG_241 <= \REG[242]\;
    REG_417 <= \REG[418]\;
    REG_57 <= \REG[58]\;
    REG_162 <= \REG[163]\;
    REG_178 <= \REG[179]\;
    REG_130 <= \REG[131]\;
    REG_258 <= \REG[259]\;
    REG_194 <= \REG[195]\;
    REG_242 <= \REG[243]\;
    REG_418 <= \REG[419]\;
    REG_58 <= \REG[59]\;
    REG_163 <= \REG[164]\;
    REG_179 <= \REG[180]\;
    REG_131 <= \REG[132]\;
    REG_259 <= \REG[260]\;
    REG_195 <= \REG[196]\;
    REG_243 <= \REG[244]\;
    REG_419 <= \REG[420]\;
    REG_59 <= \REG[60]\;
    REG_164 <= \REG[165]\;
    REG_180 <= \REG[181]\;
    REG_132 <= \REG[133]\;
    REG_260 <= \REG[261]\;
    REG_196 <= \REG[197]\;
    REG_244 <= \REG[245]\;
    REG_420 <= \REG[421]\;
    REG_60 <= \REG[61]\;
    REG_165 <= \REG[166]\;
    REG_181 <= \REG[182]\;
    REG_133 <= \REG[134]\;
    REG_261 <= \REG[262]\;
    REG_197 <= \REG[198]\;
    REG_245 <= \REG[246]\;
    REG_421 <= \REG[422]\;
    REG_61 <= \REG[62]\;
    REG_166 <= \REG[167]\;
    REG_182 <= \REG[183]\;
    REG_134 <= \REG[135]\;
    REG_262 <= \REG[263]\;
    REG_198 <= \REG[199]\;
    REG_246 <= \REG[247]\;
    REG_422 <= \REG[423]\;
    REG_455 <= \REG[456]\;
    REG_423 <= \REG[424]\;
    REG_62 <= \REG[63]\;
    REG_167 <= \REG[168]\;
    REG_183 <= \REG[184]\;
    REG_135 <= \REG[136]\;
    REG_263 <= \REG[264]\;
    REG_199 <= \REG[200]\;
    REG_247 <= \REG[248]\;
    REG_63 <= \REG[64]\;
    REG_424 <= \REG[425]\;
    REG_64 <= \REG[65]\;
    REG_425 <= \REG[426]\;
    REG_65 <= \REG[66]\;
    REG_426 <= \REG[427]\;
    REG_66 <= \REG[67]\;
    REG_427 <= \REG[428]\;
    REG_67 <= \REG[68]\;
    REG_428 <= \REG[429]\;
    REG_68 <= \REG[69]\;
    REG_429 <= \REG[430]\;
    REG_69 <= \REG[70]\;
    REG_430 <= \REG[431]\;
    REG_70 <= \REG[71]\;
    REG_431 <= \REG[432]\;
    REG_71 <= \REG[72]\;
    REG_432 <= \REG[433]\;
    REG_72 <= \REG[73]\;
    REG_433 <= \REG[434]\;
    REG_73 <= \REG[74]\;
    REG_434 <= \REG[435]\;
    REG_74 <= \REG[75]\;
    REG_435 <= \REG[436]\;
    REG_75 <= \REG[76]\;
    REG_436 <= \REG[437]\;
    REG_76 <= \REG[77]\;
    REG_437 <= \REG[438]\;
    REG_77 <= \REG[78]\;
    REG_438 <= \REG[439]\;
    REG_78 <= \REG[79]\;
    REG_439 <= \REG[440]\;
    REG_4 <= \REG[5]\;
    REG_79 <= \REG[80]\;
    TST_c_c(3) <= \TST_c_c[3]\;
    TST_c_4 <= \TST_c[4]\;
    TST_c_0 <= \TST_c[0]\;
    TST_c_5 <= \TST_c[5]\;
    TST_c_2 <= \TST_c[2]\;
    TST_c_1 <= \TST_c[1]\;
    REG_0(127) <= \REG_0[127]\;
    REG_0(126) <= \REG_0[126]\;
    REG_0(125) <= \REG_0[125]\;
    REG_0(124) <= \REG_0[124]\;
    nLBAS_c <= \nLBAS_c\;
    LB_nOE <= LB_nOE_net_1;
    MYBERR_c <= \MYBERR_c\;
    FWIMG2LOAD <= FWIMG2LOAD_net_1;
    NLBLAST_c <= \NLBLAST_c\;
    NLBRD_c <= \NLBRD_c\;
    EVREAD <= \EVREAD\;
    NRDMEB <= \NRDMEB\;
    RUN_c <= \RUN_c\;
    N_441 <= \N_441\;
    NOE16W_c <= \NOE16W_c\;
    NSELCLK_c <= \NSELCLK_c\;
    N_2613_0 <= \N_2613_0\;
    NOEAD_c_0 <= \NOEAD_c_0\;
    WDOGTO <= \WDOGTO\;
    NOEAD_c_0_0 <= \NOEAD_c_0_0\;
    RUN_c_0_0 <= \RUN_c_0_0\;

    \PIPEB_4_i[9]\ : AND2
      port map(A => DPR(9), B => N_616, Y => N_2623);
    
    \VDBi_66_0[7]\ : MUX2H
      port map(A => \REG[400]\, B => \REG[384]\, S => 
        \REGMAP[29]_net_1\, Y => N_2024);
    
    \PIPEB[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_34\, CLR => CLEAR_26, 
        Q => \PIPEB[14]_net_1\);
    
    \PIPEA1[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_577\, CLR => CLEAR_21, 
        Q => \PIPEA1[21]_net_1\);
    
    LB_s_92 : MUX2H
      port map(A => LB_in(13), B => \LB_s[13]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_92\);
    
    un4_asb_1 : XOR2FT
      port map(A => GA_c(1), B => VAD_in_28, Y => \un4_asb_1\);
    
    LB_DOUT_152 : MUX2H
      port map(A => VDB_in(4), B => \LB_DOUT[4]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_152\);
    
    \REG_1[70]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_477\, CLR => 
        \un10_hwres_30\, Q => \REG[70]\);
    
    \REG_1[281]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_294\, CLR => 
        \un10_hwres_15\, Q => \REG[281]\);
    
    PIPEB_26 : MUX2H
      port map(A => \PIPEB[6]_net_1\, B => N_2620, S => N_1996, Y
         => \PIPEB_26\);
    
    \OR_RDATA[6]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_188\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[6]_net_1\);
    
    un776_regmap_7 : OR3
      port map(A => \REGMAP[10]_net_1\, B => \REGMAP[9]_net_1\, C
         => \REGMAP_i_0_i[4]\, Y => un776_regmap_7_i);
    
    LWORDS : DFFC
      port map(CLK => CLK_c_c, D => \LWORDS_18\, CLR => 
        HWRES_c_19, Q => \LWORDS\);
    
    LB_DOUT_174 : MUX2H
      port map(A => VDB_in(26), B => \LB_DOUT[26]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_174\);
    
    REG_1_411 : MUX2H
      port map(A => VDB_in_0(5), B => \REG[446]\, S => N_3104_i, 
        Y => \REG_1_411\);
    
    WDOG_3_I_24 : XOR2
      port map(A => \WDOG_i_0_i[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => \WDOG_3[4]\);
    
    \VDBm_0[10]\ : MUX2H
      port map(A => \PIPEB[10]_net_1\, B => \PIPEA[10]_net_1\, S
         => \BLTCYC_2\, Y => N_2306);
    
    REG_1_359 : MUX2H
      port map(A => VDB_in_0(1), B => \REG[394]\, S => N_3008_i, 
        Y => \REG_1_359\);
    
    REG_0_sqmuxa_0_a3 : NOR2FT
      port map(A => \REGMAP_0[16]_net_1\, B => PULSE_0_sqmuxa_1_2, 
        Y => REG_0_sqmuxa);
    
    \LB_ADDR[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_546\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[3]_net_1\);
    
    \VDBi_92_0_iv_0[15]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[15]_net_1\, C
         => \PIPEA_m[15]_net_1\, Y => \VDBi_92_0_iv_0[15]_net_1\);
    
    REG_1_379 : MUX2H
      port map(A => VDB_in_0(5), B => \REG[414]\, S => N_3072_i, 
        Y => \REG_1_379\);
    
    REG_1_373_e_0 : OR2FT
      port map(A => \REGMAP[30]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => N_3008_i_0);
    
    un1_STATE5_18_i_0_o2 : NOR2FT
      port map(A => N_2592, B => N_66, Y => N_1837);
    
    \REG3[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_123\, CLR => 
        \un10_hwres_5\, Q => \REG[10]\);
    
    WDOG_3_I_28 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => \WDOG[1]_net_1\, 
        Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \STATE1_ns_1_iv_0_0_a2_0_1[5]\ : NAND2
      port map(A => \REGMAP[0]_net_1\, B => \STATE1[9]_net_1\, Y
         => N_573_1);
    
    \VDBi_16_1_0[3]\ : AO21TTF
      port map(A => \REGMAP[2]_net_1\, B => \REG[19]\, C => 
        N_2468, Y => \VDBi_16_1_0_i[3]\);
    
    \LB_s[14]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_93\, CLR => HWRES_c_17, 
        Q => \LB_s[14]_net_1\);
    
    \VDBi_77_d[5]\ : MUX2H
      port map(A => \REG[414]\, B => N_2057, S => \N_441\, Y => 
        \VDBi_77_d[5]_net_1\);
    
    REG_1_197 : MUX2H
      port map(A => VDB_in(4), B => \REG[157]\, S => N_2688_i, Y
         => \REG_1_197\);
    
    \PIPEA[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_613\, CLR => CLEAR_24, 
        Q => \PIPEA[24]_net_1\);
    
    LB_DOUT_173 : MUX2H
      port map(A => VDB_in(25), B => \LB_DOUT[25]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_173\);
    
    \REG_1_m[129]\ : NAND2
      port map(A => \REGMAP[16]_net_1\, B => \REG[129]\, Y => 
        \REG_1_m[129]_net_1\);
    
    \REGMAP[4]\ : DFF
      port map(CLK => CLK_c_c, D => \un21_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_0_i[4]\);
    
    LB_ADDR_547 : MUX2H
      port map(A => \LB_ADDR[4]_net_1\, B => \VAS[4]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_547\);
    
    un1_TCNT_1_I_40 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_4[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_4[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_5[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_2_0[0]\);
    
    REG_1_328 : MUX2H
      port map(A => VDB_in(18), B => \REG[363]\, S => N_2944_i, Y
         => \REG_1_328\);
    
    un102_reg_ads_0_a3_0_a2_1 : NOR2
      port map(A => \LWORDS\, B => N_659, Y => N_673);
    
    \VDBm[19]\ : MUX2H
      port map(A => N_2315, B => \VDBi[19]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_19);
    
    \PIPEA_7_i_m2[0]\ : MUX2H
      port map(A => DPR(0), B => \PIPEA1[0]_net_1\, S => N_1996_2, 
        Y => N_509);
    
    \PIPEA1_9_i[22]\ : AND2
      port map(A => DPR(22), B => N_85_3, Y => N_284);
    
    \REG_1[52]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_459\, CLR => 
        \un10_hwres_28\, Q => \REG[52]\);
    
    LB_ADDR_544 : MUX2H
      port map(A => \LB_ADDR[1]_net_1\, B => \VAS[1]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_544\);
    
    PIPEA_611 : MUX2H
      port map(A => \PIPEA_7[22]\, B => \PIPEA[22]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_611\);
    
    un1_LBUSTMO_1_I_17 : XOR2FT
      port map(A => N_66_0, B => \LBUSTMO_i_0_i[0]\, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\);
    
    \VDBi[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_626\, CLR => 
        \un10_hwres_35\, Q => \VDBi[5]_net_1\);
    
    REG_1_506 : MUX2H
      port map(A => \REG[99]\, B => VDB_in_0(10), S => N_2416_i, 
        Y => \REG_1_506\);
    
    \REG_1[197]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_237\, CLR => 
        \un10_hwres_12\, Q => \REG[197]\);
    
    \VDBi_66_0[3]\ : MUX2H
      port map(A => \REG[396]\, B => \REG[380]\, S => 
        \REGMAP[29]_net_1\, Y => N_2020);
    
    \VDBi[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_621\, CLR => 
        \un10_hwres_33\, Q => \VDBi[0]_net_1\);
    
    un11_ronlylt14_1_i_o3 : OR2
      port map(A => \VAS[13]_net_1\, B => \VAS[14]_net_1\, Y => 
        N_2369);
    
    \LB_DOUT[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_156\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[8]_net_1\);
    
    \VDBm[29]\ : MUX2H
      port map(A => N_2325, B => \VDBi[29]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_29);
    
    \VDBm_i_0_m2[21]\ : MUX2H
      port map(A => N_488, B => \VDBi[21]_net_1\, S => 
        \SINGCYC_0\, Y => N_500);
    
    \VDBi_77_0[9]\ : MUX2H
      port map(A => REG_465, B => \REG[450]\, S => 
        \REGMAP_i_i[33]\, Y => N_2061);
    
    un1_STATE2_12_0_0_1 : NAND3FFT
      port map(A => N_620_i_i, B => N_485, C => N_580, Y => 
        un1_STATE2_12_0_0_1_i);
    
    \VDBi_23_m[14]\ : AND2
      port map(A => \VDBi_9_sqmuxa_0\, B => \VDBi_23[14]_net_1\, 
        Y => \VDBi_23_m_i[14]\);
    
    \PIPEA[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_590\, CLR => CLEAR_24, 
        Q => \PIPEA[1]_net_1\);
    
    un10_hwres_32_0 : OR2
      port map(A => HWRES_c_0_0, B => WDOGTO_0, Y => 
        \un10_hwres_32_0\);
    
    \VDBi_66_0[1]\ : MUX2H
      port map(A => \REG[394]\, B => \REG[378]\, S => 
        \REGMAP[29]_net_1\, Y => N_2018);
    
    \VAS[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_62\, CLR => HWRES_c_22, 
        Q => \VAS[11]_net_1\);
    
    \VDBi_92_0_iv_0_a2_12[21]\ : NOR2
      port map(A => N_2613, B => \REGMAP_1[31]_net_1\, Y => N_669);
    
    \LB_i_6_1[14]\ : MUX2H
      port map(A => VDB_in_0(14), B => \LB_DOUT[14]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2196);
    
    REG_1_258 : MUX2H
      port map(A => VDB_in(12), B => \REG[245]\, S => N_2784_i_0, 
        Y => \REG_1_258\);
    
    REG_1_367 : MUX2H
      port map(A => VDB_in_0(9), B => \REG[402]\, S => N_3008_i_0, 
        Y => \REG_1_367\);
    
    ASBS_0 : DFFS
      port map(CLK => CLK_c_c, D => \ASBSF1\, SET => HWRES_c_13, 
        Q => \TST_c_0[0]\);
    
    \REG3[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_127\, CLR => 
        \un10_hwres_6\, Q => \REG[14]\);
    
    REG_1_278 : MUX2H
      port map(A => VDB_in(0), B => \REG[265]\, S => N_2880_i, Y
         => \REG_1_278\);
    
    REG_1_461 : MUX2H
      port map(A => VDB_in_0(6), B => \REG[54]\, S => N_3234_i, Y
         => \REG_1_461\);
    
    STATE1_tr27_i_a2 : NOR2FT
      port map(A => \WRITES_0\, B => N_2533, Y => N_2561);
    
    \STATE1[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[5]\, CLR => 
        \un10_hwres_32\, Q => \STATE1[5]_net_1\);
    
    \VDBi_60[3]\ : MUX2H
      port map(A => \VDBi_58[3]_net_1\, B => EV_RES_c, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60[3]_net_1\);
    
    un50_reg_ads_0_a2_3_a2 : NOR2FT
      port map(A => N_674, B => N_791, Y => 
        \un50_reg_ads_0_a2_3_a2\);
    
    \STATE5_0[2]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns_i_0[2]_net_1\, 
        CLR => HWRES_c_22_0, Q => \STATE5_0[2]_net_1\);
    
    \REG_1[454]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_419\, CLR => 
        \un10_hwres_25\, Q => \REG[454]\);
    
    \VDBi_60[17]\ : MUX2H
      port map(A => \VDBi_55[17]_net_1\, B => LBSP_in_17, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[17]_net_1\);
    
    un1_LBUSTMO_1_I_19 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[1]\, B => 
        \DWACT_ADD_CI_0_TMP_0[0]\, Y => I_19_0);
    
    \REG_1[369]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_334\, CLR => 
        \un10_hwres_18\, Q => \REG[369]\);
    
    REG_1_495 : MUX2H
      port map(A => \REG_88[88]_net_1\, B => \REG[88]\, S => 
        un1_STATE1_15, Y => \REG_1_495\);
    
    \REG_1[51]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_458\, CLR => 
        \un10_hwres_28\, Q => \REG[51]\);
    
    REG_1_205 : MUX2H
      port map(A => VDB_in(12), B => \REG[165]\, S => N_2688_i_0, 
        Y => \REG_1_205\);
    
    \LB_i[31]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_543\, CLR => 
        HWRES_c_16, Q => \LB_i[31]_net_1\);
    
    \LB_i_6_r[28]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_0, C => N_2210, 
        Y => \LB_i_6[28]\);
    
    \VDBi_92_0_iv_0[25]\ : OR3
      port map(A => \VDBi_92_0_iv_0_4_i[25]\, B => 
        \VDBi_92_0_iv_0_2_i[25]\, C => \VDBi_92_0_iv_0_1_i[25]\, 
        Y => \VDBi_92[25]\);
    
    \LBUSTMO[0]\ : DFFS
      port map(CLK => ALICLK_c, D => \LBUSTMO_3[0]\, SET => 
        HWRES_c_13_0, Q => \LBUSTMO_i_0_i[0]\);
    
    un1_LBUSTMO_1_I_20 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, Y => I_20_3);
    
    \REG_1[447]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_412\, CLR => 
        \un10_hwres_24\, Q => \REG[447]\);
    
    LB_i_542 : MUX2H
      port map(A => \LB_i[30]_net_1\, B => \LB_i_6[30]\, S => 
        N_2570_0, Y => \LB_i_542\);
    
    \LB_i_6_0[10]\ : AND2
      port map(A => \LB_ADDR[10]_net_1\, B => \STATE5_2[0]_net_1\, 
        Y => N_2180);
    
    \VDBm_0[6]\ : MUX2H
      port map(A => \PIPEB[6]_net_1\, B => \PIPEA[6]_net_1\, S
         => \BLTCYC\, Y => N_2302);
    
    \VDBm_0[7]\ : MUX2H
      port map(A => \PIPEB[7]_net_1\, B => \PIPEA[7]_net_1\, S
         => \BLTCYC\, Y => N_2303);
    
    \STATE2_ns_0_0_a2_0[4]\ : OR2FT
      port map(A => \STATE2[2]_net_1\, B => N_449, Y => N_725);
    
    REG_1_486 : MUX2H
      port map(A => VDB_in(31), B => \REG[79]\, S => N_3234_i_0, 
        Y => \REG_1_486\);
    
    \LB_ADDR[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_554\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[11]_net_1\);
    
    \REGMAP[15]\ : DFF
      port map(CLK => CLK_c_c, D => \un7_ronly_0_a3_0_a2\, Q => 
        \REGMAP[15]_net_1\);
    
    \PIPEA_m[22]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA[22]_net_1\, Y => 
        \PIPEA_m[22]_net_1\);
    
    \LB_ADDR[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_547\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[4]_net_1\);
    
    \VDBi_53_0_iv_2[12]\ : AOI21TTF
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[181]\, C => 
        \REG_1_m[165]_net_1\, Y => \VDBi_53_0_iv_2[12]_net_1\);
    
    REG_1_247 : MUX2H
      port map(A => VDB_in(1), B => \REG[234]\, S => N_2784_i, Y
         => \REG_1_247\);
    
    \REG_1[495]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_436\, CLR => 
        \un10_hwres_26\, Q => \REG[495]\);
    
    \LB_i_6_1[27]\ : MUX2H
      port map(A => VDB_in(27), B => \LB_DOUT[27]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2209);
    
    \VADm[21]\ : NOR2FT
      port map(A => \PIPEA[21]_net_1\, B => N_2507_0, Y => 
        VADm(21));
    
    REG_1_201 : MUX2H
      port map(A => VDB_in(8), B => \REG[161]\, S => N_2688_i_0, 
        Y => \REG_1_201\);
    
    \VDBi_77_d[15]\ : MUX2H
      port map(A => \REG[424]\, B => N_2067, S => N_441_0, Y => 
        \VDBi_77_d[15]_net_1\);
    
    VDBi_9_sqmuxa : AND3
      port map(A => \un776_regmap_23\, B => \VDBi_9_sqmuxa_1\, C
         => \VDBi_9_sqmuxa_i_1\, Y => \VDBi_9_sqmuxa\);
    
    \VDBi_92_0_iv_0[30]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[30]_net_1\, C
         => \PIPEA_m[30]_net_1\, Y => \VDBi_92_0_iv_0[30]_net_1\);
    
    \REGMAP[36]\ : DFF
      port map(CLK => CLK_c_c, D => \un8_d32_0_a3_0_a2\, Q => 
        \REGMAP[36]_net_1\);
    
    \LB_i_6_0[1]\ : AND2
      port map(A => \LB_ADDR[1]_net_1\, B => \STATE5[0]_net_1\, Y
         => N_2171);
    
    \LB_DOUT[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_169\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[21]_net_1\);
    
    un1_TCNT_1_I_34 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[7]\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => I_34_1);
    
    \PIPEA_7_r[27]\ : AND2
      port map(A => N_85_0, B => N_536, Y => \PIPEA_7[27]\);
    
    \REG_1[380]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_345\, CLR => 
        \un10_hwres_19\, Q => \REG[380]\);
    
    STATE1_tr12_7_0_o2_4 : OR3
      port map(A => STATE1_tr12_7_0_o2_2_i, B => \TCNT_i_i[0]\, C
         => \TCNT[1]_net_1\, Y => STATE1_tr12_7_0_o2_4_i);
    
    \REG_1[442]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_407\, CLR => 
        \un10_hwres_24\, Q => \REG[442]\);
    
    \VDBm[31]\ : MUX2H
      port map(A => N_2327, B => \VDBi[31]_net_1\, S => 
        \SINGCYC_0\, Y => VDBm_31);
    
    \VDBi[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_652\, CLR => 
        \un10_hwres_35\, Q => \VDBi[31]_net_1\);
    
    \PIPEA[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_602\, CLR => CLEAR_23, 
        Q => \PIPEA[13]_net_1\);
    
    \PIPEB_4_0[29]\ : OR2FT
      port map(A => N_616_0, B => DPR(29), Y => \PIPEB_4[29]\);
    
    \REG_1[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_24_16\, CLR => 
        un15_hwres_i, Q => \REG[24]\);
    
    un2_vsel_1_i_a2_0_0 : OR2
      port map(A => AMB_c(0), B => N_232, Y => 
        \un2_vsel_1_i_a2_0\);
    
    \TCNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[1]\, CLR => 
        \un10_hwres_33\, Q => \TCNT[1]_net_1\);
    
    \PIPEA1_9_i[14]\ : AND2
      port map(A => DPR(14), B => N_85_4, Y => N_268);
    
    REG_1_433 : MUX2H
      port map(A => VDB_in_0(10), B => \REG[492]\, S => 
        N_3170_i_1, Y => \REG_1_433\);
    
    \REG_1[499]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_440\, CLR => 
        \un10_hwres_27\, Q => \REG[499]\);
    
    LB_s_88 : MUX2H
      port map(A => LB_in(9), B => \LB_s[9]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_88\);
    
    un1_LBUSTMO_1_I_24 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_2[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\);
    
    un10_hwres_25 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_25\);
    
    un1_STATE2_12_0_0 : OAI21FTF
      port map(A => \STATE2[2]_net_1\, B => N_472_i_0, C => 
        un1_STATE2_12_0_0_1_i, Y => un1_STATE2_13_4);
    
    REQUESTER_1_i_0 : OA21TTF
      port map(A => N_2572_0, B => \OR_RREQ_sync\, C => N_2589, Y
         => \REQUESTER_1_i_0\);
    
    \PIPEA_7_i_m2[17]\ : MUX2H
      port map(A => DPR(17), B => \PIPEA1[17]_net_1\, S => 
        N_1996_1, Y => N_526);
    
    REG_1_405_e_1 : OR2FT
      port map(A => \REGMAP_0[31]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_3072_i_1);
    
    REG_1_454_e_0 : OR2FT
      port map(A => \REGMAP_0[13]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => N_3170_i_0);
    
    REG_1_208_e_0 : OR2FT
      port map(A => \REGMAP_0[18]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_2688_i_0);
    
    \PIPEA_7_r[9]\ : AND2
      port map(A => N_85_2, B => N_518, Y => \PIPEA_7[9]\);
    
    \LB_i_6_r[21]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_1, C => N_2203, 
        Y => \LB_i_6[21]\);
    
    un4_asb_0 : XOR2FT
      port map(A => GA_c(0), B => VAD_in_27, Y => \un4_asb_0\);
    
    un37_reg_ads_0_a2_4_a2 : NOR3
      port map(A => N_724, B => N_683_i, C => N_666, Y => 
        \un37_reg_ads_0_a2_4_a2\);
    
    REG_1_229 : MUX2H
      port map(A => VDB_in(4), B => \REG[189]\, S => N_2752_i, Y
         => \REG_1_229\);
    
    \VDBi_92_iv_0_a2_1[7]\ : NAND2
      port map(A => FBOUT(7), B => \STATE1[2]_net_1\, Y => N_596);
    
    LB_ADDR_554 : MUX2H
      port map(A => \LB_ADDR[11]_net_1\, B => \VAS[11]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_554\);
    
    un87_reg_ads_0_a3_0_a2 : NOR2FT
      port map(A => N_675, B => un13_reg_ads_1, Y => 
        \un87_reg_ads_0_a3_0_a2\);
    
    un1_TCNT_1_I_6 : AND2
      port map(A => \TCNT_i_i[2]\, B => N_83, Y => 
        \DWACT_ADD_CI_0_g_array_0_2_0[0]\);
    
    \FBOUT_m[5]\ : NAND2
      port map(A => FBOUT(5), B => \STATE1[2]_net_1\, Y => 
        \FBOUT_m[5]_net_1\);
    
    \VDBi_71[27]\ : MUX2H
      port map(A => \VDBi_60[27]_net_1\, B => \REG[436]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[27]_net_1\);
    
    \REG_1[58]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_465\, CLR => 
        \un10_hwres_29\, Q => \REG[58]\);
    
    \STATE1_ns_0_iv_0_a2_0_i[6]\ : NOR2FT
      port map(A => N_480, B => \TST_c_0[2]\, Y => N_2612);
    
    un4_asb_2 : XOR2FT
      port map(A => GA_c(2), B => VAD_in_29, Y => \un4_asb_2\);
    
    \LB_s[2]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_81\, CLR => HWRES_c_18, 
        Q => \LB_s[2]_net_1\);
    
    un1_TCNT_1_I_47 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_2_0[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\);
    
    PIPEA1_559 : MUX2H
      port map(A => N_246, B => \PIPEA1[3]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_559\);
    
    \VDBm_0[27]\ : MUX2H
      port map(A => \PIPEB[27]_net_1\, B => \PIPEA[27]_net_1\, S
         => \BLTCYC_1\, Y => N_2323);
    
    \VDBi_16_1_0[5]\ : AO21TTF
      port map(A => \REGMAP[2]_net_1\, B => REG_c_21, C => N_2474, 
        Y => \VDBi_16_1_0_i[5]\);
    
    LB_REQ_8_r : AOI21
      port map(A => \STATE1_0[8]_net_1\, B => \LB_ACK_sync\, C
         => \STATE1[10]_net_1\, Y => LB_REQ_8);
    
    REG_1_339 : MUX2H
      port map(A => VDB_in(29), B => \REG[374]\, S => N_2944_i_0, 
        Y => \REG_1_339\);
    
    \REG_1[413]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_378\, SET => 
        \un10_hwres_21\, Q => \REG[413]\);
    
    \PIPEA_m[11]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[11]_net_1\, Y => 
        \PIPEA_m[11]_net_1\);
    
    \VDBi[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_632\, CLR => 
        \un10_hwres_33\, Q => \VDBi[11]_net_1\);
    
    un1_TCNT_1_I_23 : XOR2
      port map(A => \TCNT[3]_net_1\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[3]\);
    
    \LB_DOUT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_149\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[1]_net_1\);
    
    LB_s_91 : MUX2H
      port map(A => LB_in(12), B => \LB_s[12]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_91\);
    
    \PULSE_42_f0_i_o2[1]\ : AND2
      port map(A => \REGMAP_i_0_i[4]\, B => \STATE1[8]_net_1\, Y
         => N_2417);
    
    \REG1_15[514]\ : AND2FT
      port map(A => REG1_0_sqmuxa_1, B => VDB_in(0), Y => 
        \REG1_15[514]_net_1\);
    
    \VDBi[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_634\, CLR => 
        \un10_hwres_34\, Q => \VDBi[13]_net_1\);
    
    \VDBi_92_iv_2[3]\ : AOI21TTF
      port map(A => \LB_s[3]_net_1\, B => N_7_i, C => 
        \VDBi_92_iv_1[3]_net_1\, Y => \VDBi_92_iv_2[3]_net_1\);
    
    \VDBi_53_0_iv_2[13]\ : AOI21TTF
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[182]\, C => 
        \REG_1_m[166]_net_1\, Y => \VDBi_53_0_iv_2[13]_net_1\);
    
    \PIPEA_7_r[25]\ : AND2
      port map(A => N_85_0, B => N_534, Y => \PIPEA_7[25]\);
    
    \PIPEA1_9_i[19]\ : AND2
      port map(A => DPR(19), B => N_85_4, Y => N_278);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \REG_1[234]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_247\, SET => 
        \un10_hwres_13\, Q => \REG[234]\);
    
    RAMAD_VME_12 : MUX2H
      port map(A => \VAS[9]_net_1\, B => \RAMAD_VME[8]_net_1\, S
         => N_2523_0, Y => \RAMAD_VME_12\);
    
    \LB_i_6_r[0]\ : AND3
      port map(A => N_2572_3, B => LB_i_6_sn_N_2, C => N_2182, Y
         => \LB_i_6[0]\);
    
    \VDBi[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_622\, CLR => 
        \un10_hwres_34\, Q => \VDBi[1]_net_1\);
    
    STATE1_tr25_1_0_a2_0_a2_i_o2 : OR2FT
      port map(A => \WRITES_1\, B => \REGMAP[10]_net_1\, Y => 
        N_486);
    
    \VDBi_60[0]\ : MUX2H
      port map(A => \VDBi_60_d[0]_net_1\, B => \VDBi_53[0]\, S
         => \VDBi_60_s[0]_net_1\, Y => \VDBi_60[0]_net_1\);
    
    \PIPEA1[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_570\, CLR => CLEAR_21, 
        Q => \PIPEA1[14]_net_1\);
    
    PIPEA_617 : MUX2H
      port map(A => \PIPEA_7[28]\, B => \PIPEA_i_0_i[28]\, S => 
        un1_STATE2_16_0, Y => \PIPEA_617\);
    
    \LB_i_6_r[13]\ : AND3
      port map(A => N_2572_2, B => LB_i_6_sn_N_2_1, C => N_2195, 
        Y => \LB_i_6[13]\);
    
    \PIPEB[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_43\, CLR => CLEAR_27, 
        Q => \PIPEB[23]_net_1\);
    
    un1_STATE5_8_0 : OAI21FTT
      port map(A => \STATE5_0[2]_net_1\, B => 
        \un1_STATE5_8_0_a2_0\, C => LB_i_6_sn_N_2_0, Y => 
        un1_STATE5_8);
    
    \VDBi_66[8]\ : MUX2H
      port map(A => \VDBi_60[8]_net_1\, B => N_2025, S => N_2033, 
        Y => \VDBi_66[8]_net_1\);
    
    \VDBi[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_645\, CLR => 
        \un10_hwres_35\, Q => \VDBi[24]_net_1\);
    
    un1_STATE2_8_0_0_0_o2_1 : NAND2
      port map(A => N_426, B => \STATE2_i_0[3]\, Y => N_1996_1);
    
    \REGMAP[26]\ : DFF
      port map(CLK => CLK_c_c, D => \un94_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[26]_net_1\);
    
    un776_regmap : OR3
      port map(A => N_441_0, B => un776_regmap_25_i, C => 
        un776_regmap_26_i, Y => \un776_regmap\);
    
    \VDBi_71_d[1]\ : MUX2H
      port map(A => \VDBi_66_d[1]_net_1\, B => \REG[410]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71_d[1]_net_1\);
    
    \VDBi_92_iv_2[5]\ : AOI21TTF
      port map(A => \LB_s[5]_net_1\, B => N_7_i, C => 
        \VDBi_92_iv_1[5]_net_1\, Y => \VDBi_92_iv_2[5]_net_1\);
    
    \REG_i[121]\ : INV
      port map(A => \REG[121]\, Y => REG_i_0_116);
    
    \STATE1[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[6]\, CLR => 
        \un10_hwres_32\, Q => \STATE1[4]_net_1\);
    
    REG_1_277_e : OR2FT
      port map(A => \REGMAP_0[24]_net_1\, B => PULSE_0_sqmuxa_1, 
        Y => N_2816_i_0);
    
    \PIPEA_7_i_m2[15]\ : MUX2H
      port map(A => DPR(15), B => \PIPEA1[15]_net_1\, S => 
        N_1996_1, Y => N_524);
    
    \VDBi_23_d[10]\ : MUX2H
      port map(A => \REG[58]\, B => \REG[492]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23_d[10]_net_1\);
    
    \VDBi_92_iv[4]\ : OAI21FTT
      port map(A => \VDBi_80[4]_net_1\, B => \N_2613_0\, C => 
        \VDBi_92_iv_2[4]_net_1\, Y => \VDBi_92[4]\);
    
    \VAS[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_52\, CLR => HWRES_c_22_0, 
        Q => \VAS[1]_net_1\);
    
    un1_NRDMEBi_2_sqmuxa_2_i : NOR3
      port map(A => N_7139_i, B => N_2499_i, C => 
        un1_NRDMEBi_2_sqmuxa_2_i_1_i, Y => N_42_i_0);
    
    \LB_i_6_1[16]\ : MUX2H
      port map(A => VDB_in(16), B => \LB_DOUT[16]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2198);
    
    un1_STATE2_13_i_0_o2 : OAI21
      port map(A => \STATE2[2]_net_1\, B => N_450_i, C => N_676, 
        Y => N_459);
    
    \VDBi_23_s[7]\ : OR2
      port map(A => \REGMAP_0[13]_net_1\, B => \TST_c_0[5]\, Y
         => \VDBi_23_s[7]_net_1\);
    
    \VDBi_16_r[11]\ : OA21TTF
      port map(A => N_2489_i, B => N_2488_i, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[11]\);
    
    \REG_88[85]\ : NOR2FT
      port map(A => N_2156, B => N_2566, Y => \REG_88[85]_net_1\);
    
    \PULSE_42_f0_0_a4[6]\ : NOR3FFT
      port map(A => \SINGCYC_0\, B => \STATE1_0[9]_net_1\, C => 
        N_2550_1, Y => N_2566);
    
    \PIPEA1[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_579\, CLR => CLEAR_22, 
        Q => \PIPEA1[23]_net_1\);
    
    REG_1_342 : MUX2H
      port map(A => VDB_in_0(0), B => \REG[377]\, S => N_2976_i, 
        Y => \REG_1_342\);
    
    \PIPEB_4_i_a2[0]\ : NAND2
      port map(A => N_428, B => \STATE2_i_0[3]\, Y => N_616);
    
    \LB_DOUT[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_158\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[10]_net_1\);
    
    \VDBi_80_s[2]\ : OR2
      port map(A => \REGMAP[35]_net_1\, B => N_441_0, Y => 
        \VDBi_80_s[2]_net_1\);
    
    \VDBi_21[0]\ : MUX2H
      port map(A => \VDBi_18[0]_net_1\, B => \REG[80]\, S => 
        \REGMAP[9]_net_1\, Y => \VDBi_21[0]_net_1\);
    
    REG_1_448 : MUX2H
      port map(A => VDB_in(25), B => \REG[507]\, S => N_3170_i_0, 
        Y => \REG_1_448\);
    
    \REG_m[106]\ : NAND2
      port map(A => \REGMAP[12]_net_1\, B => REG_105, Y => 
        \REG_m[106]_net_1\);
    
    \VDBi_92_0_iv_1[18]\ : AOI21TTF
      port map(A => \LB_s[18]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[18]_net_1\, Y => 
        \VDBi_92_0_iv_1[18]_net_1\);
    
    \RAMDTS[5]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(5), CLR => HWRES_c_21, 
        Q => \RAMDTS[5]_net_1\);
    
    \VDBi_53_0_iv_1[11]\ : AO21TTF
      port map(A => \REGMAP_i_i[23]\, B => \REG[244]\, C => 
        \REG_1_m[196]_net_1\, Y => \VDBi_53_0_iv_1_i[11]\);
    
    \VDBi_92_0_iv_1[29]\ : AOI21TTF
      port map(A => \LB_s[29]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[29]_net_1\, Y => 
        \VDBi_92_0_iv_1[29]_net_1\);
    
    \PIPEA_7_i_m2[5]\ : MUX2H
      port map(A => DPR(5), B => \PIPEA1[5]_net_1\, S => N_1996_2, 
        Y => N_514);
    
    REG_1_238 : MUX2H
      port map(A => VDB_in(13), B => \REG[198]\, S => N_2752_i_0, 
        Y => \REG_1_238\);
    
    REG_1_456 : MUX2H
      port map(A => VDB_in_0(1), B => \REG[49]\, S => N_3234_i, Y
         => \REG_1_456\);
    
    REG_1_346 : MUX2H
      port map(A => VDB_in_0(4), B => \REG[381]\, S => N_2976_i, 
        Y => \REG_1_346\);
    
    REG_1_309_e_0 : OR2FT
      port map(A => \REGMAP[25]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => N_2880_i_0);
    
    \PIPEA1_9_i[2]\ : AND2
      port map(A => DPR(2), B => N_85, Y => N_244);
    
    un1_STATE5_15_i : OR3
      port map(A => N_2606_i_i, B => N_2601_i, C => N_2602_i, Y
         => N_2569);
    
    REG_1_300 : MUX2H
      port map(A => VDB_in(22), B => \REG[287]\, S => N_2880_i_0, 
        Y => \REG_1_300\);
    
    REG_1_476 : MUX2H
      port map(A => VDB_in(21), B => \REG[69]\, S => N_3234_i_0, 
        Y => \REG_1_476\);
    
    un1_TCNT_1_I_12 : XOR2
      port map(A => \TCNT[1]_net_1\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_0[0]\);
    
    REG3_126 : MUX2H
      port map(A => \REG[13]\, B => VDB_in(13), S => 
        REG1_0_sqmuxa_0, Y => \REG3_126\);
    
    \VDBi_16_1_a2[14]\ : AND2
      port map(A => N_2511_0, B => REG_45, Y => N_2494_i);
    
    \LB_nOE\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_nOE_15\, CLR => 
        HWRES_c_17, Q => LB_nOE_net_1);
    
    \REG_1[381]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_346\, CLR => 
        \un10_hwres_19\, Q => \REG[381]\);
    
    REG_1_240 : MUX2H
      port map(A => VDB_in(15), B => \REG[200]\, S => N_2752_i_0, 
        Y => \REG_1_240\);
    
    \VDBi_92_iv_2[1]\ : AOI21TTF
      port map(A => \LB_s[1]_net_1\, B => N_7_i, C => 
        \VDBi_92_iv_1[1]_net_1\, Y => \VDBi_92_iv_2[1]_net_1\);
    
    \LB_i_6_1[7]\ : MUX2H
      port map(A => VDB_in_0(7), B => \LB_DOUT[7]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2189);
    
    \REGMAP[33]\ : DFF
      port map(CLK => CLK_c_c, D => \un114_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_i[33]\);
    
    REG_1_129 : MUX2H
      port map(A => \REG[121]\, B => VDB_in(0), S => REG_0_sqmuxa, 
        Y => \REG_1_129\);
    
    \VDBi_53_0_iv_3[0]\ : AO21TTF
      port map(A => \REGMAP[18]_net_1\, B => \REG[153]\, C => 
        \REG_1_m[121]_net_1\, Y => \VDBi_53_0_iv_3_i[0]\);
    
    \LB_i[7]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_519\, CLR => 
        HWRES_c_16, Q => \LB_i[7]_net_1\);
    
    \REG3[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_119\, CLR => 
        \un10_hwres_6_0\, Q => \REG[6]\);
    
    un1_STATE1_29_0 : NAND2
      port map(A => N_446, B => N_2420, Y => un1_STATE1_29);
    
    \VDBi_92_0_iv_0_a2_0[31]\ : NAND2
      port map(A => N_723, B => \REG[440]\, Y => N_610);
    
    \PIPEA_7_i[31]\ : MUX2H
      port map(A => DPR(31), B => \PIPEA1[31]_net_1\, S => 
        N_1996_0, Y => N_366);
    
    \VDBi_53_0_iv_0[11]\ : AO21TTF
      port map(A => \REGMAP[12]_net_1\, B => REG_115, C => 
        \REG_1_m[260]_net_1\, Y => \VDBi_53_0_iv_0_i[11]\);
    
    LB_DOUT_172 : MUX2H
      port map(A => VDB_in(24), B => \LB_DOUT[24]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_172\);
    
    \PIPEB[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_30\, CLR => CLEAR_26, 
        Q => \PIPEB[10]_net_1\);
    
    \LB_i_6[9]\ : MUX2H
      port map(A => N_2179, B => N_2191, S => LB_i_6_sn_N_2, Y
         => N_2225);
    
    \PIPEB_4_i[23]\ : AND2
      port map(A => DPR(23), B => N_616_0, Y => N_225);
    
    \VDBi_16_1_0[0]\ : AOI21TTF
      port map(A => EVRDY_c, B => \REGMAP[2]_net_1\, C => N_2380, 
        Y => \VDBi_16_1_0[0]_net_1\);
    
    \REG3[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_128\, CLR => 
        \un10_hwres_6\, Q => \REG[15]\);
    
    LB_s_82 : MUX2H
      port map(A => LB_in(3), B => \LB_s[3]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_82\);
    
    un10_hwres_24 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_24\);
    
    \VADm[26]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[26]_net_1\, Y => 
        VADm(26));
    
    VDBi_80_m_0_m4_0_a2 : NOR3
      port map(A => VDBi_80_m_0_m4_0_a2_1_i, B => \N_2613_0\, C
         => N_441_0, Y => \VDBi_80_m_0_m4_0_a2\);
    
    \REG_1_m[197]\ : NAND2
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[197]\, Y => 
        \REG_1_m[197]_net_1\);
    
    \REG_i[80]\ : INV
      port map(A => \REG[80]\, Y => REG_i_0_75);
    
    VDBi_651 : MUX2H
      port map(A => \VDBi_92[30]\, B => \VDBi[30]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_651\);
    
    VAS_63 : MUX2H
      port map(A => \VAS[12]_net_1\, B => VAD_in_11, S => 
        \TST_c_0[1]\, Y => \VAS_63\);
    
    \REG_1[403]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_368\, CLR => 
        \un10_hwres_20\, Q => \REG[403]\);
    
    LB_i_536 : MUX2H
      port map(A => \LB_i[24]_net_1\, B => \LB_i_6[24]\, S => 
        N_2570_0, Y => \LB_i_536\);
    
    REG_1_213 : MUX2H
      port map(A => VDB_in(4), B => \REG[173]\, S => N_2720_i, Y
         => \REG_1_213\);
    
    \STATE1_ns_0_iv_0_0[4]\ : OAI21TTF
      port map(A => N_573_1, B => N_2413, C => N_570_i, Y => 
        \STATE1_ns[4]\);
    
    REG_1_226 : MUX2H
      port map(A => VDB_in(1), B => \REG[186]\, S => N_2752_i, Y
         => \REG_1_226\);
    
    \VDBi_18[18]\ : AND2
      port map(A => \REG[66]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[18]_net_1\);
    
    \OR_RDATA_5_i[9]\ : AND2
      port map(A => N_2572_3, B => LB_in(9), Y => N_33);
    
    \REG_1[66]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_473\, CLR => 
        \un10_hwres_29\, Q => \REG[66]\);
    
    \REG_1[372]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_337\, CLR => 
        \un10_hwres_18\, Q => \REG[372]\);
    
    \REG_1[512]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_453\, SET => 
        \un10_hwres_28\, Q => \REG[512]\);
    
    \VDBi_80_d[3]\ : MUX2H
      port map(A => \VDBi_77_d[3]_net_1\, B => REG_475, S => 
        \REGMAP[35]_net_1\, Y => \VDBi_80_d[3]_net_1\);
    
    \REG_1[190]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_230\, CLR => 
        \un10_hwres_12\, Q => \REG[190]\);
    
    \PULSE_42_f0_0_tz[6]\ : OR3
      port map(A => N_2566, B => N_2430, C => \PULSE[6]\, Y => 
        \PULSE_42_tz[6]\);
    
    \PIPEA[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_609\, CLR => CLEAR_24, 
        Q => \PIPEA[20]_net_1\);
    
    un1_STATE5_14_i_0 : NAND2
      port map(A => LB_i_6_sn_N_2, B => N_2592, Y => N_1828);
    
    \PIPEA[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_605\, CLR => CLEAR_24, 
        Q => \PIPEA[16]_net_1\);
    
    \VDBi_92_0_iv[22]\ : OAI21FTT
      port map(A => \VDBi_71[22]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[22]_net_1\, Y => \VDBi_92[22]\);
    
    \REG_88_0[88]\ : MUX2H
      port map(A => VDB_in_0(7), B => \REG[88]\, S => N_20, Y => 
        N_2159);
    
    REG_1_511 : MUX2H
      port map(A => \REG[104]\, B => VDB_in_0(15), S => N_2416_i, 
        Y => \REG_1_511\);
    
    REG_1_217 : MUX2H
      port map(A => VDB_in(8), B => \REG[177]\, S => N_2720_i_0, 
        Y => \REG_1_217\);
    
    LB_DOUT_156 : MUX2H
      port map(A => VDB_in(8), B => \LB_DOUT[8]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_156\);
    
    un57_reg_ads_0_a3_0_a2 : NOR3FTT
      port map(A => \VAS[3]_net_1\, B => N_678, C => N_791, Y => 
        \un57_reg_ads_0_a3_0_a2\);
    
    un17_reg_ads_0_a3_0_a2 : NOR3
      port map(A => N_662, B => un17_reg_ads_1, C => N_671, Y => 
        \un17_reg_ads_0_a3_0_a2\);
    
    \REGMAP[30]\ : DFF
      port map(CLK => CLK_c_c, D => \un108_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[30]_net_1\);
    
    \VDBi_60[28]\ : MUX2H
      port map(A => \VDBi_55[28]_net_1\, B => LBSP_in_28, S => 
        \REGMAP_0[28]_net_1\, Y => \VDBi_60[28]_net_1\);
    
    \STATE1_ns_1_iv_0_0_a2_0_0[5]\ : OR2FT
      port map(A => \BLTCYC_0\, B => N_573_1, Y => 
        \STATE1_ns_1_iv_0_0_a2_0_0[5]_net_1\);
    
    \REG_1[376]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_341\, CLR => 
        \un10_hwres_18\, Q => \REG[376]\);
    
    \REG_1[157]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_197\, CLR => 
        \un10_hwres_9\, Q => \REG[157]\);
    
    \VDBi_92_0_iv[30]\ : OAI21FTT
      port map(A => \VDBi_71[30]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[30]_net_1\, Y => \VDBi_92[30]\);
    
    un1_STATE2_8_0_0_0_o2_2 : NAND2
      port map(A => N_426, B => \STATE2_i_0[3]\, Y => N_1996_2);
    
    \VDBi_66_d[6]\ : MUX2H
      port map(A => L1R_c_c, B => N_2023, S => N_2033, Y => 
        \VDBi_66_d[6]_net_1\);
    
    \VDBi_53_0_iv_2[7]\ : AOI21TTF
      port map(A => \REGMAP[19]_net_1\, B => \REG[176]\, C => 
        \REG_1_m[160]_net_1\, Y => \VDBi_53_0_iv_2[7]_net_1\);
    
    un4_asb_NE : NOR3
      port map(A => \un4_asb_0\, B => \un4_asb_1\, C => 
        \un4_asb_NE_0\, Y => \un4_asb_NE\);
    
    \VDBi_23_m[3]\ : AND2
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[3]_net_1\, Y
         => \VDBi_23_m_i[3]\);
    
    \REG_1[440]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_405\, CLR => 
        \un10_hwres_24\, Q => \REG[440]\);
    
    un1_TCNT_1_I_25 : XOR2
      port map(A => \TCNT[5]_net_1\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum[5]\);
    
    REG_1_388 : MUX2H
      port map(A => VDB_in_0(14), B => \REG[423]\, S => 
        N_3072_i_1, Y => \REG_1_388\);
    
    \VDBi_92_0_iv[18]\ : OAI21FTT
      port map(A => \VDBi_71[18]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[18]_net_1\, Y => \VDBi_92[18]\);
    
    PIPEB_43 : MUX2H
      port map(A => \PIPEB[23]_net_1\, B => N_225, S => N_1996_3, 
        Y => \PIPEB_43\);
    
    \VDBi_23[19]\ : MUX2H
      port map(A => \VDBi_18[19]_net_1\, B => \REG[501]\, S => 
        \REGMAP_1[13]_net_1\, Y => \VDBi_23[19]_net_1\);
    
    un776_regmap_26 : OR3
      port map(A => un776_regmap_23_2_i, B => un776_regmap_21_i, 
        C => un776_regmap_20_i, Y => un776_regmap_26_i);
    
    un2_nlbrdy_0_a2 : OR3
      port map(A => un2_nlbrdy_0_a2_2_i, B => \LBUSTMO_i_0_i[3]\, 
        C => \LBUSTMO[4]_net_1\, Y => un2_nlbrdy_i_0);
    
    \PIPEA1_9_i[16]\ : AND2
      port map(A => DPR(16), B => N_85_4, Y => N_272);
    
    \REG_1[345]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_310\, CLR => 
        \un10_hwres_17\, Q => \REG[345]\);
    
    \REGMAP[23]\ : DFF
      port map(CLK => CLK_c_c, D => \un78_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_i[23]\);
    
    \VDBi_55[3]\ : OA21TTF
      port map(A => \VDBi_23_m_i[3]\, B => \VDBi_53_0_iv_5_i[3]\, 
        C => \REGMAP[26]_net_1\, Y => \VDBi_55[3]_net_1\);
    
    \REG_i[293]\ : INV
      port map(A => \REG[293]\, Y => REG_i_0_288);
    
    LB_ADDR_0_sqmuxa_i_0_o2 : OR2FT
      port map(A => \WRITES_0\, B => N_2532, Y => N_2535);
    
    \VDBi_92_iv_2[4]\ : AOI21TTF
      port map(A => \LB_s[4]_net_1\, B => N_7_i, C => 
        \VDBi_92_iv_1[4]_net_1\, Y => \VDBi_92_iv_2[4]_net_1\);
    
    \VAS[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_57\, CLR => HWRES_c_23, 
        Q => \VAS[6]_net_1\);
    
    PIPEA_620 : MUX2H
      port map(A => \PIPEA_7[31]\, B => \PIPEA[31]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_620\);
    
    EVREAD_DS_145 : MUX2H
      port map(A => \EVREAD_DS\, B => \TST_c_i_0[2]\, S => 
        un1_EVREAD_DS_1_sqmuxa_1, Y => \EVREAD_DS_145\);
    
    REG_1_309_e : OR2FT
      port map(A => \REGMAP[25]_net_1\, B => PULSE_0_sqmuxa_1, Y
         => N_2880_i);
    
    \REGMAP_1[31]\ : DFF
      port map(CLK => CLK_c_c, D => \un111_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_1[31]_net_1\);
    
    \VDBi_16_1_0[6]\ : AO21TTF
      port map(A => \REGMAP[2]_net_1\, B => REG_c_22, C => N_2477, 
        Y => \VDBi_16_1_0_i[6]\);
    
    \LB_i_6_r[5]\ : AND2
      port map(A => N_2221, B => N_2572_3, Y => \LB_i_6[5]_net_1\);
    
    \VDBi_53_0_iv_2[14]\ : AOI21TTF
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[183]\, C => 
        \REG_1_m[167]_net_1\, Y => \VDBi_53_0_iv_2[14]_net_1\);
    
    \VDBi_18[30]\ : NAND2
      port map(A => \REG[78]\, B => \TST_c_0[5]\, Y => 
        \VDBi_18[30]_net_1\);
    
    un117_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_684_i, B => un98_reg_ads_1, Y => 
        \un117_reg_ads_0_a3_0_a2\);
    
    CYCS : DFFC
      port map(CLK => CLK_c_c, D => \CYCSF1\, CLR => HWRES_c_13, 
        Q => \CYCS\);
    
    PIPEA1_562 : MUX2H
      port map(A => N_252, B => \PIPEA1[6]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_562\);
    
    \PIPEA_m[9]\ : NAND2
      port map(A => N_457_i_0, B => \PIPEA[9]_net_1\, Y => 
        \PIPEA_m[9]_net_1\);
    
    \PIPEA1[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_567\, CLR => CLEAR_20, 
        Q => \PIPEA1[11]_net_1\);
    
    \VDBi_92_0_iv_0[19]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[19]_net_1\, C
         => \PIPEA_m[19]_net_1\, Y => \VDBi_92_0_iv_0[19]_net_1\);
    
    REG_1_301 : MUX2H
      port map(A => VDB_in(23), B => \REG[288]\, S => N_2880_i_0, 
        Y => \REG_1_301\);
    
    \VDBi_55[30]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[30]_net_1\, Y => \VDBi_55[30]_net_1\);
    
    \PIPEA_7_s[30]\ : OR2FT
      port map(A => N_85_0, B => N_539, Y => \PIPEA_7[30]\);
    
    VAS_54 : MUX2H
      port map(A => \VAS[3]_net_1\, B => VAD_in_2, S => 
        \TST_c[1]\, Y => \VAS_54\);
    
    PIPEB_46 : MUX2H
      port map(A => \PIPEB[26]_net_1\, B => N_2636, S => N_1996_3, 
        Y => \PIPEB_46\);
    
    REG_1_263 : MUX2H
      port map(A => VDB_in(1), B => \REG[250]\, S => N_2816_i_0, 
        Y => \REG_1_263\);
    
    \RAMAD_VME[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_4\, CLR => 
        \un10_hwres_4\, Q => \RAMAD_VME[0]_net_1\);
    
    \VDBi_92_0_iv_0_a2_2[31]\ : NAND2
      port map(A => N_793, B => \REG[513]\, Y => N_612);
    
    \PIPEA_7_i_m2[22]\ : MUX2H
      port map(A => DPR(22), B => \PIPEA1[22]_net_1\, S => 
        N_1996_0, Y => N_531);
    
    \REG3[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_125\, CLR => 
        \un10_hwres_6\, Q => \REG[12]\);
    
    \PIPEB[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_46\, CLR => CLEAR_27, 
        Q => \PIPEB[26]_net_1\);
    
    \VADm[4]\ : NOR2FT
      port map(A => \PIPEA[4]_net_1\, B => N_2507_0, Y => VADm(4));
    
    REG3_122 : MUX2H
      port map(A => \REG[9]\, B => VDB_in(9), S => 
        REG1_0_sqmuxa_0, Y => \REG3_122\);
    
    \LB_i_6_r[15]\ : AND3
      port map(A => N_2572_2, B => LB_i_6_sn_N_2_1, C => N_2197, 
        Y => \LB_i_6[15]\);
    
    VDBi_642 : MUX2H
      port map(A => \VDBi_92[21]\, B => \VDBi[21]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_642\);
    
    \PIPEA_m[24]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA[24]_net_1\, Y => 
        \PIPEA_m[24]_net_1\);
    
    REG_1_509 : MUX2H
      port map(A => \REG[102]\, B => VDB_in_0(13), S => N_2416_i, 
        Y => \REG_1_509\);
    
    un1_TCNT_1_I_11 : AND2
      port map(A => \TCNT[3]_net_1\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_3_0[0]\);
    
    \REG_1[433]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_398\, CLR => 
        \un10_hwres_23\, Q => \REG[433]\);
    
    \PIPEA_7_i_m2[13]\ : MUX2H
      port map(A => DPR(13), B => \PIPEA1[13]_net_1\, S => 
        N_1996_1, Y => N_522);
    
    \REG_1[455]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_420\, CLR => 
        \un10_hwres_25\, Q => \REG[455]\);
    
    OR_RDATA_187 : MUX2H
      port map(A => N_25, B => \OR_RDATA[5]_net_1\, S => N_1832, 
        Y => \OR_RDATA_187\);
    
    REG_1_267 : MUX2H
      port map(A => VDB_in(5), B => \REG[254]\, S => N_2816_i_0, 
        Y => \REG_1_267\);
    
    PIPEA_602 : MUX2H
      port map(A => \PIPEA_7[13]\, B => \PIPEA[13]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_602\);
    
    \PIPEA_m[18]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[18]_net_1\, Y => 
        \PIPEA_m[18]_net_1\);
    
    REG_1_344 : MUX2H
      port map(A => VDB_in_0(2), B => \REG[379]\, S => N_2976_i, 
        Y => \REG_1_344\);
    
    un1_STATE5_10_i : OAI21FTT
      port map(A => \LB_WRITE_sync\, B => N_66, C => N_2603, Y
         => N_2570);
    
    LB_DOUT_159 : MUX2H
      port map(A => VDB_in(11), B => \LB_DOUT[11]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_159\);
    
    PULSE_1_75 : MUX2H
      port map(A => \PULSE[3]\, B => N_2391, S => N_2454, Y => 
        \PULSE_1_75\);
    
    \LB_i_6[11]\ : MUX2H
      port map(A => N_2181, B => N_2193, S => LB_i_6_sn_N_2_1, Y
         => N_2227);
    
    \VDBi_77_s[3]\ : NOR2
      port map(A => \N_441\, B => \VDBi_71_s[4]_net_1\, Y => 
        \VDBi_77_s[3]_net_1\);
    
    \VDBi_16_1_a2_0[14]\ : AND2
      port map(A => N_2512_0, B => \REG[14]\, Y => N_2495_i);
    
    \STATE5_ns_0_0_a2_3[1]\ : NOR2
      port map(A => \STATE5[1]_net_1\, B => \STATE5[2]_net_1\, Y
         => N_2607);
    
    \REGMAP_0[23]\ : DFF
      port map(CLK => CLK_c_c, D => \un78_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_i_0[23]\);
    
    \LB_i[22]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_534\, CLR => 
        HWRES_c_15, Q => \LB_i[22]_net_1\);
    
    un8_d32_0_a3_0_a2_0 : OR2
      port map(A => N_2369, B => \VAS[15]_net_1\, Y => N_656);
    
    \REG_1[162]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_202\, CLR => 
        \un10_hwres_9\, Q => \REG[162]\);
    
    \REG_i[395]\ : INV
      port map(A => \REG[395]\, Y => REG_i_0_390);
    
    REG_1_447 : MUX2H
      port map(A => VDB_in(24), B => \REG[506]\, S => N_3170_i_0, 
        Y => \REG_1_447\);
    
    \PIPEA_7_r[24]\ : AND2
      port map(A => N_85_1, B => N_533, Y => \PIPEA_7[24]\);
    
    REG_1_424 : MUX2H
      port map(A => VDB_in_0(1), B => \REG[483]\, S => N_3170_i, 
        Y => \REG_1_424\);
    
    \REGMAP[20]\ : DFF
      port map(CLK => CLK_c_c, D => \un67_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[20]_net_1\);
    
    PIPEA_591 : MUX2H
      port map(A => \PIPEA_7[2]\, B => \PIPEA[2]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_591\);
    
    \REG_1[164]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_204\, CLR => 
        \un10_hwres_9\, Q => \REG[164]\);
    
    \VDBm_0[18]\ : MUX2H
      port map(A => \PIPEB[18]_net_1\, B => \PIPEA[18]_net_1\, S
         => \BLTCYC_2\, Y => N_2314);
    
    \VDBi_92_0_iv_0[11]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[11]_net_1\, C
         => \PIPEA_m[11]_net_1\, Y => \VDBi_92_0_iv_0[11]_net_1\);
    
    \LB_i_6_1[2]\ : MUX2H
      port map(A => VDB_in_0(2), B => \LB_DOUT[2]_net_1\, S => 
        \STATE5[0]_net_1\, Y => N_2184);
    
    \LB_i[20]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_532\, CLR => 
        HWRES_c_15, Q => \LB_i[20]_net_1\);
    
    REG_1_436 : MUX2H
      port map(A => VDB_in_0(13), B => \REG[495]\, S => 
        N_3170_i_1, Y => \REG_1_436\);
    
    \REGMAP_0[8]\ : DFF
      port map(CLK => CLK_c_c, D => \un37_reg_ads_0_a2_4_a2\, Q
         => \TST_c_0[5]\);
    
    \VDBi_53_0_iv_2[10]\ : AOI21TTF
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[179]\, C => 
        \REG_1_m[163]_net_1\, Y => \VDBi_53_0_iv_2[10]_net_1\);
    
    PIPEA_593 : MUX2H
      port map(A => \PIPEA_7[4]\, B => \PIPEA[4]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_593\);
    
    N_2522_i_i_o2_0 : AND3
      port map(A => N_425, B => \STATE1_0[9]_net_1\, C => 
        \REGMAP[0]_net_1\, Y => N_457_i_0_0);
    
    \REG_1[166]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_206\, CLR => 
        \un10_hwres_10\, Q => \REG[166]\);
    
    \REG3[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_122\, CLR => 
        \un10_hwres_7\, Q => \REG[9]\);
    
    \REG_1[502]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_443\, SET => 
        \un10_hwres_27\, Q => \REG[502]\);
    
    \TCNT_10_0_a2[0]\ : AND2
      port map(A => N_2397, B => \DWACT_ADD_CI_0_partial_sum[0]\, 
        Y => \TCNT_10[0]\);
    
    un1_STATE1_17_0 : OR3FFT
      port map(A => \un1_STATE1_17_0_1\, B => N_446, C => 
        \STATE1_0[1]_net_1\, Y => un1_STATE1_17);
    
    \REG_1_m[192]\ : NAND2
      port map(A => \REGMAP[20]_net_1\, B => \REG[192]\, Y => 
        \REG_1_m[192]_net_1\);
    
    \VDBi_53_0_iv_0[7]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_143, C => 
        \REG_1_m[256]_net_1\, Y => \VDBi_53_0_iv_0_i[7]\);
    
    un46_reg_ads_0_a3_0_a2 : NOR3
      port map(A => N_689_i, B => N_694, C => \VAS[3]_net_1\, Y
         => \un46_reg_ads_0_a3_0_a2\);
    
    N_7_i_0_a2 : NOR2FT
      port map(A => \STATE1[9]_net_1\, B => N_425, Y => N_7_i);
    
    LB_DOUT_150 : MUX2H
      port map(A => VDB_in(2), B => \LB_DOUT[2]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_150\);
    
    \REG_1[383]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_348\, CLR => 
        \un10_hwres_19\, Q => \REG[383]\);
    
    \VDBi_66[12]\ : MUX2H
      port map(A => \VDBi_66_d[12]_net_1\, B => 
        \VDBi_58[12]_net_1\, S => \VDBi_66_s[1]_net_1\, Y => 
        \VDBi_66[12]_net_1\);
    
    un1_STATE5_8_0_a2_0 : OR2
      port map(A => \STATE5[1]_net_1\, B => \LB_WRITE_sync\, Y
         => \un1_STATE5_8_0_a2_0\);
    
    LB_s_106 : MUX2H
      port map(A => LB_in(27), B => \LB_s[27]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_106\);
    
    \LB_i_6_1[22]\ : MUX2H
      port map(A => VDB_in(22), B => \LB_DOUT[22]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2204);
    
    REG_1_418 : MUX2H
      port map(A => VDB_in_0(12), B => \REG[453]\, S => 
        N_3104_i_0, Y => \REG_1_418\);
    
    REG_1_442 : MUX2H
      port map(A => VDB_in(19), B => \REG[501]\, S => N_3170_i_1, 
        Y => \REG_1_442\);
    
    REG_1_295 : MUX2H
      port map(A => VDB_in(17), B => \REG[282]\, S => N_2880_i, Y
         => \REG_1_295\);
    
    CYCSF1_17_i : INV
      port map(A => \TST_c[0]\, Y => \TST_c_i_0[0]\);
    
    REG_1_240_e : OR2FT
      port map(A => \REGMAP_0[20]_net_1\, B => PULSE_0_sqmuxa_1_2, 
        Y => N_2752_i);
    
    \REG_1[91]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_498\, CLR => 
        \un10_hwres_31\, Q => \REG[91]\);
    
    \VDBi_53_0_iv[2]\ : AO21TTF
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[2]_net_1\, C
         => \VDBi_53_0_iv_5[2]_net_1\, Y => \VDBi_53[2]\);
    
    \VDBi_16_1_a2_0[1]\ : AND2
      port map(A => N_2511, B => REG_32, Y => N_2461_i);
    
    \VDBi_71[13]\ : MUX2H
      port map(A => \VDBi_66[13]_net_1\, B => \REG[422]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71[13]_net_1\);
    
    \VDBi_66_0[15]\ : MUX2H
      port map(A => \REG[408]\, B => \REG[392]\, S => 
        \REGMAP_0[29]_net_1\, Y => N_2032);
    
    \REG_i[286]\ : INV
      port map(A => \REG[286]\, Y => REG_i_0_281);
    
    LB_s_90 : MUX2H
      port map(A => LB_in(11), B => \LB_s[11]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_90\);
    
    \VDBi_92_0_iv_0[29]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[29]_net_1\, C
         => \PIPEA_m[29]_net_1\, Y => \VDBi_92_0_iv_0[29]_net_1\);
    
    OR_RDATA_188 : MUX2H
      port map(A => N_2568, B => \OR_RDATA[6]_net_1\, S => N_1832, 
        Y => \OR_RDATA_188\);
    
    END_PK_1_0_i_a2_0_a2_4 : NAND2
      port map(A => \EVREAD_DS\, B => \STATE2[1]_net_1\, Y => 
        N_85_4);
    
    un84_reg_ads_0_a3_0_a2_1 : NAND2
      port map(A => N_682, B => N_690, Y => un84_reg_ads_1);
    
    \WDOG[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \WDOG_3[1]\, CLR => 
        un15_hwres_i, Q => \WDOG[1]_net_1\);
    
    \PULSE_42_f0_0[6]\ : NOR3FFT
      port map(A => N_2524, B => \PULSE_42_tz[6]\, C => 
        \STATE1_0[7]_net_1\, Y => \PULSE_42[6]\);
    
    WDOG_3_I_26 : XOR2
      port map(A => \WDOG[5]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => \WDOG_3[5]\);
    
    \REG_1[416]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_381\, CLR => 
        \un10_hwres_22\, Q => \REG[416]\);
    
    \PULSE_1[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_244\, CLR => 
        \un10_hwres_4\, Q => \PULSE[9]\);
    
    REG_1_210 : MUX2H
      port map(A => VDB_in(1), B => \REG[170]\, S => N_2720_i, Y
         => \REG_1_210\);
    
    \VDBi_53_0_iv_0[8]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_144, C => 
        \REG_m[113]_net_1\, Y => \VDBi_53_0_iv_0_i[8]\);
    
    PIPEA1_583 : MUX2H
      port map(A => N_294, B => \PIPEA1[27]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_583\);
    
    \REGMAP_0[13]\ : DFF
      port map(CLK => CLK_c_c, D => \un84_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[13]_net_1\);
    
    \LB_i_6_1[17]\ : MUX2H
      port map(A => VDB_in(17), B => \LB_DOUT[17]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2199);
    
    \VDBi_92_0_iv_0_a2_5[25]\ : NAND2
      port map(A => \LB_s[25]_net_1\, B => N_7_i_0, Y => N_608);
    
    \REG_1[421]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_386\, CLR => 
        \un10_hwres_22\, Q => \REG[421]\);
    
    \VDBi_92_iv_2[6]\ : AOI21TTF
      port map(A => \LB_s[6]_net_1\, B => N_7_i, C => 
        \VDBi_92_iv_1[6]_net_1\, Y => \VDBi_92_iv_2[6]_net_1\);
    
    \VDBi_92_0_iv_0_a2_9[21]\ : NOR3FTT
      port map(A => \TST_c_0[5]\, B => \REGMAP_0[13]_net_1\, C
         => N_680, Y => N_790);
    
    \VDBi_53_0_iv_1[15]\ : AO21TTF
      port map(A => \REGMAP_i_i[23]\, B => \REG[248]\, C => 
        \REG_1_m[200]_net_1\, Y => \VDBi_53_0_iv_1_i[15]\);
    
    \REG_1[295]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_308\, CLR => 
        \un10_hwres_17\, Q => \REG[295]\);
    
    VDBi_66_sn_m1 : OR2
      port map(A => \REGMAP_0[29]_net_1\, B => \REGMAP[30]_net_1\, 
        Y => N_2033);
    
    \STATE1_ns_0_iv_0_a2_0_1[9]\ : OR2FT
      port map(A => \un776_regmap\, B => \REGMAP[36]_net_1\, Y
         => N_2552_1);
    
    \VDBi_77_0[14]\ : MUX2H
      port map(A => REG_470, B => \REG[455]\, S => 
        \REGMAP_i_i[33]\, Y => N_2066);
    
    NRDMEBi_588 : MUX2H
      port map(A => \NRDMEB\, B => N_42_i_0, S => 
        \un1_NRDMEBi_2_sqmuxa_1_i_a3_i\, Y => \NRDMEBi_588\);
    
    LB_s_81 : MUX2H
      port map(A => LB_in(2), B => \LB_s[2]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_81\);
    
    REG_1_358 : MUX2H
      port map(A => VDB_in_0(0), B => \REG[393]\, S => N_3008_i, 
        Y => \REG_1_358\);
    
    \REG_1[374]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_339\, CLR => 
        \un10_hwres_18\, Q => \REG[374]\);
    
    WDOG_3_I_15 : XOR2
      port map(A => \WDOG[0]_net_1\, B => TICK(2), Y => 
        \DWACT_ADD_CI_0_partial_sum_1[0]\);
    
    \REG_i[510]\ : INV
      port map(A => \REG[510]\, Y => \REG_i[510]_net_1\);
    
    \VDBm_0[30]\ : MUX2H
      port map(A => \PIPEB[30]_net_1\, B => \PIPEA[30]_net_1\, S
         => \BLTCYC_0\, Y => N_2326);
    
    \REG_i[499]\ : INV
      port map(A => \REG[499]\, Y => \REG_i[499]_net_1\);
    
    \REG_i[393]\ : INV
      port map(A => \REG[393]\, Y => REG_i_0_388);
    
    REG_1_378 : MUX2H
      port map(A => VDB_in_0(4), B => \REG[413]\, S => N_3072_i, 
        Y => \REG_1_378\);
    
    \PIPEA[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_606\, CLR => CLEAR_24, 
        Q => \PIPEA[17]_net_1\);
    
    \VDBi_92_0_iv_0_a2_13[21]\ : OR3FTT
      port map(A => N_669, B => \REGMAP_0[26]_net_1\, C => 
        \REGMAP_0[28]_net_1\, Y => N_680);
    
    \VDBm_0[25]\ : MUX2H
      port map(A => \PIPEB[25]_net_1\, B => \PIPEA[25]_net_1\, S
         => \BLTCYC_1\, Y => N_2321);
    
    \VDBm_i_m2[11]\ : MUX2H
      port map(A => N_2540, B => \VDBi[11]_net_1\, S => 
        \SINGCYC_0\, Y => VDBm_i_m2(11));
    
    un1_LBUSTMO_1_I_22 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\, Y => I_22_1);
    
    \REG_1[238]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_251\, SET => 
        \un10_hwres_13\, Q => \REG[238]\);
    
    \PIPEA1[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_561\, CLR => CLEAR_23, 
        Q => \PIPEA1[5]_net_1\);
    
    \VDBi_53_0_iv_5[1]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[1]\, B => \REG_1_m_i[234]\, 
        C => \REG_1_m_i[250]\, Y => \VDBi_53_0_iv_5_i[1]\);
    
    \TCNT_10_0_o2_0[6]\ : OAI21
      port map(A => PULSE_0_sqmuxa_1_1, B => \REGMAP[10]_net_1\, 
        C => N_2455, Y => \TCNT_10_0_o2_0_i[6]\);
    
    MBLTCYC : DFFC
      port map(CLK => CLK_c_c, D => \MBLTCYC_78\, CLR => 
        HWRES_c_19, Q => \MBLTCYC\);
    
    \REG_1[291]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_304\, CLR => 
        \un10_hwres_16\, Q => \REG[291]\);
    
    \VDBi_92_iv[5]\ : OAI21FTT
      port map(A => \VDBi_80[5]_net_1\, B => \N_2613_0\, C => 
        \VDBi_92_iv_2[5]_net_1\, Y => \VDBi_92[5]\);
    
    \VAS[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_55\, CLR => HWRES_c_22_0, 
        Q => \VAS[4]_net_1\);
    
    \VDBi_53_0_iv_5[8]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[8]\, B => \REG_1_m_i[241]\, 
        C => \REG_1_m_i[257]\, Y => \VDBi_53_0_iv_5_i[8]\);
    
    \VDBi_53_0_iv_5[2]\ : NOR3
      port map(A => \VDBi_53_0_iv_3_i[2]\, B => 
        \VDBi_53_0_iv_0_i[2]\, C => \VDBi_53_0_iv_1_i[2]\, Y => 
        \VDBi_53_0_iv_5[2]_net_1\);
    
    REG_1_132 : MUX2H
      port map(A => \REG_0[124]\, B => VDB_in(3), S => 
        REG_0_sqmuxa, Y => \REG_1_132\);
    
    un12_wdog_0_a3_1 : NAND2
      port map(A => \WDOG[0]_net_1\, B => \WDOG[3]_net_1\, Y => 
        un12_wdog_0_a3_1_i);
    
    REG_1_362 : MUX2H
      port map(A => VDB_in_0(4), B => \REG[397]\, S => N_3008_i, 
        Y => \REG_1_362\);
    
    un1_TCNT_1_I_28 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum_0[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, Y => I_28);
    
    un1_STATE1_4_i_a2_0_o2_i_o2 : NOR2
      port map(A => \STATE1[2]_net_1\, B => \STATE1[3]_net_1\, Y
         => N_2524);
    
    PIPEA_594 : MUX2H
      port map(A => \PIPEA_7[5]\, B => \PIPEA[5]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_594\);
    
    \VDBi_53_0_iv_0[15]\ : AO21TTF
      port map(A => \REGMAP[12]_net_1\, B => REG_119, C => 
        \REG_1_m[264]_net_1\, Y => \VDBi_53_0_iv_0_i[15]\);
    
    \VDBi_18[20]\ : NAND2
      port map(A => \REG[68]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[20]_net_1\);
    
    \VDBi_71[29]\ : MUX2H
      port map(A => \VDBi_60[29]_net_1\, B => \REG[438]\, S => 
        \REGMAP_0[31]_net_1\, Y => \VDBi_71[29]_net_1\);
    
    REG_1_134 : MUX2H
      port map(A => \REG_0[126]\, B => VDB_in(5), S => 
        REG_0_sqmuxa, Y => \REG_1_134\);
    
    REG_1_468 : MUX2H
      port map(A => VDB_in_0(13), B => \REG[61]\, S => N_3234_i_1, 
        Y => \REG_1_468\);
    
    \VDBi_53_0_iv_1[7]\ : AO21TTF
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[240]\, C => 
        \REG_1_m[192]_net_1\, Y => \VDBi_53_0_iv_1_i[7]\);
    
    un1_MYBERRi_1_sqmuxa_0 : AO21TTF
      port map(A => N_2612, B => \PURGED\, C => N_2424, Y => 
        un1_MYBERRi_1_sqmuxa);
    
    \PIPEB_4_0[28]\ : OR2FT
      port map(A => N_616_0, B => DPR(28), Y => \PIPEB_4[28]\);
    
    \TCNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[2]\, CLR => 
        \un10_hwres_33\, Q => \TCNT_i_i[2]\);
    
    \VDBi_58[7]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[7]\, B => \VDBi_23_m_i[7]\, 
        C => \VDBi_58_0[9]\, Y => \VDBi_58[7]_net_1\);
    
    \OR_RDATA_5_i_o2_1[0]\ : OR2
      port map(A => N_66_0, B => \STATE5_0[2]_net_1\, Y => 
        N_2572_1);
    
    \TCNT[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[7]\, CLR => 
        \un10_hwres_33\, Q => \TCNT[7]_net_1\);
    
    REG_1_136 : MUX2H
      port map(A => \REG[128]\, B => VDB_in(7), S => REG_0_sqmuxa, 
        Y => \REG_1_136\);
    
    \VDBi_60[20]\ : MUX2H
      port map(A => \VDBi_55[20]_net_1\, B => LBSP_in_20, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[20]_net_1\);
    
    REG_1_366 : MUX2H
      port map(A => VDB_in_0(8), B => \REG[401]\, S => N_3008_i_0, 
        Y => \REG_1_366\);
    
    \VDBi_23_m[15]\ : AND2
      port map(A => \VDBi_9_sqmuxa_0\, B => \VDBi_23[15]_net_1\, 
        Y => \VDBi_23_m_i[15]\);
    
    \VDBi[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_630\, CLR => 
        \un10_hwres\, Q => \VDBi[9]_net_1\);
    
    un1_STATE2_12_0_o2_2_i_a2_0 : NOR2
      port map(A => \PIPEB[29]_net_1\, B => \PIPEB[31]_net_1\, Y
         => un1_STATE2_12_0_o2_2_i_a2_0_i);
    
    \REG_1[98]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_505\, CLR => 
        \un10_hwres_31\, Q => \REG[98]\);
    
    \LB_s[22]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_101\, CLR => 
        HWRES_c_18, Q => \LB_s[22]_net_1\);
    
    \VDBi_77_d[4]\ : MUX2H
      port map(A => \VDBi_71_d[4]_net_1\, B => N_2056, S => 
        \N_441\, Y => \VDBi_77_d[4]_net_1\);
    
    \PULSE_42_f0_i[9]\ : OA21FTF
      port map(A => N_2816_i_0_0, B => \PULSE[9]\, C => 
        \STATE1[7]_net_1\, Y => N_2387);
    
    \STATE5[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns[0]\, CLR => 
        HWRES_c_21_0, Q => \STATE5[0]_net_1\);
    
    LB_s_96 : MUX2H
      port map(A => LB_in(17), B => \LB_s[17]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_96\);
    
    TCNT_0_sqmuxa_i_s_0 : OR3FFT
      port map(A => \REGMAP[15]_net_1\, B => \WRITES_0\, C => 
        N_1898, Y => N_2523_0);
    
    REG_1_260 : MUX2H
      port map(A => VDB_in(14), B => \REG[247]\, S => N_2784_i_0, 
        Y => \REG_1_260\);
    
    LB_i_522 : MUX2H
      port map(A => \LB_i[10]_net_1\, B => \LB_i_6[10]_net_1\, S
         => N_2570_1, Y => \LB_i_522\);
    
    N_7_i_0_a2_0 : NOR2FT
      port map(A => \STATE1_0[9]_net_1\, B => N_425, Y => N_7_i_0);
    
    \VDBi_71[16]\ : MUX2H
      port map(A => \VDBi_60[16]_net_1\, B => \REG[425]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[16]_net_1\);
    
    \REG_1[59]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_466\, CLR => 
        \un10_hwres_29\, Q => \REG[59]\);
    
    un1_STATE1_17_0_1 : NOR3FFT
      port map(A => \STATE1_i_0[5]\, B => N_462, C => 
        \STATE1[0]_net_1\, Y => \un1_STATE1_17_0_1\);
    
    \VDBm[0]\ : MUX2H
      port map(A => N_2296, B => \VDBi[0]_net_1\, S => \SINGCYC\, 
        Y => VDBm_0);
    
    \LB_s[20]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_99\, CLR => HWRES_c_18, 
        Q => \LB_s[20]_net_1\);
    
    \REG_1[387]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_352\, CLR => 
        \un10_hwres_19\, Q => \REG[387]\);
    
    PIPEA1_572 : MUX2H
      port map(A => N_272, B => \PIPEA1[16]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_572\);
    
    \REG_1[244]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_257\, SET => 
        \un10_hwres_13\, Q => \REG[244]\);
    
    \VDBi_53_0_iv_1[3]\ : AO21TTF
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[236]\, C => 
        \REG_1_m[188]_net_1\, Y => \VDBi_53_0_iv_1_i[3]\);
    
    \STATE2_ns_0_0[3]\ : OAI21
      port map(A => \EVREAD_DS\, B => N_426, C => 
        \STATE2_ns_0_0_0[3]_net_1\, Y => \STATE2_ns[3]\);
    
    \REG_1[242]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_255\, SET => 
        \un10_hwres_13\, Q => \REG[242]\);
    
    un1_STATE1_15_0_i2_0_a2_i_o2 : NAND2
      port map(A => \STATE1[8]_net_1\, B => \WRITES\, Y => N_446);
    
    \PIPEB[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_47\, CLR => CLEAR_27, 
        Q => \PIPEB[27]_net_1\);
    
    \REG_1[481]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_422\, CLR => 
        \un10_hwres_25\, Q => \REG[481]\);
    
    \REG_1[123]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_131\, CLR => 
        \un10_hwres_7_0\, Q => \REG[123]\);
    
    \VDBi_66_0[8]\ : MUX2H
      port map(A => \REG[401]\, B => \NSELCLK_c\, S => 
        \REGMAP[29]_net_1\, Y => N_2025);
    
    REG_1_303 : MUX2H
      port map(A => VDB_in(25), B => \REG[290]\, S => N_2880_i_0, 
        Y => \REG_1_303\);
    
    \REG_1[368]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_333\, CLR => 
        \un10_hwres_18\, Q => \REG[368]\);
    
    \VDBi_23[13]\ : MUX2H
      port map(A => \VDBi_16[13]\, B => \VDBi_23_d[13]_net_1\, S
         => \VDBi_23_s[7]_net_1\, Y => \VDBi_23[13]_net_1\);
    
    un10_hwres_15 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_15\);
    
    un1_STATE2_10_i_0 : OAI21FTF
      port map(A => \STATE2[1]_net_1\, B => \STATE2[2]_net_1\, C
         => N_86, Y => N_16);
    
    \PULSE_1[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_73\, CLR => 
        \un10_hwres_4\, Q => \PULSE[1]\);
    
    un1_TCNT_1_I_9 : AND2
      port map(A => \TCNT[5]_net_1\, B => N_83, Y => 
        \DWACT_ADD_CI_0_g_array_0_5[0]\);
    
    \PIPEA[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_598\, CLR => CLEAR_26, 
        Q => \PIPEA[9]_net_1\);
    
    \VDBi_71_s[4]\ : OR2
      port map(A => \REGMAP_0[31]_net_1\, B => N_2033_0, Y => 
        \VDBi_71_s[4]_net_1\);
    
    \VDBi_92_0_iv_0_a2_5[31]\ : NAND2
      port map(A => \LB_s[31]_net_1\, B => N_7_i_0, Y => N_615);
    
    \VDBi_66[13]\ : MUX2H
      port map(A => \VDBi_60[13]_net_1\, B => N_2030, S => 
        N_2033_0, Y => \VDBi_66[13]_net_1\);
    
    un1_STATE2_16_0_0_0 : OAI21FTF
      port map(A => \STATE2[5]_net_1\, B => DTEST_FIFO, C => 
        \STATE2[2]_net_1\, Y => un1_STATE2_16_0_0_0_i);
    
    \REG_1[406]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_371\, CLR => 
        \un10_hwres_21\, Q => \REG[406]\);
    
    \REG_1[175]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_215\, CLR => 
        \un10_hwres_10\, Q => \REG[175]\);
    
    \VAS[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_63\, CLR => HWRES_c_22, 
        Q => \VAS[12]_net_1\);
    
    un1_LBUSTMO_1_I_13 : XOR2FT
      port map(A => N_66, B => \LBUSTMO[4]_net_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[4]\);
    
    \PIPEA_m[30]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA[30]_net_1\, Y => 
        \PIPEA_m[30]_net_1\);
    
    \PIPEA_m[29]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA[29]_net_1\, Y => 
        \PIPEA_m[29]_net_1\);
    
    \LB_i_6[5]\ : MUX2H
      port map(A => N_2175, B => N_2187, S => LB_i_6_sn_N_2, Y
         => N_2221);
    
    \VDBm_0[2]\ : MUX2H
      port map(A => \PIPEB[2]_net_1\, B => \PIPEA[2]_net_1\, S
         => \BLTCYC\, Y => N_2298);
    
    REQUESTER : DFFC
      port map(CLK => ALICLK_c, D => \REQUESTER_1_i_0\, CLR => 
        HWRES_c_21, Q => \REQUESTER\);
    
    \VDBi[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_642\, CLR => 
        \un10_hwres_34\, Q => \VDBi[21]_net_1\);
    
    \PIPEA1[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_569\, CLR => CLEAR_21, 
        Q => \PIPEA1[13]_net_1\);
    
    \REG_1[505]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_446\, CLR => 
        \un10_hwres_27\, Q => \REG[505]\);
    
    \LB_s[9]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_88\, CLR => HWRES_c_19, 
        Q => \LB_s[9]_net_1\);
    
    \VADm[11]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[11]_net_1\, Y => VADm(11));
    
    REG_1_390 : MUX2H
      port map(A => VDB_in(16), B => \REG[425]\, S => N_3072_i_1, 
        Y => \REG_1_390\);
    
    LB_DOUT_176 : MUX2H
      port map(A => VDB_in(28), B => \LB_DOUT[28]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_176\);
    
    PIPEA1_558 : MUX2H
      port map(A => N_244, B => \PIPEA1[2]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_558\);
    
    \PIPEA1[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_587\, CLR => CLEAR_22, 
        Q => \PIPEA1[31]_net_1\);
    
    VDBi_626 : MUX2H
      port map(A => \VDBi_92[5]\, B => \VDBi[5]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_626\);
    
    \VDBi_58[14]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[14]\, B => 
        \VDBi_23_m_i[14]\, C => \VDBi_58_0[9]\, Y => 
        \VDBi_58[14]_net_1\);
    
    \VDBi[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_644\, CLR => 
        \un10_hwres_34\, Q => \VDBi[23]_net_1\);
    
    \VDBi_92_0_iv_1[15]\ : AOI21TTF
      port map(A => \LB_s[15]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[15]_net_1\, Y => 
        \VDBi_92_0_iv_1[15]_net_1\);
    
    REG_1_259 : MUX2H
      port map(A => VDB_in(13), B => \REG[246]\, S => N_2784_i_0, 
        Y => \REG_1_259\);
    
    PULSE_1_72 : MUX2H
      port map(A => \PULSE[0]\, B => N_2392, S => N_2454, Y => 
        \PULSE_1_72\);
    
    \REG_1_m[195]\ : NAND2
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[195]\, Y => 
        \REG_1_m[195]_net_1\);
    
    \VDBi_80_d[1]\ : MUX2H
      port map(A => N_2053, B => REG_473, S => \REGMAP[35]_net_1\, 
        Y => \VDBi_80_d[1]_net_1\);
    
    \LB_DOUT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_151\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[3]_net_1\);
    
    REG_1_279 : MUX2H
      port map(A => VDB_in(1), B => \REG[266]\, S => N_2880_i, Y
         => \REG_1_279\);
    
    un1_anycyc_i_0_o2_i_a2 : OR2
      port map(A => \SINGCYC_0\, B => \BLTCYC_0\, Y => N_2507);
    
    \VDBi_92_0_iv_0_0[21]\ : OR3
      port map(A => \VDBi_92_0_iv_0_0_4_i[21]\, B => 
        \VDBi_92_0_iv_0_0_2_i[21]\, C => 
        \VDBi_92_0_iv_0_0_1_i[21]\, Y => \VDBi_92[21]\);
    
    REG_1_417 : MUX2H
      port map(A => VDB_in_0(11), B => \REG[452]\, S => 
        N_3104_i_0, Y => \REG_1_417\);
    
    PIPEA1_566 : MUX2H
      port map(A => N_260, B => \PIPEA1[10]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_566\);
    
    \REG3[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_117\, CLR => 
        \un10_hwres_6_0\, Q => \REG[4]\);
    
    RAMAD_VME_5 : MUX2H
      port map(A => \VAS[2]_net_1\, B => \RAMAD_VME[1]_net_1\, S
         => \TCNT_0_sqmuxa_i_s\, Y => \RAMAD_VME_5\);
    
    \VDBi_55[4]\ : OA21TTF
      port map(A => \VDBi_23_m_i[4]\, B => \VDBi_53_0_iv_5_i[4]\, 
        C => \REGMAP[26]_net_1\, Y => \VDBi_55[4]_net_1\);
    
    \VDBi_18[23]\ : NAND2
      port map(A => \REG[71]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[23]_net_1\);
    
    END_PK : DFFC
      port map(CLK => CLK_c_c, D => \END_PK_555\, CLR => CLEAR_20, 
        Q => \END_PK\);
    
    \REG_1[390]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_355\, CLR => 
        \un10_hwres_19\, Q => \REG[390]\);
    
    \VDBi_92_0_iv_0_a2_10[21]\ : AND2
      port map(A => N_669, B => \REGMAP_1[28]_net_1\, Y => N_792);
    
    \VDBi_53_0_iv_0[0]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_136, C => 
        \REG_m[105]_net_1\, Y => \VDBi_53_0_iv_0_i[0]\);
    
    \OR_RDATA_5_i[5]\ : AND2
      port map(A => N_2572, B => LB_in(5), Y => N_25);
    
    \REG_1[183]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_223\, CLR => 
        \un10_hwres_11\, Q => \REG[183]\);
    
    \VDBi_92_0_iv_0_1[12]\ : AOI21TTF
      port map(A => \LB_s[12]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0_0[12]_net_1\, Y => 
        \VDBi_92_0_iv_0_1[12]_net_1\);
    
    un1_STATE2_16_0_0_2 : NAND3FTT
      port map(A => un1_STATE2_16_0_0_0_i, B => N_79, C => N_580, 
        Y => un1_STATE2_16_1);
    
    \PULSE_42_f0_i_o2[2]\ : AND2
      port map(A => \REGMAP[5]_net_1\, B => \STATE1[8]_net_1\, Y
         => N_2418);
    
    BLTCYC_1 : DFFC
      port map(CLK => CLK_c_c, D => \BLTCYC_77\, CLR => 
        HWRES_c_13_0, Q => \BLTCYC_1\);
    
    un22_bltcyc_0_a2_0_a2 : OR2
      port map(A => \MBLTCYC\, B => \BLTCYC_0\, Y => un22_bltcyc);
    
    \TCNT_10_0_o2[6]\ : OAI21FTF
      port map(A => PULSE_0_sqmuxa_1_2, B => \LB_ADDR_0_sqmuxa_1\, 
        C => \TCNT_10_0_o2_0_i[6]\, Y => N_2397);
    
    \VDBi_23[8]\ : MUX2H
      port map(A => \VDBi_18[8]_net_1\, B => \REG[490]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23[8]_net_1\);
    
    \REG_1[168]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_208\, CLR => 
        \un10_hwres_10\, Q => \REG[168]\);
    
    \VDBm[16]\ : MUX2H
      port map(A => N_2312, B => \VDBi[16]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_16);
    
    END_PK_1_0_i_a2_0_a2_2 : NAND2
      port map(A => \EVREAD_DS\, B => \STATE2[1]_net_1\, Y => 
        N_85_2);
    
    REG_1_440 : MUX2H
      port map(A => VDB_in(17), B => \REG[499]\, S => N_3170_i_1, 
        Y => \REG_1_440\);
    
    \REG_1[510]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_451\, SET => 
        \un10_hwres_28\, Q => \REG[510]\);
    
    REG_1_338 : MUX2H
      port map(A => VDB_in(28), B => \REG[373]\, S => N_2944_i_0, 
        Y => \REG_1_338\);
    
    REG_1_412 : MUX2H
      port map(A => VDB_in_0(6), B => \REG[447]\, S => N_3104_i, 
        Y => \REG_1_412\);
    
    \REG_1_m[187]\ : NAND2
      port map(A => \REGMAP[20]_net_1\, B => \REG[187]\, Y => 
        \REG_1_m[187]_net_1\);
    
    \VDBm[4]\ : MUX2H
      port map(A => N_2300, B => \VDBi[4]_net_1\, S => \SINGCYC\, 
        Y => VDBm_4);
    
    \REG_1[57]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_464\, CLR => 
        \un10_hwres_28\, Q => \REG[57]\);
    
    \PIPEA_7_r[31]\ : AND2
      port map(A => N_85_0, B => N_366, Y => \PIPEA_7[31]\);
    
    un1_STATE2_8_0_0_0_o2_3 : NAND2
      port map(A => N_426, B => \STATE2_i_0[3]\, Y => N_1996_3);
    
    REG_1_345 : MUX2H
      port map(A => VDB_in_0(3), B => \REG[380]\, S => N_2976_i, 
        Y => \REG_1_345\);
    
    \PIPEA_7_i_m2[27]\ : MUX2H
      port map(A => DPR(27), B => \PIPEA1[27]_net_1\, S => 
        N_1996_0, Y => N_536);
    
    WDOG_3_I_33 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    \VDBi_77_0[15]\ : MUX2H
      port map(A => REG_471, B => \REG[456]\, S => 
        \REGMAP_i_i[33]\, Y => N_2067);
    
    un3_noe32wi_i_s_0 : OR2
      port map(A => \LWORDS\, B => \NOE16W_c\, Y => NOE32W_c);
    
    PIPEA1_587 : MUX2H
      port map(A => N_296, B => \PIPEA1[31]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_587\);
    
    \LB_i_6_r[29]\ : AND3
      port map(A => N_2572_0, B => LB_i_6_sn_N_2_0, C => N_2211, 
        Y => \LB_i_6[29]\);
    
    REG_1_307 : MUX2H
      port map(A => VDB_in(29), B => \REG[294]\, S => N_2880_i_0, 
        Y => \REG_1_307\);
    
    \REG_1[102]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_509\, CLR => 
        \un10_hwres_7\, Q => \REG[102]\);
    
    \OR_RDATA[3]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_185\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[3]_net_1\);
    
    \STATE1_ns_0_iv_0[9]\ : OAI21TTF
      port map(A => N_2552_1, B => 
        \STATE1_ns_0_iv_0_a2_0_1[9]_net_1\, C => N_2551_i, Y => 
        \STATE1_ns[9]\);
    
    PIPEB_22 : MUX2H
      port map(A => \PIPEB[2]_net_1\, B => N_2616, S => N_1996, Y
         => \PIPEB_22\);
    
    \LB_DOUT[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_172\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[24]_net_1\);
    
    \VDBm_0[0]\ : MUX2H
      port map(A => \PIPEB[0]_net_1\, B => \PIPEA[0]_net_1\, S
         => \BLTCYC\, Y => N_2296);
    
    \REG_1[436]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_401\, CLR => 
        \un10_hwres_23\, Q => \REG[436]\);
    
    DSS_0 : DFFS
      port map(CLK => CLK_c_c, D => \DSSF1\, SET => HWRES_c_0, Q
         => \TST_c_0[2]\);
    
    \VDBm[26]\ : MUX2H
      port map(A => N_2322, B => \VDBi[26]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_26);
    
    REG_1_401 : MUX2H
      port map(A => VDB_in(27), B => \REG[436]\, S => N_3072_i_0, 
        Y => \REG_1_401\);
    
    \REG_1[104]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_511\, CLR => 
        \un10_hwres_7\, Q => \REG[104]\);
    
    \REGMAP[29]\ : DFF
      port map(CLK => CLK_c_c, D => \un105_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[29]_net_1\);
    
    LB_DOUT_161 : MUX2H
      port map(A => VDB_in(13), B => \LB_DOUT[13]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_161\);
    
    REG_1_364 : MUX2H
      port map(A => VDB_in_0(6), B => \REG[399]\, S => N_3008_i, 
        Y => \REG_1_364\);
    
    \PULSE_1[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_75\, CLR => 
        \un10_hwres_4\, Q => \PULSE[3]\);
    
    \VDBi_66_0[13]\ : MUX2H
      port map(A => \REG[406]\, B => \REG[390]\, S => 
        \REGMAP_0[29]_net_1\, Y => N_2030);
    
    LB_s_79 : MUX2H
      port map(A => LB_in(0), B => \LB_s[0]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_79\);
    
    LB_DOUT_179 : MUX2H
      port map(A => VDB_in(31), B => \LB_DOUT[31]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_179\);
    
    \RAMAD_VME[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_9\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[5]_net_1\);
    
    \VDBm[9]\ : MUX2H
      port map(A => N_2305, B => \VDBi[9]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_9);
    
    LB_REQ_67 : MUX2H
      port map(A => \LB_REQ\, B => LB_REQ_8, S => N_2384, Y => 
        \LB_REQ_67\);
    
    \REGMAP_0[26]\ : DFF
      port map(CLK => CLK_c_c, D => \un94_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[26]_net_1\);
    
    \PULSE_42_f0_i[2]\ : OA21TTF
      port map(A => N_2418, B => \PULSE[2]\, C => 
        \STATE1[7]_net_1\, Y => N_2390);
    
    un1_STATE5_10_i_0 : OAI21FTT
      port map(A => \LB_WRITE_sync\, B => N_66_0, C => N_2603, Y
         => N_2570_0);
    
    REG_1_467 : MUX2H
      port map(A => VDB_in_0(12), B => \REG[60]\, S => N_3234_i_1, 
        Y => \REG_1_467\);
    
    ASBSF1 : DFFS
      port map(CLK => CLK_c_c, D => ASB_c, SET => HWRES_c_13, Q
         => \ASBSF1\);
    
    VDBi_9_sqmuxa_i_0 : NOR2
      port map(A => \REGMAP_i_i[23]\, B => \REGMAP[24]_net_1\, Y
         => \VDBi_9_sqmuxa_i_0\);
    
    \LBUSTMO_3_0[4]\ : OR2FT
      port map(A => N_2572_0, B => I_22_1, Y => \LBUSTMO_3[4]\);
    
    un10_hwres_14 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_14\);
    
    un111_reg_ads_0_a3_0_a2_1 : OR2FT
      port map(A => N_688, B => N_666, Y => un111_reg_ads_1);
    
    REG3_117 : MUX2H
      port map(A => \REG[4]\, B => VDB_in(4), S => REG1_0_sqmuxa, 
        Y => \REG3_117\);
    
    \VDBi_77[11]\ : MUX2H
      port map(A => \VDBi_71[11]_net_1\, B => N_2063, S => 
        N_441_0, Y => \VDBi_77[11]_net_1\);
    
    \REG_1_m[257]\ : AND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[257]\, Y => 
        \REG_1_m_i[257]\);
    
    \VDBi_58_0[7]\ : NOR2
      port map(A => \REGMAP[26]_net_1\, B => \REGMAP[27]_net_1\, 
        Y => \VDBi_58_0[9]\);
    
    \PIPEB_4_i[11]\ : AND2
      port map(A => DPR(11), B => N_616_1, Y => N_2625);
    
    LWORDS_18 : MUX2H
      port map(A => \LWORDS\, B => LWORDB_in, S => \TST_c[1]\, Y
         => \LWORDS_18\);
    
    un1_REG_0_sqmuxa_i : OR3
      port map(A => N_66, B => N_2577_i, C => N_2576_i, Y => N_11);
    
    \REG_1_m[252]\ : NAND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[252]\, Y => 
        \REG_1_m[252]_net_1\);
    
    \LB_DOUT[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_179\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[31]_net_1\);
    
    \VDBi_23_m[10]\ : AND2
      port map(A => \VDBi_9_sqmuxa_0\, B => \VDBi_23[10]_net_1\, 
        Y => \VDBi_23_m_i[10]\);
    
    WRITES_2 : MUX2H
      port map(A => \WRITES\, B => WRITEB_c, S => \TST_c[1]\, Y
         => \WRITES_2\);
    
    un1_REG_0_sqmuxa_i_o2_0 : OR2
      port map(A => \STATE5_0[0]_net_1\, B => \STATE5[1]_net_1\, 
        Y => N_66_0);
    
    \OR_RDATA_5_i_o2[0]\ : OR2
      port map(A => N_66_0, B => \STATE5_0[2]_net_1\, Y => N_2572);
    
    un776_regmap_6 : OR3
      port map(A => un776_regmap_0_i, B => \REGMAP_i_0_i[3]\, C
         => \REGMAP[5]_net_1\, Y => un776_regmap_6_i);
    
    LB_DOUT_170 : MUX2H
      port map(A => VDB_in(22), B => \LB_DOUT[22]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_170\);
    
    REG_1_484 : MUX2H
      port map(A => VDB_in(29), B => \REG[77]\, S => N_3234_i_0, 
        Y => \REG_1_484\);
    
    \VDBi_53_0_iv_0[6]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_142, C => 
        \REG_1_m[255]_net_1\, Y => \VDBi_53_0_iv_0_i[6]\);
    
    un111_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_716, B => un111_reg_ads_1, Y => 
        \un111_reg_ads_0_a3_0_a2\);
    
    \PIPEA_7_i_m2[25]\ : MUX2H
      port map(A => DPR(25), B => \PIPEA1[25]_net_1\, S => 
        N_1996_0, Y => N_534);
    
    \VDBi_23[9]\ : MUX2H
      port map(A => \VDBi_16[9]\, B => \VDBi_23_d[9]_net_1\, S
         => \VDBi_23_s[7]_net_1\, Y => \VDBi_23[9]_net_1\);
    
    REG_1_425 : MUX2H
      port map(A => VDB_in_0(2), B => \REG[484]\, S => N_3170_i, 
        Y => \REG_1_425\);
    
    \REG_88[82]\ : NOR2FT
      port map(A => N_2153, B => N_2566, Y => \REG_88[82]_net_1\);
    
    \STATE1_ns_1_iv_0_a2_2_i_o2[5]\ : NOR2FT
      port map(A => \STATE1[5]_net_1\, B => \TST_c[0]\, Y => 
        N_480);
    
    REG_1_462 : MUX2H
      port map(A => VDB_in_0(7), B => \REG[55]\, S => N_3234_i, Y
         => \REG_1_462\);
    
    \PIPEA1[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_583\, CLR => CLEAR_22, 
        Q => \PIPEA1[27]_net_1\);
    
    \STATE2[3]\ : DFFS
      port map(CLK => CLK_c_c, D => \STATE2_i[4]_net_1\, SET => 
        CLEAR, Q => \STATE2_i_0[3]\);
    
    \VDBi_92_iv_0[1]\ : AOI21TTF
      port map(A => \RAMDTS[1]_net_1\, B => \STATE1[1]_net_1\, C
         => \FBOUT_m[1]_net_1\, Y => \VDBi_92_iv_0[1]_net_1\);
    
    REG_1_391 : MUX2H
      port map(A => VDB_in(17), B => \REG[426]\, S => N_3072_i_1, 
        Y => \REG_1_391\);
    
    NOEDTKi : DFFS
      port map(CLK => CLK_c_c, D => \NOEDTKi_192\, SET => 
        \un10_hwres_4\, Q => \TST_c_c[3]\);
    
    LB_i_512 : MUX2H
      port map(A => \LB_i[0]_net_1\, B => \LB_i_6[0]\, S => 
        N_2570, Y => \LB_i_512\);
    
    un1_EVREAD_DS_1_sqmuxa_1_0_a2_2_a2_0 : AND2
      port map(A => \MBLTCYC\, B => N_652, Y => N_665);
    
    \VDBi_53_0_iv_5[7]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[7]\, B => 
        \VDBi_53_0_iv_0_i[7]\, C => \VDBi_53_0_iv_1_i[7]\, Y => 
        \VDBi_53_0_iv_5_i[7]\);
    
    VDBi_644 : MUX2H
      port map(A => \VDBi_92[23]\, B => \VDBi[23]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_644\);
    
    \TCNT_10_0_a2_1_0_a2[6]\ : OR2
      port map(A => N_486, B => N_1898, Y => N_2455_1);
    
    \REG_i[508]\ : INV
      port map(A => \REG[508]\, Y => \REG_i[508]_net_1\);
    
    \VDBm_0[26]\ : MUX2H
      port map(A => \PIPEB[26]_net_1\, B => \PIPEA[26]_net_1\, S
         => \BLTCYC_1\, Y => N_2322);
    
    \PIPEA1[28]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEA1_584\, SET => CLEAR_22, 
        Q => \PIPEA1[28]_net_1\);
    
    VDBi_649 : MUX2H
      port map(A => \VDBi_92[28]\, B => \VDBi[28]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_649\);
    
    \VDBm[8]\ : MUX2H
      port map(A => N_2304, B => \VDBi[8]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_8);
    
    \PULSE_42_f0_i[1]\ : OA21TTF
      port map(A => N_2417, B => \PULSE[1]\, C => 
        \STATE1[7]_net_1\, Y => N_2389);
    
    \VDBm_0[1]\ : MUX2H
      port map(A => \PIPEB[1]_net_1\, B => \PIPEA[1]_net_1\, S
         => \BLTCYC\, Y => N_2297);
    
    \REG_1_m[163]\ : NAND2
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[163]\, Y => 
        \REG_1_m[163]_net_1\);
    
    \REG_1[513]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_454\, CLR => 
        \un10_hwres_28\, Q => \REG[513]\);
    
    \REG_1[375]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_340\, CLR => 
        \un10_hwres_18\, Q => \REG[375]\);
    
    \PIPEB_4_i[4]\ : AND2
      port map(A => DPR(4), B => N_616, Y => N_2618);
    
    LB_s_80 : MUX2H
      port map(A => LB_in(1), B => \LB_s[1]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_80\);
    
    un43_reg_ads_0_a3_0_a2_1 : NAND2
      port map(A => N_463, B => \VAS[1]_net_1\, Y => 
        un43_reg_ads_1);
    
    \VDBi_53_0_iv_5[6]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[6]\, B => 
        \VDBi_53_0_iv_0_i[6]\, C => \VDBi_53_0_iv_1_i[6]\, Y => 
        \VDBi_53_0_iv_5_i[6]\);
    
    REG_1_138 : MUX2H
      port map(A => \REG[130]\, B => VDB_in(9), S => 
        REG_0_sqmuxa_0, Y => \REG_1_138\);
    
    \REG_1[443]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_408\, CLR => 
        \un10_hwres_24\, Q => \REG[443]\);
    
    \REGMAP_0[16]\ : DFF
      port map(CLK => CLK_c_c, D => \un54_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[16]_net_1\);
    
    REG_1_373_e : OR2FT
      port map(A => \REGMAP[30]_net_1\, B => PULSE_0_sqmuxa_1, Y
         => N_3008_i);
    
    LB_s_97 : MUX2H
      port map(A => LB_in(18), B => \LB_s[18]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_97\);
    
    \VDBi_60_s[0]\ : NOR2FT
      port map(A => \VDBi_58_0[9]\, B => \REGMAP_0[28]_net_1\, Y
         => \VDBi_60_s[0]_net_1\);
    
    \VDBi[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_629\, CLR => 
        \un10_hwres\, Q => \VDBi[8]_net_1\);
    
    \REG_i[280]\ : INV
      port map(A => \REG[280]\, Y => REG_i_0_275);
    
    LB_DOUT_168 : MUX2H
      port map(A => VDB_in(20), B => \LB_DOUT[20]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_168\);
    
    un29_reg_ads_0_a2_0_a2_2 : OR3
      port map(A => N_658, B => N_656, C => 
        \un29_reg_ads_0_a2_0_a2_2_0\, Y => N_659);
    
    REG_1_429 : MUX2H
      port map(A => VDB_in_0(6), B => \REG[488]\, S => N_3170_i, 
        Y => \REG_1_429\);
    
    \REG_1[255]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_268\, CLR => 
        \un10_hwres_14\, Q => \REG[255]\);
    
    REG_1_256 : MUX2H
      port map(A => VDB_in(10), B => \REG[243]\, S => N_2784_i_0, 
        Y => \REG_1_256\);
    
    un776_regmap_14_i_0_o2_0 : OR2
      port map(A => \REGMAP_i_i[33]\, B => \REGMAP[34]_net_1\, Y
         => N_441_0);
    
    \REG_1[391]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_356\, CLR => 
        \un10_hwres_19\, Q => \REG[391]\);
    
    \REG_1[132]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_140\, CLR => 
        \un10_hwres_8\, Q => \REG[132]\);
    
    REG_1_276 : MUX2H
      port map(A => VDB_in(14), B => \REG[263]\, S => 
        N_2816_i_0_0, Y => \REG_1_276\);
    
    PIPEA_610 : MUX2H
      port map(A => \PIPEA_7[21]\, B => \PIPEA[21]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_610\);
    
    \REG_88[87]\ : NOR2FT
      port map(A => N_2158, B => N_2566, Y => \REG_88[87]_net_1\);
    
    PULSE_1_244 : MUX2H
      port map(A => N_2387, B => \PULSE[9]\, S => un1_STATE1_17, 
        Y => \PULSE_1_244\);
    
    \PULSE_42_f0_i_o2[7]\ : NOR2FT
      port map(A => \REGMAP_i_0_i[11]\, B => PULSE_0_sqmuxa_1_2, 
        Y => N_2416_i);
    
    OR_RDATA_189 : MUX2H
      port map(A => N_29, B => \OR_RDATA[7]_net_1\, S => N_1832, 
        Y => \OR_RDATA_189\);
    
    \VAS[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_61\, CLR => HWRES_c_22, 
        Q => \VAS[10]_net_1\);
    
    un87_reg_ads_0_a3_0_a2_0 : NOR2FT
      port map(A => \VAS[2]_net_1\, B => N_198, Y => N_675);
    
    \REGMAP_0[29]\ : DFF
      port map(CLK => CLK_c_c, D => \un105_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[29]_net_1\);
    
    \REG_1[134]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_142\, CLR => 
        \un10_hwres_8_0\, Q => \REG[134]\);
    
    \LB_i_6_r[20]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_1, C => N_2202, 
        Y => \LB_i_6[20]\);
    
    \REG_i[285]\ : INV
      port map(A => \REG[285]\, Y => REG_i_0_280);
    
    \VDBi_18[1]\ : MUX2H
      port map(A => \VDBi_16[1]\, B => \REG[49]\, S => \TST_c[5]\, 
        Y => \VDBi_18[1]_net_1\);
    
    \REG_1[500]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_441\, SET => 
        \un10_hwres_27\, Q => \REG[500]\);
    
    \WDOG[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \WDOG_3[3]\, CLR => 
        un15_hwres_i, Q => \WDOG[3]_net_1\);
    
    \REG_1[136]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_144\, CLR => 
        \un10_hwres_8_0\, Q => \REG[136]\);
    
    un1_LB_DOUT_0_sqmuxa_0_1 : OR3FTT
      port map(A => N_2429, B => \STATE1[0]_net_1\, C => N_2408, 
        Y => un1_LB_DOUT_0_sqmuxa_0_1_i);
    
    CYCSF1 : DFFC
      port map(CLK => CLK_c_c, D => \CYCSF1_17\, CLR => 
        HWRES_c_13, Q => \CYCSF1\);
    
    \VDBi_16_1_a2_2[1]\ : NOR2FT
      port map(A => \REGMAP[6]_net_1\, B => \REGMAP_0[2]_net_1\, 
        Y => N_2511);
    
    \REG_1[251]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_264\, CLR => 
        \un10_hwres_14\, Q => \REG[251]\);
    
    \VADm[16]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[16]_net_1\, Y => VADm(16));
    
    \VDBi_66_0[0]\ : MUX2H
      port map(A => \REG[393]\, B => \REG[377]\, S => 
        \REGMAP[29]_net_1\, Y => N_2017);
    
    \LB_i[5]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_517\, CLR => 
        HWRES_c_16, Q => \LB_i[5]_net_1\);
    
    \VDBi_66[0]\ : MUX2H
      port map(A => \VDBi_60[0]_net_1\, B => N_2017, S => N_2033, 
        Y => \VDBi_66[0]_net_1\);
    
    STATE1_tr12_7_0_o2_0 : OR2
      port map(A => \TCNT_i_i[6]\, B => \TCNT[7]_net_1\, Y => 
        STATE1_tr12_7_0_o2_0_i);
    
    un1_STATE1_34_0_1 : AO21TTF
      port map(A => N_2535, B => \STATE1_0[9]_net_1\, C => 
        \un1_STATE1_34_0_0\, Y => un1_STATE1_34_1);
    
    \LB_ADDR[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_545\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[2]_net_1\);
    
    REG_1_239 : MUX2H
      port map(A => VDB_in(14), B => \REG[199]\, S => N_2752_i_0, 
        Y => \REG_1_239\);
    
    \VDBm_0[20]\ : MUX2H
      port map(A => \PIPEB[20]_net_1\, B => \PIPEA[20]_net_1\, S
         => \BLTCYC_1\, Y => N_2316);
    
    VDBi_632 : MUX2H
      port map(A => \VDBi_92[11]\, B => \VDBi[11]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_632\);
    
    LB_ADDR_0_sqmuxa_2_0 : AO21TTF
      port map(A => \LB_ADDR_0_sqmuxa_1\, B => \REGMAP[36]_net_1\, 
        C => LB_DOUT_0_sqmuxa_0, Y => LB_ADDR_0_sqmuxa_2);
    
    \REG_1[169]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_209\, CLR => 
        \un10_hwres_10\, Q => \REG[169]\);
    
    LB_DOUT_157 : MUX2H
      port map(A => VDB_in(9), B => \LB_DOUT[9]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_157\);
    
    \VDBi_66[9]\ : MUX2H
      port map(A => \VDBi_60[9]_net_1\, B => N_2026, S => N_2033, 
        Y => \VDBi_66[9]_net_1\);
    
    \VDBi_16_1_a2[15]\ : AND2
      port map(A => N_2511_0, B => REG_46, Y => N_2496_i);
    
    \PIPEA_m[23]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA[23]_net_1\, Y => 
        \PIPEA_m[23]_net_1\);
    
    \LB_i_6_1[12]\ : MUX2H
      port map(A => VDB_in_0(12), B => \LB_DOUT[12]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2194);
    
    \LB_i[12]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_524\, CLR => 
        HWRES_c_14, Q => \LB_i[12]_net_1\);
    
    \VADm[1]\ : NOR2FT
      port map(A => \PIPEA[1]_net_1\, B => N_2507_0, Y => VADm(1));
    
    \VDBi_16_r[15]\ : OA21TTF
      port map(A => N_2497_i, B => N_2496_i, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[15]\);
    
    STATE1_tr12_7_0_o2_2 : OR2
      port map(A => \TCNT_i_i[2]\, B => \TCNT[3]_net_1\, Y => 
        STATE1_tr12_7_0_o2_2_i);
    
    un1_STATE1_34_0_a2_0 : OR2FT
      port map(A => \STATE1_0[7]_net_1\, B => \TST_c_0[2]\, Y => 
        N_2542);
    
    \PIPEA1_9_i[31]\ : AND2
      port map(A => DPR(31), B => N_85_0, Y => N_296);
    
    PIPEA1_576 : MUX2H
      port map(A => N_280, B => \PIPEA1[20]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_576\);
    
    \PIPEA1[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_564\, CLR => CLEAR_23, 
        Q => \PIPEA1[8]_net_1\);
    
    \VDBi_92_iv_0_2[7]\ : AOI21TTF
      port map(A => \LB_s[7]_net_1\, B => N_7_i, C => 
        \VDBi_92_iv_0_1[7]_net_1\, Y => \VDBi_92_iv_0_2[7]_net_1\);
    
    un1_STATE1_20_i_a2_0_a2 : AND3FTT
      port map(A => N_83_0, B => \un1_STATE1_20_i_a2_0_a2_2\, C
         => N_446, Y => N_2454);
    
    \VDBi_23[17]\ : MUX2H
      port map(A => \VDBi_18[17]_net_1\, B => \REG_i[499]_net_1\, 
        S => \REGMAP_1[13]_net_1\, Y => \VDBi_23[17]_net_1\);
    
    \LB_i[10]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_522\, CLR => 
        HWRES_c_14, Q => \LB_i[10]_net_1\);
    
    un1_LBUSTMO_1_I_9 : XOR2FT
      port map(A => N_66_0, B => \LBUSTMO_i_0_i[1]\, Y => 
        \DWACT_ADD_CI_0_pog_array_0[0]\);
    
    \REGMAP[11]\ : DFF
      port map(CLK => CLK_c_c, D => \un46_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_0_i[11]\);
    
    PIPEA_619 : MUX2H
      port map(A => \PIPEA_7[30]\, B => \PIPEA[30]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_619\);
    
    \PIPEB_4_i[10]\ : AND2
      port map(A => DPR(10), B => N_616_1, Y => N_2624);
    
    \PIPEA1_9_i[18]\ : AND2
      port map(A => DPR(18), B => N_85_4, Y => N_276);
    
    \REG_1_m[255]\ : NAND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[255]\, Y => 
        \REG_1_m[255]_net_1\);
    
    \VDBi_55[22]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[22]_net_1\, Y => \VDBi_55[22]_net_1\);
    
    un1_STATE1_20_i_a2_0_a2_2 : AND2FT
      port map(A => N_1698, B => \un1_STATE1_17_0_1\, Y => 
        \un1_STATE1_20_i_a2_0_a2_2\);
    
    \LB_i_6_r[31]\ : AND3
      port map(A => N_2572_0, B => LB_i_6_sn_N_2_0, C => N_2213, 
        Y => \LB_i_6[31]\);
    
    \REGMAP_0[19]\ : DFF
      port map(CLK => CLK_c_c, D => \un64_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[19]_net_1\);
    
    LB_s_86 : MUX2H
      port map(A => LB_in(7), B => \LB_s[7]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_86\);
    
    \REG_1[266]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_279\, CLR => 
        \un10_hwres_15\, Q => \REG[266]\);
    
    un105_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_683_i, B => un105_reg_ads_1_0, Y => 
        \un105_reg_ads_0_a3_0_a2\);
    
    STATE1_tr27_i_o2 : OR2FT
      port map(A => \SINGCYC_0\, B => N_2565, Y => N_2532);
    
    SINGCYC_0 : DFFC
      port map(CLK => CLK_c_c, D => \SINGCYC_147\, CLR => 
        HWRES_c_21_0, Q => \SINGCYC_0\);
    
    \VDBi_53_0_iv_2[0]\ : AO21TTF
      port map(A => \REGMAP[20]_net_1\, B => \REG[185]\, C => 
        \REG_1_m[169]_net_1\, Y => \VDBi_53_0_iv_2_i[0]\);
    
    \VDBi_53_0_iv_5[3]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[3]\, B => 
        \VDBi_53_0_iv_0_i[3]\, C => \VDBi_53_0_iv_1_i[3]\, Y => 
        \VDBi_53_0_iv_5_i[3]\);
    
    REG3_125 : MUX2H
      port map(A => \REG[12]\, B => VDB_in(12), S => 
        REG1_0_sqmuxa_0, Y => \REG3_125\);
    
    \VDBi_23[16]\ : MUX2H
      port map(A => \VDBi_18[16]_net_1\, B => \REG_i[498]_net_1\, 
        S => \REGMAP_1[13]_net_1\, Y => \VDBi_23[16]_net_1\);
    
    un25_reg_ads_0_a3_0_a2_0 : OR2
      port map(A => N_678, B => \WRITES\, Y => N_694);
    
    EVREADi : DFFC
      port map(CLK => CLK_c_c, D => \EVREADi_181\, CLR => 
        CLEAR_20, Q => \EVREAD\);
    
    \STATE1_0[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[2]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1_0[8]_net_1\);
    
    \PIPEB[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_31\, CLR => CLEAR_26, 
        Q => \PIPEB[11]_net_1\);
    
    un90_reg_ads_0_a3_0_a2_0 : OR2
      port map(A => N_671, B => \WRITES_1\, Y => 
        un90_reg_ads_0_a3_0_a2_0_i);
    
    \LB_i_6_r[9]\ : AND2
      port map(A => N_2225, B => N_2572_2, Y => \LB_i_6[9]_net_1\);
    
    \REG_1[248]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_261\, SET => 
        \un10_hwres_14\, Q => \REG[248]\);
    
    \STATE1_ns_0_iv_0_0_a2_1[1]\ : OR3FTT
      port map(A => \REGMAP[36]_net_1\, B => \LB_ACK_sync\, C => 
        N_2455_1, Y => N_629);
    
    un1_STATE1_6_i_a2_0_o2_0 : OR2FT
      port map(A => N_2524, B => \STATE1_0[1]_net_1\, Y => N_83_0);
    
    un1_LBUSTMO_1_I_16 : XOR2FT
      port map(A => N_66, B => \LBUSTMO_i_0_i[1]\, Y => 
        \DWACT_ADD_CI_0_partial_sum[1]\);
    
    \REG_1[283]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_296\, CLR => 
        \un10_hwres_16\, Q => \REG[283]\);
    
    \LB_s[31]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_110\, CLR => 
        HWRES_c_19, Q => \LB_s[31]_net_1\);
    
    REG_1_454 : MUX2H
      port map(A => VDB_in(31), B => \REG[513]\, S => N_3170_i_0, 
        Y => \REG_1_454\);
    
    \REG_1[503]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_444\, CLR => 
        \un10_hwres_27\, Q => \REG[503]\);
    
    REG_1_410 : MUX2H
      port map(A => VDB_in_0(4), B => \REG[445]\, S => N_3104_i, 
        Y => \REG_1_410\);
    
    \VAS[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_58\, CLR => HWRES_c_23, 
        Q => \VAS[7]_net_1\);
    
    REG_1_474 : MUX2H
      port map(A => VDB_in(19), B => \REG[67]\, S => N_3234_i_1, 
        Y => \REG_1_474\);
    
    \VDBi_53_0_iv_3[3]\ : AO21TTF
      port map(A => \REGMAP[16]_net_1\, B => \REG_0[124]\, C => 
        \VDBi_53_0_iv_2[3]_net_1\, Y => \VDBi_53_0_iv_3_i[3]\);
    
    un1_STATE1_32_0_3 : AOI21TTF
      port map(A => N_83_0, B => N_2531, C => \un1_STATE1_32_0_2\, 
        Y => \un1_STATE1_32_0_3\);
    
    \VDBi_18[27]\ : NAND2
      port map(A => \REG[75]\, B => \TST_c_0[5]\, Y => 
        \VDBi_18[27]_net_1\);
    
    \REGMAP_0[20]\ : DFF
      port map(CLK => CLK_c_c, D => \un67_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[20]_net_1\);
    
    VDBi_650 : MUX2H
      port map(A => \VDBi_92[29]\, B => \VDBi[29]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_650\);
    
    \REG_1[287]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_300\, CLR => 
        \un10_hwres_16\, Q => \REG[287]\);
    
    un2_vsel_1_i_a2_1 : NAND3FFT
      port map(A => un2_vsel_1_i_a2_1_0_i, B => 
        un2_vsel_1_i_a2_1_1_i, C => N_2403, Y => N_237);
    
    \PIPEA[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_610\, CLR => CLEAR_24, 
        Q => \PIPEA[21]_net_1\);
    
    \LB_DOUT[28]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_176\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[28]_net_1\);
    
    \VDBm[18]\ : MUX2H
      port map(A => N_2314, B => \VDBi[18]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_18);
    
    VAS_62 : MUX2H
      port map(A => \VAS[11]_net_1\, B => VAD_in_10, S => 
        \TST_c_0[1]\, Y => \VAS_62\);
    
    \LB_i_6[3]\ : MUX2H
      port map(A => N_2173, B => N_2185, S => LB_i_6_sn_N_2, Y
         => N_2219);
    
    un1_TCNT_1_I_45 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_5[0]\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_6[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    \STATE1_ns_0_iv_0_0_a2[4]\ : NOR2FT
      port map(A => \STATE1[6]_net_1\, B => \TST_c_0[2]\, Y => 
        N_570_i);
    
    REG_1_139 : MUX2H
      port map(A => \REG[131]\, B => VDB_in(10), S => 
        REG_0_sqmuxa_0, Y => \REG_1_139\);
    
    \STATE5_ns_0_0_a2_1_1[1]\ : AND2
      port map(A => \OR_RREQ_sync\, B => \STATE5[1]_net_1\, Y => 
        N_2597_1);
    
    \PIPEA1_9_i[15]\ : AND2
      port map(A => DPR(15), B => N_85_4, Y => N_270);
    
    \VDBi_77_0[10]\ : MUX2H
      port map(A => REG_466, B => \REG[451]\, S => 
        \REGMAP_i_i[33]\, Y => N_2062);
    
    \PIPEA_7_r[16]\ : AND2
      port map(A => N_85_1, B => N_525, Y => \PIPEA_7[16]\);
    
    \LB_s[8]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_87\, CLR => HWRES_c_19, 
        Q => \LB_s[8]_net_1\);
    
    \FBOUT_m[3]\ : NAND2
      port map(A => FBOUT(3), B => \STATE1[2]_net_1\, Y => 
        \FBOUT_m[3]_net_1\);
    
    \PIPEA_7_i_m2[23]\ : MUX2H
      port map(A => DPR(23), B => \PIPEA1[23]_net_1\, S => 
        N_1996_0, Y => N_532);
    
    un776_regmap_23_2 : OR3FFT
      port map(A => \un776_regmap_14\, B => \un776_regmap_19\, C
         => \TST_c_0[5]\, Y => un776_regmap_23_2_i);
    
    \VDBm[30]\ : MUX2H
      port map(A => N_2326, B => \VDBi[30]_net_1\, S => 
        \SINGCYC_0\, Y => VDBm_30);
    
    \VDBi[30]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_651\, CLR => 
        \un10_hwres_35\, Q => \VDBi[30]_net_1\);
    
    \VDBi_23[1]\ : MUX2H
      port map(A => \VDBi_18[1]_net_1\, B => \REG[483]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23[1]_net_1\);
    
    \LB_i_6_r[2]\ : AND2
      port map(A => N_2218, B => N_2572_3, Y => \LB_i_6[2]_net_1\);
    
    \VDBi_80[5]\ : MUX2H
      port map(A => \VDBi_77[5]_net_1\, B => REG_477, S => 
        \REGMAP[35]_net_1\, Y => \VDBi_80[5]_net_1\);
    
    N_28_i_i_0 : NAND2
      port map(A => N_425, B => N_479, Y => \N_2613_0\);
    
    \LB_i_6_r[7]\ : AND2
      port map(A => N_2223, B => N_2572_3, Y => \LB_i_6[7]_net_1\);
    
    un10_hwres_22 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_22\);
    
    \VDBm[28]\ : MUX2H
      port map(A => N_2324, B => \VDBi[28]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_28);
    
    \REG_1[99]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_506\, CLR => 
        \un10_hwres_32\, Q => \REG[99]\);
    
    \PULSE_42_f0_i[8]\ : OA21TTF
      port map(A => \PULSE[8]\, B => REG_0_sqmuxa_0, C => 
        \STATE1_0[7]_net_1\, Y => N_2386);
    
    \LB_i_6_1[3]\ : MUX2H
      port map(A => VDB_in_0(3), B => \LB_DOUT[3]_net_1\, S => 
        \STATE5[0]_net_1\, Y => N_2185);
    
    \VDBi_18[26]\ : NAND2
      port map(A => \REG[74]\, B => \TST_c_0[5]\, Y => 
        \VDBi_18[26]_net_1\);
    
    \RAMAD_VME[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_6\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[2]_net_1\);
    
    \REG_1[428]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_393\, CLR => 
        \un10_hwres_23\, Q => \REG[428]\);
    
    REG3_121 : MUX2H
      port map(A => \REG[8]\, B => VDB_in(8), S => 
        REG1_0_sqmuxa_0, Y => \REG3_121\);
    
    \VDBi_92_iv_0_1[7]\ : AOI21TTF
      port map(A => N_457_i_0, B => \PIPEA[7]_net_1\, C => 
        \VDBi_92_iv_0_0[7]_net_1\, Y => \VDBi_92_iv_0_1[7]_net_1\);
    
    un776_regmap_4 : NOR2
      port map(A => \REGMAP[15]_net_1\, B => \REGMAP[14]_net_1\, 
        Y => \un776_regmap_4\);
    
    REG_1_405_e_0 : OR2FT
      port map(A => \REGMAP_0[31]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_3072_i_0);
    
    REG_1_393 : MUX2H
      port map(A => VDB_in(19), B => \REG[428]\, S => N_3072_i_1, 
        Y => \REG_1_393\);
    
    \PIPEA[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_601\, CLR => CLEAR_23, 
        Q => \PIPEA[12]_net_1\);
    
    \VDBi_66_d[12]\ : MUX2H
      port map(A => SPULSE1_c_c, B => N_2029, S => N_2033_0, Y
         => \VDBi_66_d[12]_net_1\);
    
    VAS_58 : MUX2H
      port map(A => \VAS[7]_net_1\, B => VAD_in_6, S => 
        \TST_c_0[1]\, Y => \VAS_58\);
    
    REG_1_224_e : OR2FT
      port map(A => \REGMAP_0[19]_net_1\, B => PULSE_0_sqmuxa_1_2, 
        Y => N_2720_i);
    
    \STATE5_0[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns[0]\, CLR => 
        HWRES_c_21_0, Q => \STATE5_0[0]_net_1\);
    
    \VDBi_53_0_iv_2[2]\ : AOI21TTF
      port map(A => \REGMAP[19]_net_1\, B => \REG[171]\, C => 
        \REG_1_m[155]_net_1\, Y => \VDBi_53_0_iv_2[2]_net_1\);
    
    PIPEA1_580 : MUX2H
      port map(A => N_288, B => \PIPEA1[24]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_580\);
    
    \OR_RDATA[9]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_191\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[9]_net_1\);
    
    \LB_i_6_r[1]\ : AND2
      port map(A => N_2217, B => N_2572_3, Y => \LB_i_6[1]_net_1\);
    
    \LB_i_6_1[5]\ : MUX2H
      port map(A => VDB_in_0(5), B => \LB_DOUT[5]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2187);
    
    \PIPEB[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_39\, CLR => CLEAR_26, 
        Q => \PIPEB[19]_net_1\);
    
    \VDBi_23[14]\ : MUX2H
      port map(A => \VDBi_16[14]\, B => \VDBi_23_d[14]_net_1\, S
         => \VDBi_23_s[7]_net_1\, Y => \VDBi_23[14]_net_1\);
    
    \OR_RACK\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RACK_1_sqmuxa_i_i_a2\, 
        CLR => HWRES_c_19, Q => OR_RACK);
    
    \VDBi_55[6]\ : OA21TTF
      port map(A => \VDBi_23_m_i[6]\, B => \VDBi_53_0_iv_5_i[6]\, 
        C => \REGMAP[26]_net_1\, Y => \VDBi_55[6]_net_1\);
    
    un98_reg_ads_0_a3_0_a2 : NOR3FFT
      port map(A => \WRITES_1\, B => N_682, C => un98_reg_ads_1, 
        Y => \un98_reg_ads_0_a3_0_a2\);
    
    REG_1_236 : MUX2H
      port map(A => VDB_in(11), B => \REG[196]\, S => N_2752_i_0, 
        Y => \REG_1_236\);
    
    PIPEB_34 : MUX2H
      port map(A => \PIPEB[14]_net_1\, B => N_2628, S => N_1996_4, 
        Y => \PIPEB_34\);
    
    \VDBi_92_iv[6]\ : OAI21FTT
      port map(A => \VDBi_80[6]_net_1\, B => \N_2613_0\, C => 
        \VDBi_92_iv_2[6]_net_1\, Y => \VDBi_92[6]\);
    
    un776_regmap_20 : OR3
      port map(A => \REGMAP_0[29]_net_1\, B => 
        \REGMAP_0[7]_net_1\, C => \REGMAP_0[13]_net_1\, Y => 
        un776_regmap_20_i);
    
    un1_STATE1_28_i_a2_1_0 : AND2
      port map(A => \WRITES\, B => \REGMAP[36]_net_1\, Y => 
        \un1_STATE1_28_i_a2_1_0\);
    
    REG_1_460 : MUX2H
      port map(A => VDB_in_0(5), B => \REG[53]\, S => N_3234_i, Y
         => \REG_1_460\);
    
    \OR_RDATA_5_i[2]\ : AND2
      port map(A => N_2572, B => LB_in(2), Y => N_19);
    
    ADACKCYC_76 : MUX2H
      port map(A => \ADACKCYC\, B => \TST_c_0[1]\, S => N_59, Y
         => \ADACKCYC_76\);
    
    REG_1_224_e_0 : OR2FT
      port map(A => \REGMAP_0[19]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_2720_i_0);
    
    un1_LB_DOUT_0_sqmuxa_0_o2 : OR2FT
      port map(A => N_462, B => \STATE1_0[7]_net_1\, Y => N_2408);
    
    REG_1_365 : MUX2H
      port map(A => VDB_in_0(7), B => \REG[400]\, S => N_3008_i, 
        Y => \REG_1_365\);
    
    \REG_1[393]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_358\, CLR => 
        \un10_hwres_20\, Q => \REG[393]\);
    
    \REG_1[161]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_201\, CLR => 
        \un10_hwres_9\, Q => \REG[161]\);
    
    un1_STATE2_12_0_0_0 : OAI21FTF
      port map(A => \STATE2[2]_net_1\, B => N_472_i_0, C => 
        un1_STATE2_12_0_0_1_i, Y => un1_STATE2_13_4_0);
    
    \LB_i_6[10]\ : MUX2H
      port map(A => N_2180, B => N_2192, S => LB_i_6_sn_N_2_1, Y
         => N_2226);
    
    \VDBi_60[29]\ : MUX2H
      port map(A => \VDBi_55[29]_net_1\, B => LBSP_in_29, S => 
        \REGMAP_0[28]_net_1\, Y => \VDBi_60[29]_net_1\);
    
    REG_1_240_e_0 : OR2FT
      port map(A => \REGMAP_0[20]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_2752_i_0);
    
    \REG_1[83]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_490\, CLR => 
        \un10_hwres_31\, Q => \REG[83]\);
    
    \VDBi[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_631\, CLR => 
        \un10_hwres_33\, Q => \VDBi[10]_net_1\);
    
    \PIPEB_4_i[7]\ : AND2
      port map(A => DPR(7), B => N_616, Y => N_2621);
    
    \PIPEA_7_r[19]\ : AND2
      port map(A => N_85_1, B => N_528, Y => \PIPEA_7[19]\);
    
    \VDBi_55[26]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[26]_net_1\, Y => \VDBi_55[26]_net_1\);
    
    un123_reg_ads_0_a2_3_a2 : NOR2
      port map(A => N_672, B => un84_reg_ads_1, Y => 
        \un123_reg_ads_0_a2_3_a2\);
    
    \PIPEA[29]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEA_618\, SET => CLEAR_25, 
        Q => \PIPEA[29]_net_1\);
    
    \REG_i[296]\ : INV
      port map(A => \REG[296]\, Y => REG_i_0_291);
    
    \LBUSTMO_3_0[1]\ : OR2FT
      port map(A => N_2572_0, B => I_19_0, Y => \LBUSTMO_3[1]\);
    
    \VDBi_60[13]\ : MUX2H
      port map(A => \VDBi_58[13]_net_1\, B => SPULSE2_c_c, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[13]_net_1\);
    
    PIPEB_27 : MUX2H
      port map(A => \PIPEB[7]_net_1\, B => N_2621, S => N_1996, Y
         => \PIPEB_27\);
    
    \REG_1_m[262]\ : NAND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[262]\, Y => 
        \REG_1_m[262]_net_1\);
    
    un10_hwres_9 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_9\);
    
    \PIPEB[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_26\, CLR => CLEAR_28, 
        Q => \PIPEB[6]_net_1\);
    
    \LB_i[2]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_514\, CLR => 
        HWRES_c_16, Q => \LB_i[2]_net_1\);
    
    REG_1_203 : MUX2H
      port map(A => VDB_in(10), B => \REG[163]\, S => N_2688_i_0, 
        Y => \REG_1_203\);
    
    \VDBi_92_0_iv_1[19]\ : AOI21TTF
      port map(A => \LB_s[19]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[19]_net_1\, Y => 
        \VDBi_92_0_iv_1[19]_net_1\);
    
    un1_STATE2_16_0_o2_0_o2 : AND2FT
      port map(A => \STATE2[0]_net_1\, B => N_584, Y => N_79);
    
    RAMAD_VME_9 : MUX2H
      port map(A => \VAS[6]_net_1\, B => \RAMAD_VME[5]_net_1\, S
         => N_2523_0, Y => \RAMAD_VME_9\);
    
    \REG_1_m[157]\ : NAND2
      port map(A => \REGMAP[18]_net_1\, B => \REG[157]\, Y => 
        \REG_1_m[157]_net_1\);
    
    \VDBi_80_s[3]\ : NOR2FT
      port map(A => \VDBi_77_s[3]_net_1\, B => \REGMAP[35]_net_1\, 
        Y => \VDBi_80_s[3]_net_1\);
    
    \PIPEA1_9_i[20]\ : AND2
      port map(A => DPR(20), B => N_85_3, Y => N_280);
    
    un776_regmap_0 : OR2
      port map(A => \REGMAP_i_0_i[11]\, B => \REGMAP[25]_net_1\, 
        Y => un776_regmap_0_i);
    
    un1_TCNT_1_I_22 : XOR2
      port map(A => \TCNT[7]_net_1\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum[7]\);
    
    \VDBi_16_1_a3_2_1[0]\ : NOR2
      port map(A => \REGMAP[2]_net_1\, B => \REGMAP[6]_net_1\, Y
         => N_2380_1);
    
    \PIPEB[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_42\, CLR => CLEAR_27, 
        Q => \PIPEB[22]_net_1\);
    
    un21_reg_ads_0_a3_0_a2 : NOR3FTT
      port map(A => N_682, B => \WRITES_1\, C => N_681_i, Y => 
        \un21_reg_ads_0_a3_0_a2\);
    
    \VDBi_16_r[6]\ : OA21TTF
      port map(A => \VDBi_16_1_0_i[6]\, B => N_2476_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[6]\);
    
    \REG_1[382]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_347\, CLR => 
        \un10_hwres_19\, Q => \REG[382]\);
    
    BLTCYC_0 : DFFC
      port map(CLK => CLK_c_c, D => \BLTCYC_77\, CLR => 
        HWRES_c_13_0, Q => \BLTCYC_0\);
    
    un102_reg_ads_0_a3_0_a2_0 : AND2
      port map(A => N_673, B => \VAS[6]_net_1\, Y => N_688);
    
    un1_LBUSTMO_1_I_21 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, Y => I_21_1);
    
    NDTKIN : OR2
      port map(A => \CLOSEDTK\, B => \TST_c_c[3]\, Y => NDTKIN_c);
    
    \REG_1[84]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_491\, CLR => 
        \un10_hwres_31\, Q => \REG[84]\);
    
    REG_1_207 : MUX2H
      port map(A => VDB_in(14), B => \REG[167]\, S => N_2688_i_0, 
        Y => \REG_1_207\);
    
    PIPEB_38 : MUX2H
      port map(A => \PIPEB[18]_net_1\, B => N_199, S => N_1996_4, 
        Y => \PIPEB_38\);
    
    \VDBi_16_1_a2[10]\ : AND2
      port map(A => N_2511_0, B => REG_41, Y => N_2486_i);
    
    \REG_1[73]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_480\, CLR => 
        \un10_hwres_30\, Q => \REG[73]\);
    
    \VDBi_23_d[4]\ : MUX2H
      port map(A => \REG[52]\, B => \REG[486]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23_d[4]_net_1\);
    
    \REG_1[488]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_429\, SET => 
        \un10_hwres_26\, Q => \REG[488]\);
    
    un10_hwres_27 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_27\);
    
    \VAS[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_59\, CLR => HWRES_c_23, 
        Q => \VAS[8]_net_1\);
    
    \PIPEA_m[20]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[20]_net_1\, Y => 
        \PIPEA_m[20]_net_1\);
    
    VDBi_648 : MUX2H
      port map(A => \VDBi_92[27]\, B => \VDBi[27]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_648\);
    
    \LB_DOUT[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_160\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[12]_net_1\);
    
    \REGMAP[35]\ : DFF
      port map(CLK => CLK_c_c, D => \un123_reg_ads_0_a2_3_a2\, Q
         => \REGMAP[35]_net_1\);
    
    un10_hwres_2 : OR2
      port map(A => HWRES_c_0_6, B => \WDOGTO\, Y => 
        \un10_hwres_2\);
    
    un1_STATE2_13_i_0_a2_1_0_0 : OR2
      port map(A => DPR(29), B => DPR(31), Y => 
        \un1_STATE2_13_i_0_a2_1_0_0\);
    
    \PIPEB[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_22\, CLR => CLEAR_27, 
        Q => \PIPEB[2]_net_1\);
    
    STATE5_0_sqmuxa_0_a3_0_a2 : NAND2FT
      port map(A => N_2608, B => N_2606_i_i, Y => STATE5_0_sqmuxa);
    
    \REG_1[386]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_351\, CLR => 
        \un10_hwres_19\, Q => \REG[386]\);
    
    un10_hwres_23 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_23\);
    
    nLBLAST_112 : MUX2H
      port map(A => \STATE5_i_0[0]\, B => \NLBLAST_c\, S => 
        N_1828, Y => \nLBLAST_112\);
    
    \VDBi_77_0_i_m2[7]\ : MUX2H
      port map(A => REG_463, B => \REG[448]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_493);
    
    BLTCYC_2 : DFFC
      port map(CLK => CLK_c_c, D => \BLTCYC_77\, CLR => 
        HWRES_c_13_0, Q => \BLTCYC_2\);
    
    \PIPEA1_9_i[1]\ : AND2
      port map(A => DPR(1), B => N_85, Y => N_242);
    
    \LB_i[25]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_537\, CLR => 
        HWRES_c_15, Q => \LB_i[25]_net_1\);
    
    \REG_1[280]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_293\, CLR => 
        \un10_hwres_15\, Q => \REG[280]\);
    
    \VDBi_92_0_iv_1[11]\ : AOI21TTF
      port map(A => \LB_s[11]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[11]_net_1\, Y => 
        \VDBi_92_0_iv_1[11]_net_1\);
    
    \REG3[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_121\, CLR => 
        \un10_hwres_7\, Q => \REG[8]\);
    
    \LB_i_6_1[28]\ : MUX2H
      port map(A => VDB_in(28), B => \LB_DOUT[28]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2210);
    
    \REG_1[97]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_504\, CLR => 
        \un10_hwres_31\, Q => \REG[97]\);
    
    \REG_88_0[86]\ : MUX2H
      port map(A => VDB_in_0(5), B => \REG[86]\, S => N_20, Y => 
        N_2157);
    
    REG_1_397 : MUX2H
      port map(A => VDB_in(23), B => \REG[432]\, S => N_3072_i_0, 
        Y => \REG_1_397\);
    
    MYBERRi_19 : MUX2H
      port map(A => \MYBERR_c\, B => \TST_c[2]\, S => 
        un1_MYBERRi_1_sqmuxa, Y => \MYBERRi_19\);
    
    \REG_1[446]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_411\, CLR => 
        \un10_hwres_24\, Q => \REG[446]\);
    
    \VDBi_16_1_a3_0[0]\ : AND2
      port map(A => N_2511, B => REG_31, Y => N_2377_i);
    
    \VDBi_92_iv_1[2]\ : AOI21TTF
      port map(A => N_457_i_0, B => \PIPEA[2]_net_1\, C => 
        \VDBi_92_iv_0[2]_net_1\, Y => \VDBi_92_iv_1[2]_net_1\);
    
    \VDBi_66_0[5]\ : MUX2H
      port map(A => \REG[398]\, B => \REG[382]\, S => 
        \REGMAP[29]_net_1\, Y => N_2022);
    
    \PIPEA[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_607\, CLR => CLEAR_24, 
        Q => \PIPEA[18]_net_1\);
    
    REG_1_491 : MUX2H
      port map(A => \REG_88[84]_net_1\, B => \REG[84]\, S => 
        un1_STATE1_15, Y => \REG_1_491\);
    
    REG_1_485 : MUX2H
      port map(A => VDB_in(30), B => \REG[78]\, S => N_3234_i_0, 
        Y => \REG_1_485\);
    
    LB_i_533 : MUX2H
      port map(A => \LB_i[21]_net_1\, B => \LB_i_6[21]\, S => 
        N_2570_0, Y => \LB_i_533\);
    
    REG_1_434 : MUX2H
      port map(A => VDB_in_0(11), B => \REG[493]\, S => 
        N_3170_i_1, Y => \REG_1_434\);
    
    PULSE_1_241 : MUX2H
      port map(A => \PULSE_42[6]\, B => \PULSE[6]\, S => 
        un1_STATE1_17, Y => \PULSE_1_241\);
    
    \VDBm[1]\ : MUX2H
      port map(A => N_2297, B => \VDBi[1]_net_1\, S => \SINGCYC\, 
        Y => VDBm_1);
    
    \REG_1[74]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_481\, CLR => 
        \un10_hwres_30\, Q => \REG[74]\);
    
    \REG_1[239]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_252\, SET => 
        \un10_hwres_13\, Q => \REG[239]\);
    
    LB_s_87 : MUX2H
      port map(A => LB_in(8), B => \LB_s[8]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_87\);
    
    \PIPEA1_9_i[11]\ : AND2
      port map(A => DPR(11), B => N_85_4, Y => N_262);
    
    REG_1_131 : MUX2H
      port map(A => \REG[123]\, B => VDB_in(2), S => REG_0_sqmuxa, 
        Y => \REG_1_131\);
    
    \REG3_0_0[514]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_514_180\, CLR => 
        \un10_hwres_6_0\, Q => \RUN_c_0_0\);
    
    WRITES_1 : DFFC
      port map(CLK => CLK_c_c, D => \WRITES_2\, CLR => 
        HWRES_c_23_0, Q => \WRITES_1\);
    
    un2_vsel_1_i_a2_0 : OR2
      port map(A => AMB_c(1), B => N_228, Y => N_232);
    
    \PIPEA_m[27]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA[27]_net_1\, Y => 
        \PIPEA_m[27]_net_1\);
    
    un2_vsel_2_i_a2_1 : NAND2FT
      port map(A => N_237, B => AMB_c(0), Y => N_2434_1);
    
    PIPEB_42 : MUX2H
      port map(A => \PIPEB[22]_net_1\, B => N_2634, S => N_1996_3, 
        Y => \PIPEB_42\);
    
    \VDBi_16_1_a2_1[7]\ : NAND2
      port map(A => N_2512, B => \REG[7]\, Y => N_2480);
    
    SINGCYC_147 : OA21TTF
      port map(A => N_2436_i, B => \SINGCYC_0\, C => \TST_c_0[0]\, 
        Y => \SINGCYC_147\);
    
    nLBASi : DFFS
      port map(CLK => ALICLK_c, D => \nLBASi_3\, SET => 
        HWRES_c_23, Q => \nLBAS_c\);
    
    \LB_i_6_r[14]\ : AND3
      port map(A => N_2572_2, B => LB_i_6_sn_N_2_1, C => N_2196, 
        Y => \LB_i_6[14]\);
    
    \VDBi_77_0[4]\ : MUX2H
      port map(A => REG_460, B => \REG[445]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_2056);
    
    \REG_1[397]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_362\, CLR => 
        \un10_hwres_20\, Q => \REG[397]\);
    
    REG_1_486_e_0 : OR2FT
      port map(A => N_2409, B => un1_STATE1_15, Y => N_3234_i_0);
    
    \VDBi_92_0_iv_0_a2_0[25]\ : NAND2
      port map(A => N_723, B => \REG[434]\, Y => N_603);
    
    un1_TCNT_1_I_48 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_3[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_4[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    un10_hwres_28 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_0, Y => 
        \un10_hwres_28\);
    
    REQUESTER_1_i_0_a2 : NOR2FT
      port map(A => N_2572_0, B => \REQUESTER\, Y => N_2589);
    
    \REG_1[491]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_432\, CLR => 
        \un10_hwres_26\, Q => \REG[491]\);
    
    \PIPEA_7_r[5]\ : AND2
      port map(A => N_85_2, B => N_514, Y => \PIPEA_7[5]\);
    
    un776_regmap_13 : NOR3
      port map(A => \REGMAP[12]_net_1\, B => \REGMAP[27]_net_1\, 
        C => un776_regmap_6_i, Y => \un776_regmap_13\);
    
    REG_1_443 : MUX2H
      port map(A => VDB_in(20), B => \REG[502]\, S => N_3170_i_1, 
        Y => \REG_1_443\);
    
    PIPEB_30 : MUX2H
      port map(A => \PIPEB[10]_net_1\, B => N_2624, S => N_1996_4, 
        Y => \PIPEB_30\);
    
    \VDBi_92_0_iv[24]\ : OAI21FTT
      port map(A => \VDBi_71[24]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[24]_net_1\, Y => \VDBi_92[24]\);
    
    N_1897_o5_0_o2 : NAND2
      port map(A => \SINGCYC\, B => \STATE1[9]_net_1\, Y => 
        N_1898);
    
    \WDOG[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \WDOG_3[2]\, CLR => 
        un15_hwres_i, Q => \WDOG[2]_net_1\);
    
    REG_1_489 : MUX2H
      port map(A => \REG_88[82]_net_1\, B => \REG[82]\, S => 
        un1_STATE1_15, Y => \REG_1_489\);
    
    PIPEB_50 : MUX2H
      port map(A => \PIPEB[30]_net_1\, B => \PIPEB_4[30]\, S => 
        N_1996_3, Y => \PIPEB_50\);
    
    \VDBi_23_d[13]\ : MUX2H
      port map(A => \REG[61]\, B => \REG[495]\, S => 
        \REGMAP_1[13]_net_1\, Y => \VDBi_23_d[13]_net_1\);
    
    LB_DOUT_177 : MUX2H
      port map(A => VDB_in(29), B => \LB_DOUT[29]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_177\);
    
    PIPEB_21 : MUX2H
      port map(A => \PIPEB[1]_net_1\, B => N_2615, S => N_1996, Y
         => \PIPEB_21\);
    
    REG_1_214 : MUX2H
      port map(A => VDB_in(5), B => \REG[174]\, S => N_2720_i, Y
         => \REG_1_214\);
    
    REG_1_261_e_0 : OR2FT
      port map(A => \REGMAP_i_i_0[23]\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_2784_i_0);
    
    REG_1_212 : MUX2H
      port map(A => VDB_in(3), B => \REG[172]\, S => N_2720_i, Y
         => \REG_1_212\);
    
    \REG_1[414]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_379\, CLR => 
        \un10_hwres_21\, Q => \REG[414]\);
    
    \STATE1_ns_0_iv_0_0_a2[1]\ : OR2FT
      port map(A => \STATE1[9]_net_1\, B => N_436, Y => N_627);
    
    VDBi_643 : MUX2H
      port map(A => \VDBi_92[22]\, B => \VDBi[22]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_643\);
    
    un10_hwres_8_0 : OR2
      port map(A => HWRES_c_0_0, B => WDOGTO_0, Y => 
        \un10_hwres_8_0\);
    
    \STATE1_0[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[9]\, CLR => 
        \un10_hwres_32\, Q => \STATE1_0[1]_net_1\);
    
    \VDBi_53_0_iv_2[5]\ : AOI21TTF
      port map(A => \REGMAP[19]_net_1\, B => \REG[174]\, C => 
        \REG_1_m[158]_net_1\, Y => \VDBi_53_0_iv_2[5]_net_1\);
    
    REG_1_225 : MUX2H
      port map(A => VDB_in(0), B => \REG[185]\, S => N_2752_i, Y
         => \REG_1_225\);
    
    \REGMAP[25]\ : DFF
      port map(CLK => CLK_c_c, D => \un90_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[25]_net_1\);
    
    un779_regmap_i_0_a2 : NOR2
      port map(A => \REGMAP[36]_net_1\, B => \un776_regmap\, Y
         => N_2565);
    
    \REG_1[427]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_392\, CLR => 
        \un10_hwres_22\, Q => \REG[427]\);
    
    \PIPEA[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_596\, CLR => CLEAR_25, 
        Q => \PIPEA[7]_net_1\);
    
    \LB_i_6_1[21]\ : MUX2H
      port map(A => VDB_in(21), B => \LB_DOUT[21]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2203);
    
    \VDBi_80[6]\ : MUX2H
      port map(A => \VDBi_71[6]_net_1\, B => \VDBi_80_d[6]_net_1\, 
        S => \VDBi_80_s[2]_net_1\, Y => \VDBi_80[6]_net_1\);
    
    PIPEA_618 : MUX2H
      port map(A => \PIPEA_7[29]\, B => \PIPEA[29]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_618\);
    
    LB_i_6_sn_m1 : XOR2FT
      port map(A => \STATE5[1]_net_1\, B => \STATE5[0]_net_1\, Y
         => LB_i_6_sn_N_2);
    
    \LB_i[23]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_535\, CLR => 
        HWRES_c_15, Q => \LB_i[23]_net_1\);
    
    un1_TCNT_1_I_14 : XOR2
      port map(A => \TCNT[5]_net_1\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_4[0]\);
    
    un29_reg_ads_0_a2_0_a2_2_0 : OR2
      port map(A => \VAS[7]_net_1\, B => \VAS[8]_net_1\, Y => 
        \un29_reg_ads_0_a2_0_a2_2_0\);
    
    \LB_i_6_r[8]\ : AND2
      port map(A => N_2224, B => N_2572_3, Y => \LB_i_6[8]_net_1\);
    
    EVREADi_181 : MUX2H
      port map(A => \EVREAD\, B => \STATE2[2]_net_1\, S => N_16, 
        Y => \EVREADi_181\);
    
    \REG_1[62]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_469\, CLR => 
        \un10_hwres_29\, Q => \REG[62]\);
    
    \PIPEB[28]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEB_48\, SET => CLEAR_27, 
        Q => \PIPEB_i_i[28]\);
    
    \PIPEA_7_r[17]\ : AND2
      port map(A => N_85_1, B => N_526, Y => \PIPEA_7[17]\);
    
    REG_1_349 : MUX2H
      port map(A => VDB_in_0(7), B => \REG[384]\, S => N_2976_i, 
        Y => \REG_1_349\);
    
    un1_TCNT_1_I_1 : AND2
      port map(A => \TCNT_i_i[0]\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_TMP_1[0]\);
    
    PIPEB_35 : MUX2H
      port map(A => \PIPEB[15]_net_1\, B => N_2629, S => N_1996_4, 
        Y => \PIPEB_35\);
    
    \VDBi_60[26]\ : MUX2H
      port map(A => \VDBi_55[26]_net_1\, B => LBSP_in_26, S => 
        \REGMAP_0[28]_net_1\, Y => \VDBi_60[26]_net_1\);
    
    \VADm[9]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[9]_net_1\, Y => VADm(9));
    
    \PIPEA1[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_573\, CLR => CLEAR_21, 
        Q => \PIPEA1[17]_net_1\);
    
    REG_1_302 : MUX2H
      port map(A => VDB_in(24), B => \REG[289]\, S => N_2880_i_0, 
        Y => \REG_1_302\);
    
    \PIPEA_m[26]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA[26]_net_1\, Y => 
        \PIPEA_m[26]_net_1\);
    
    \OR_RDATA[4]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_186\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[4]_net_1\);
    
    un117_reg_ads_0_a3_0_a2_1 : NAND2
      port map(A => N_660, B => \VAS[6]_net_1\, Y => N_672);
    
    \VDBi_58[13]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[13]\, B => 
        \VDBi_23_m_i[13]\, C => \VDBi_58_0[9]\, Y => 
        \VDBi_58[13]_net_1\);
    
    \PIPEA1[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_574\, CLR => CLEAR_21, 
        Q => \PIPEA1[18]_net_1\);
    
    PIPEA1_585 : MUX2H
      port map(A => \PIPEA1_9[29]\, B => \PIPEA1[29]_net_1\, S
         => un1_STATE2_13_4_0, Y => \PIPEA1_585\);
    
    \VDBi_60[9]\ : MUX2H
      port map(A => \VDBi_58[9]_net_1\, B => \RUN_c_0_0\, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60[9]_net_1\);
    
    \STATE1_ns_1_iv_0[3]\ : OAI21FTT
      port map(A => N_2565, B => N_1898, C => 
        \STATE1_ns_1_iv_0_1[3]_net_1\, Y => \STATE1_ns[3]\);
    
    \RAMAD_VME[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_7\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[3]_net_1\);
    
    REG_1_408 : MUX2H
      port map(A => VDB_in_0(2), B => \REG[443]\, S => N_3104_i, 
        Y => \REG_1_408\);
    
    REG_1_221 : MUX2H
      port map(A => VDB_in(12), B => \REG[181]\, S => N_2720_i_0, 
        Y => \REG_1_221\);
    
    REG_1_193 : MUX2H
      port map(A => VDB_in(0), B => \REG[153]\, S => N_2688_i, Y
         => \REG_1_193\);
    
    \VDBi_58[10]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[10]\, B => 
        \VDBi_23_m_i[10]\, C => \VDBi_58_0[9]\, Y => 
        \VDBi_58[10]_net_1\);
    
    \VDBm[15]\ : MUX2H
      port map(A => N_2311, B => \VDBi[15]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_15);
    
    \VDBm_i_0_m2_0[21]\ : MUX2H
      port map(A => \PIPEB[21]_net_1\, B => \PIPEA[21]_net_1\, S
         => \BLTCYC_0\, Y => N_488);
    
    \LB_ADDR[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_549\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[6]_net_1\);
    
    \VDBi_92_iv[1]\ : OAI21FTT
      port map(A => \VDBi_80[1]_net_1\, B => \N_2613_0\, C => 
        \VDBi_92_iv_2[1]_net_1\, Y => \VDBi_92[1]\);
    
    \REG_1_m[121]\ : NAND2
      port map(A => \REGMAP[16]_net_1\, B => \REG[121]\, Y => 
        \REG_1_m[121]_net_1\);
    
    \VDBi_66_0[14]\ : MUX2H
      port map(A => \REG[407]\, B => \REG[391]\, S => 
        \REGMAP_0[29]_net_1\, Y => N_2031);
    
    \REG_1[55]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_462\, CLR => 
        \un10_hwres_28\, Q => \REG[55]\);
    
    un1_STATE5_10_i_1 : OAI21FTT
      port map(A => \LB_WRITE_sync\, B => N_66_0, C => N_2603, Y
         => N_2570_1);
    
    \REG_1[422]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_387\, SET => 
        \un10_hwres_22\, Q => \REG[422]\);
    
    REG_1_306 : MUX2H
      port map(A => VDB_in(28), B => \REG[293]\, S => N_2880_i_0, 
        Y => \REG_1_306\);
    
    un1_TCNT_1_I_21 : XOR2
      port map(A => \TCNT_i_i[2]\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[2]\);
    
    un105_reg_ads_0_a3_0_a2_0 : OR2
      port map(A => N_667, B => \VAS[1]_net_1\, Y => N_683_i);
    
    VDBi_634 : MUX2H
      port map(A => \VDBi_92[13]\, B => \VDBi[13]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_634\);
    
    N_28_i_i : NAND2
      port map(A => N_425, B => N_479, Y => N_2613);
    
    VDBi_639 : MUX2H
      port map(A => \VDBi_92[18]\, B => \VDBi[18]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_639\);
    
    \LB_i[1]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_513\, CLR => 
        HWRES_c_15, Q => \LB_i[1]_net_1\);
    
    REG_1_200 : MUX2H
      port map(A => VDB_in(7), B => \REG[160]\, S => N_2688_i, Y
         => \REG_1_200\);
    
    PIPEA1_563 : MUX2H
      port map(A => N_254, B => \PIPEA1[7]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_563\);
    
    \VDBm[25]\ : MUX2H
      port map(A => N_2321, B => \VDBi[25]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_25);
    
    \REG_1[193]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_233\, CLR => 
        \un10_hwres_12\, Q => \REG[193]\);
    
    \LB_s[25]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_104\, CLR => 
        HWRES_c_18, Q => \LB_s[25]_net_1\);
    
    un1_STATE1_32_0_a2_0 : OAI21
      port map(A => \PURGED\, B => \TST_c[2]\, C => N_480, Y => 
        N_2451);
    
    REG_1_507 : MUX2H
      port map(A => \REG[100]\, B => VDB_in_0(11), S => N_2416_i, 
        Y => \REG_1_507\);
    
    \VDBi_16_1_a3_1_0[0]\ : AND2
      port map(A => \RUN_c\, B => \REGMAP[14]_net_1\, Y => 
        \VDBi_16_1_a3_1_0[0]_net_1\);
    
    REG_1_264 : MUX2H
      port map(A => VDB_in(2), B => \REG[251]\, S => N_2816_i_0, 
        Y => \REG_1_264\);
    
    \REG_1[61]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_468\, CLR => 
        \un10_hwres_29\, Q => \REG[61]\);
    
    REG_1_262 : MUX2H
      port map(A => VDB_in(0), B => \REG[249]\, S => N_2816_i_0, 
        Y => \REG_1_262\);
    
    \LB_DOUT[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_171\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[23]_net_1\);
    
    \PIPEA_7_i_m2[9]\ : MUX2H
      port map(A => DPR(9), B => \PIPEA1[9]_net_1\, S => N_1996_2, 
        Y => N_518);
    
    \REG_1[384]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_349\, CLR => 
        \un10_hwres_19\, Q => \REG[384]\);
    
    \VAS[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_64\, CLR => HWRES_c_22, 
        Q => \VAS[13]_net_1\);
    
    N_2407_i_i_o2 : NOR2FT
      port map(A => \STATE1_0[9]_net_1\, B => \REGMAP[0]_net_1\, 
        Y => N_479);
    
    REG_1_248 : MUX2H
      port map(A => VDB_in(2), B => \REG[235]\, S => N_2784_i, Y
         => \REG_1_248\);
    
    \VDBi_16_1_a2_3[1]\ : NOR2FT
      port map(A => \VDBi_16_1_a2_3_0[1]_net_1\, B => 
        \REGMAP_0[2]_net_1\, Y => N_2512);
    
    RAMAD_VME_7 : MUX2H
      port map(A => \VAS[4]_net_1\, B => \RAMAD_VME[3]_net_1\, S
         => \TCNT_0_sqmuxa_i_s\, Y => \RAMAD_VME_7\);
    
    \PIPEA_7_r[15]\ : AND2
      port map(A => N_85_1, B => N_524, Y => \PIPEA_7[15]\);
    
    nLBRD : DFFS
      port map(CLK => ALICLK_c, D => \nLBRD_146\, SET => 
        HWRES_c_23_0, Q => \NLBRD_c\);
    
    LB_s_104 : MUX2H
      port map(A => LB_in(25), B => \LB_s[25]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_104\);
    
    \VDBi_71[14]\ : MUX2H
      port map(A => \VDBi_66[14]_net_1\, B => \REG[423]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[14]_net_1\);
    
    \REG_i[5]\ : INV
      port map(A => \REG[5]\, Y => REG_i_0_0);
    
    \REG_1[487]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_428\, CLR => 
        \un10_hwres_25\, Q => \REG[487]\);
    
    \VDBi_77[8]\ : MUX2H
      port map(A => \VDBi_66[8]_net_1\, B => \VDBi_77_d[8]_net_1\, 
        S => \VDBi_77_s[8]_net_1\, Y => \VDBi_77[8]_net_1\);
    
    REG_1_455 : MUX2H
      port map(A => VDB_in_0(0), B => \REG[48]\, S => N_3234_i, Y
         => \REG_1_455\);
    
    \REG_1[50]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_457\, CLR => 
        \un10_hwres_28\, Q => \REG[50]\);
    
    PIPEA1_581 : MUX2H
      port map(A => N_290, B => \PIPEA1[25]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_581\);
    
    VDBi_645 : MUX2H
      port map(A => \VDBi_92[24]\, B => \VDBi[24]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_645\);
    
    REG_1_475 : MUX2H
      port map(A => VDB_in(20), B => \REG[68]\, S => N_3234_i_1, 
        Y => \REG_1_475\);
    
    \VDBi_18[15]\ : MUX2H
      port map(A => \VDBi_16[15]\, B => \REG[63]\, S => 
        \TST_c_1[5]\, Y => \VDBi_18[15]_net_1\);
    
    \REG_1[236]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_249\, SET => 
        \un10_hwres_13\, Q => \REG[236]\);
    
    PIPEA_590 : MUX2H
      port map(A => \PIPEA_7[1]\, B => \PIPEA[1]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_590\);
    
    \REGMAP[9]\ : DFF
      port map(CLK => CLK_c_c, D => \un40_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[9]_net_1\);
    
    \REG_1_m[177]\ : NAND2
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[177]\, Y => 
        \REG_1_m[177]_net_1\);
    
    \REG_1[379]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_344\, CLR => 
        \un10_hwres_18\, Q => \REG[379]\);
    
    \REG_1[125]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_133\, CLR => 
        \un10_hwres_7_0\, Q => REG_124);
    
    \REG_1[167]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_207\, CLR => 
        \un10_hwres_10\, Q => \REG[167]\);
    
    PULSE_1_242 : MUX2H
      port map(A => N_2388, B => \PULSE[7]\, S => un1_STATE1_17, 
        Y => \PULSE_1_242\);
    
    LB_i_526 : MUX2H
      port map(A => \LB_i[14]_net_1\, B => \LB_i_6[14]\, S => 
        N_2570_1, Y => \LB_i_526\);
    
    \VDBi_80_d[6]\ : MUX2H
      port map(A => N_2058, B => REG_478, S => \REGMAP[35]_net_1\, 
        Y => \VDBi_80_d[6]_net_1\);
    
    \LB_s[4]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_83\, CLR => HWRES_c_19, 
        Q => \LB_s[4]_net_1\);
    
    VDBi_647 : MUX2H
      port map(A => \VDBi_92[26]\, B => \VDBi[26]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_647\);
    
    un1_STATE2_8_0_0_0_o2_0 : NAND2
      port map(A => N_426, B => \STATE2_i_0[3]\, Y => N_1996_0);
    
    un10_reg_ads_0_a2_1_a2 : NOR2FT
      port map(A => N_674, B => N_681_i, Y => 
        \un10_reg_ads_0_a2_1_a2\);
    
    \REG_1[404]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_369\, CLR => 
        \un10_hwres_21\, Q => \REG[404]\);
    
    LB_REQ_sync : DFFC
      port map(CLK => ALICLK_c, D => \LB_REQ\, CLR => HWRES_c_14, 
        Q => \LB_REQ_sync\);
    
    un1_TCNT_1_I_30 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum_0[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, Y => I_30_2);
    
    \VDBm_0[28]\ : MUX2H
      port map(A => \PIPEB_i_i[28]\, B => \PIPEA_i_0_i[28]\, S
         => \BLTCYC_1\, Y => N_2324);
    
    LB_s_110 : MUX2H
      port map(A => LB_in(31), B => \LB_s[31]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_110\);
    
    \VDBi_53_0_iv_2[11]\ : AOI21TTF
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[180]\, C => 
        \REG_1_m[164]_net_1\, Y => \VDBi_53_0_iv_2[11]_net_1\);
    
    \VDBi_53_0_iv_6[1]\ : NOR3
      port map(A => \VDBi_53_0_iv_5_i[1]\, B => 
        \VDBi_53_0_iv_2_i[1]\, C => \VDBi_53_0_iv_0_i[1]\, Y => 
        \VDBi_53_0_iv_6[1]_net_1\);
    
    REG_1_459 : MUX2H
      port map(A => VDB_in_0(4), B => \REG[52]\, S => N_3234_i, Y
         => \REG_1_459\);
    
    \PIPEA_7_r[21]\ : AND2
      port map(A => N_85_1, B => N_530, Y => \PIPEA_7[21]\);
    
    \REG_1[101]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_508\, CLR => 
        \un10_hwres_7\, Q => \REG[101]\);
    
    \PULSE_42_f0_i[7]\ : OA21TTF
      port map(A => \PULSE[7]\, B => N_2416_i, C => 
        \STATE1_0[7]_net_1\, Y => N_2388);
    
    \VDBi_77_0[1]\ : MUX2H
      port map(A => REG_457, B => \REG[442]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_2053);
    
    REG_1_479 : MUX2H
      port map(A => VDB_in(24), B => \REG[72]\, S => N_3234_i_0, 
        Y => \REG_1_479\);
    
    \REG_1[482]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_423\, SET => 
        \un10_hwres_25\, Q => \REG[482]\);
    
    LB_nOE_1_sqmuxa_0_o2 : NOR2
      port map(A => \LB_WRITE_sync\, B => N_1861, Y => N_2573);
    
    \LB_i_6_r[16]\ : AND3
      port map(A => N_2572_2, B => LB_i_6_sn_N_2_1, C => N_2198, 
        Y => \LB_i_6[16]\);
    
    VDBi_66_sn_m1_0 : OR2
      port map(A => \REGMAP_0[29]_net_1\, B => \REGMAP[30]_net_1\, 
        Y => N_2033_0);
    
    \PIPEA1_9_i[7]\ : AND2
      port map(A => DPR(7), B => N_85, Y => N_254);
    
    un1_WDOGRES_0_sqmuxa_0 : OAI21
      port map(A => un1_WDOGRES_0_sqmuxa_0_a2_0_2_i, B => 
        un1_WDOGRES_0_sqmuxa_0_a2_0_3_i, C => N_2431, Y => 
        un1_WDOGRES_0_sqmuxa);
    
    \LB_i_6_0[5]\ : MUX2H
      port map(A => OR_RADDR(3), B => \LB_ADDR[5]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2175);
    
    LB_DOUT_148 : MUX2H
      port map(A => VDB_in(0), B => \LB_DOUT[0]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_148\);
    
    un40_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_681_i, B => N_716, Y => 
        \un40_reg_ads_0_a3_0_a2\);
    
    un2_vsel_2_i_a2_0 : OR2
      port map(A => AMB_c(2), B => AMB_c(5), Y => N_228);
    
    \VDBi_92_iv_0_m2_0[7]\ : MUX2H
      port map(A => N_492, B => N_493, S => \N_441\, Y => N_476);
    
    \VDBi_53_0_iv_2[3]\ : AOI21TTF
      port map(A => \REGMAP[19]_net_1\, B => \REG[172]\, C => 
        \REG_1_m[156]_net_1\, Y => \VDBi_53_0_iv_2[3]_net_1\);
    
    \VDBm_0[13]\ : MUX2H
      port map(A => \PIPEB[13]_net_1\, B => \PIPEA[13]_net_1\, S
         => \BLTCYC_2\, Y => N_2309);
    
    \RAMAD_VME[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_11\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[7]_net_1\);
    
    \VDBi_23[15]\ : MUX2H
      port map(A => \VDBi_18[15]_net_1\, B => \REG[497]\, S => 
        \REGMAP_1[13]_net_1\, Y => \VDBi_23[15]_net_1\);
    
    \VDBi_16_1_a2_3_1[1]\ : NOR2FT
      port map(A => \VDBi_16_1_a2_3_0[1]_net_1\, B => 
        \REGMAP_0[2]_net_1\, Y => N_2512_0);
    
    \LB_s[23]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_102\, CLR => 
        HWRES_c_18, Q => \LB_s[23]_net_1\);
    
    un37_reg_ads_0_a2_4_a2_0 : OR2FT
      port map(A => N_673, B => \VAS[6]_net_1\, Y => N_724);
    
    \RAMDTS[2]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(2), CLR => HWRES_c_21, 
        Q => \RAMDTS[2]_net_1\);
    
    \REG_1[68]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_475\, CLR => 
        \un10_hwres_29\, Q => \REG[68]\);
    
    \TCNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[3]\, CLR => 
        \un10_hwres_33\, Q => \TCNT[3]_net_1\);
    
    \PIPEB_4_i[26]\ : AND2
      port map(A => DPR(26), B => N_616_0, Y => N_2636);
    
    \REG_1_m[167]\ : NAND2
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[167]\, Y => 
        \REG_1_m[167]_net_1\);
    
    \VADm[22]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[22]_net_1\, Y => 
        VADm(22));
    
    un1_LB_DOUT_0_sqmuxa_0_a2_0 : NOR2FT
      port map(A => \REGMAP[10]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_2430);
    
    \REG_i[282]\ : INV
      port map(A => \REG[282]\, Y => REG_i_0_277);
    
    \VDBm_0[14]\ : MUX2H
      port map(A => \PIPEB[14]_net_1\, B => \PIPEA[14]_net_1\, S
         => \BLTCYC_2\, Y => N_2310);
    
    un1_STATE1_29_0_m2 : MUX2H
      port map(A => \STATE1[7]_net_1\, B => \REGMAP_i_0_i[4]\, S
         => \STATE1[8]_net_1\, Y => N_2420);
    
    \STATE5_3[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns[0]\, CLR => 
        HWRES_c_21_0, Q => \STATE5_3[0]_net_1\);
    
    \VDBm[12]\ : MUX2H
      port map(A => N_2308, B => \VDBi[12]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_12);
    
    REG3_123 : MUX2H
      port map(A => \REG[10]\, B => VDB_in(10), S => 
        REG1_0_sqmuxa_0, Y => \REG3_123\);
    
    un43_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_681_i, B => un43_reg_ads_1, Y => 
        \un43_reg_ads_0_a3_0_a2\);
    
    un1_LBUSTMO_1_I_25 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_0[0]\);
    
    \REGMAP[17]\ : DFF
      port map(CLK => CLK_c_c, D => \un57_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_i[17]\);
    
    \REG_i[290]\ : INV
      port map(A => \REG[290]\, Y => REG_i_0_285);
    
    \VDBi_23_d[9]\ : MUX2H
      port map(A => \REG[57]\, B => \REG[491]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23_d[9]_net_1\);
    
    un10_hwres_21 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_21\);
    
    \VDBi_77_0[8]\ : MUX2H
      port map(A => REG_464, B => \REG[449]\, S => 
        \REGMAP_i_i[33]\, Y => N_2060);
    
    \VDBi_92_0_iv[16]\ : OAI21FTT
      port map(A => \VDBi_71[16]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[16]_net_1\, Y => \VDBi_92[16]\);
    
    VAS_66 : MUX2H
      port map(A => \VAS[15]_net_1\, B => VAD_in_14, S => 
        \TST_c_0[1]\, Y => \VAS_66\);
    
    un1_REG_0_sqmuxa_i_a2 : AND2
      port map(A => \STATE5[2]_net_1\, B => un2_nlbrdy_i_0, Y => 
        N_2576_i);
    
    \VDBi_58[15]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[15]\, B => 
        \VDBi_23_m_i[15]\, C => \VDBi_58_0[9]\, Y => 
        \VDBi_58[15]_net_1\);
    
    \REG_1[185]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_225\, CLR => 
        \un10_hwres_11\, Q => \REG[185]\);
    
    un776_regmap_8_0 : OR3
      port map(A => \REGMAP[30]_net_1\, B => \REGMAP[32]_net_1\, 
        C => \REGMAP[0]_net_1\, Y => un776_regmap_8_0_i);
    
    LB_ADDR_553 : MUX2H
      port map(A => \LB_ADDR[10]_net_1\, B => \VAS[10]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_553\);
    
    \VDBm[22]\ : MUX2H
      port map(A => N_2318, B => \VDBi[22]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_22);
    
    REG_1_413 : MUX2H
      port map(A => VDB_in_0(7), B => \REG[448]\, S => N_3104_i, 
        Y => \REG_1_413\);
    
    \LB_i[26]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_538\, CLR => 
        HWRES_c_15, Q => \LB_i[26]_net_1\);
    
    \PIPEB[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_35\, CLR => CLEAR_26, 
        Q => \PIPEB[15]_net_1\);
    
    LB_i_6_sn_m1_0 : XOR2FT
      port map(A => \STATE5[1]_net_1\, B => \STATE5_0[0]_net_1\, 
        Y => LB_i_6_sn_N_2_0);
    
    \VDBi_92_0_iv[27]\ : OAI21FTT
      port map(A => \VDBi_71[27]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[27]_net_1\, Y => \VDBi_92[27]\);
    
    \REG_i[295]\ : INV
      port map(A => \REG[295]\, Y => REG_i_0_290);
    
    PIPEA_615 : MUX2H
      port map(A => \PIPEA_7[26]\, B => \PIPEA[26]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_615\);
    
    \VADm[7]\ : NOR2FT
      port map(A => \PIPEA[7]_net_1\, B => N_2507_0, Y => VADm(7));
    
    \LB_i[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_512\, CLR => 
        HWRES_c_14, Q => \LB_i[0]_net_1\);
    
    \VDBi_53_0_iv_2[6]\ : AOI21TTF
      port map(A => \REGMAP[19]_net_1\, B => \REG[175]\, C => 
        \REG_1_m[159]_net_1\, Y => \VDBi_53_0_iv_2[6]_net_1\);
    
    un1_STATE1_32_0_1 : OA21FTT
      port map(A => N_2408, B => \TST_c_0[2]\, C => N_2451, Y => 
        \un1_STATE1_32_0_1\);
    
    REG_1_304 : MUX2H
      port map(A => VDB_in(26), B => \REG[291]\, S => N_2880_i_0, 
        Y => \REG_1_304\);
    
    \PIPEA_7_i_m2[1]\ : MUX2H
      port map(A => DPR(1), B => \PIPEA1[1]_net_1\, S => N_1996_2, 
        Y => N_510);
    
    \PIPEA_7_r[3]\ : AND2
      port map(A => N_85_2, B => N_512, Y => \PIPEA_7[3]\);
    
    NSELCLK_c_i : INV
      port map(A => \NSELCLK_c\, Y => NSELCLK_c_i_0);
    
    REG_1_137 : MUX2H
      port map(A => \REG[129]\, B => VDB_in(8), S => 
        REG_0_sqmuxa_0, Y => \REG_1_137\);
    
    \VDBi_80[1]\ : MUX2H
      port map(A => \VDBi_71[1]_net_1\, B => \VDBi_80_d[1]_net_1\, 
        S => \VDBi_80_s[2]_net_1\, Y => \VDBi_80[1]_net_1\);
    
    \REG_88[86]\ : NOR2FT
      port map(A => N_2157, B => N_2566, Y => \REG_88[86]_net_1\);
    
    \VDBi_23_m[7]\ : AND2
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[7]_net_1\, Y
         => \VDBi_23_m_i[7]\);
    
    \REGMAP[12]\ : DFF
      port map(CLK => CLK_c_c, D => \un50_reg_ads_0_a2_3_a2\, Q
         => \REGMAP[12]_net_1\);
    
    \REG_1[434]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_399\, CLR => 
        \un10_hwres_23\, Q => \REG[434]\);
    
    REG_1_407 : MUX2H
      port map(A => VDB_in_0(1), B => \REG[442]\, S => N_3104_i, 
        Y => \REG_1_407\);
    
    \LB_DOUT[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_174\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[26]_net_1\);
    
    PIPEA_614 : MUX2H
      port map(A => \PIPEA_7[25]\, B => \PIPEA[25]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_614\);
    
    \VDBi_92_0_iv_0_2[31]\ : AO21TTF
      port map(A => N_792, B => LBSP_in_31, C => 
        \VDBi_92_0_iv_0_0[31]_net_1\, Y => 
        \VDBi_92_0_iv_0_2_i[31]\);
    
    \VDBi_53_0_iv_3[8]\ : AO21TTF
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[161]\, C => 
        \REG_1_m[129]_net_1\, Y => \VDBi_53_0_iv_3_i[8]\);
    
    un64_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_684_i, B => N_689_i, Y => 
        \un64_reg_ads_0_a3_0_a2\);
    
    \REG_1[131]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_139\, CLR => 
        \un10_hwres_8\, Q => \REG[131]\);
    
    \VDBi_92_iv_0_0[7]\ : AOI21TTF
      port map(A => \RAMDTS[7]_net_1\, B => \STATE1_0[1]_net_1\, 
        C => N_596, Y => \VDBi_92_iv_0_0[7]_net_1\);
    
    \PIPEB_4_i_a2_0[0]\ : NAND2
      port map(A => N_428, B => \STATE2_i_0[3]\, Y => N_616_0);
    
    \REG_1_m[155]\ : NAND2
      port map(A => \REGMAP[18]_net_1\, B => \REG[155]\, Y => 
        \REG_1_m[155]_net_1\);
    
    WDOGCLEAR : DFFC
      port map(CLK => CLK_c_c, D => \WDOGCLEAR_69\, CLR => 
        \un10_hwres\, Q => \WDOGCLEAR\);
    
    un1_NRDMEBi_2_sqmuxa_2_i_1 : NAND3
      port map(A => N_79, B => N_2500, C => \STATE2_i_0[3]\, Y
         => un1_NRDMEBi_2_sqmuxa_2_i_1_i);
    
    un2_vsel_2_i_a2 : AND3FFT
      port map(A => N_2434_1, B => N_228, C => AMB_c(1), Y => 
        N_2434_i);
    
    \REG_1_m[200]\ : NAND2
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[200]\, Y => 
        \REG_1_m[200]_net_1\);
    
    \PIPEA[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_614\, CLR => CLEAR_24, 
        Q => \PIPEA[25]_net_1\);
    
    \STATE2_ns_a3_0[0]\ : NOR2FT
      port map(A => \EVREAD_DS\, B => N_426, Y => N_1762);
    
    \PIPEA_7_r[20]\ : AND2
      port map(A => N_85_1, B => N_529, Y => \PIPEA_7[20]\);
    
    \LB_s_m[0]\ : AND2
      port map(A => \LB_s[0]_net_1\, B => N_7_i, Y => 
        \LB_s_m_i[0]\);
    
    un1_LBUSTMO_1_I_14 : XOR2FT
      port map(A => N_66, B => \LBUSTMO_i_0_i[3]\, Y => 
        \DWACT_ADD_CI_0_partial_sum[3]\);
    
    \STATE1[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[2]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1[8]_net_1\);
    
    \VDBi_53_0_iv_0[9]\ : AO21TTF
      port map(A => \REGMAP[12]_net_1\, B => REG_113, C => 
        \REG_1_m[258]_net_1\, Y => \VDBi_53_0_iv_0_i[9]\);
    
    \REGMAP[18]\ : DFF
      port map(CLK => CLK_c_c, D => \un61_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[18]_net_1\);
    
    \STATE2[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE2_ns[4]\, CLR => 
        CLEAR_28, Q => \STATE2[1]_net_1\);
    
    un25_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_681_i, B => un17_reg_ads_1, Y => 
        \un25_reg_ads_0_a3_0_a2\);
    
    un10_hwres_12 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_12\);
    
    LB_ADDR_545 : MUX2H
      port map(A => \LB_ADDR[2]_net_1\, B => \VAS[2]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_545\);
    
    un1_NRDMEBi_2_sqmuxa_1_i_a3_i : OR2
      port map(A => N_584, B => N_1756_1, Y => 
        \un1_NRDMEBi_2_sqmuxa_1_i_a3_i\);
    
    PIPEA1_573 : MUX2H
      port map(A => N_274, B => \PIPEA1[17]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_573\);
    
    un1_STATE2_13_i_0_a2 : NAND3
      port map(A => N_583, B => N_459, C => N_582_1, Y => N_581);
    
    REG_1_402 : MUX2H
      port map(A => VDB_in(28), B => \REG[437]\, S => N_3072_i_0, 
        Y => \REG_1_402\);
    
    un33_reg_ads_0_a2_0_a2_1 : OR2FT
      port map(A => N_685, B => N_662, Y => un33_reg_ads_1);
    
    REG_1_277_e_0 : OR2FT
      port map(A => \REGMAP_0[24]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => N_2816_i_0_0);
    
    un1_STATE2_13_i_0_a2_0_0 : NOR2FT
      port map(A => N_582_1, B => \STATE2[2]_net_1\, Y => 
        \un1_STATE2_13_i_0_a2_0_0\);
    
    \REG_1[420]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_385\, CLR => 
        \un10_hwres_22\, Q => \REG[420]\);
    
    VAS_65 : MUX2H
      port map(A => \VAS[14]_net_1\, B => VAD_in_13, S => 
        \TST_c_0[1]\, Y => \VAS_65\);
    
    REG_1_293 : MUX2H
      port map(A => VDB_in(15), B => \REG[280]\, S => N_2880_i, Y
         => \REG_1_293\);
    
    PIPEA1_567 : MUX2H
      port map(A => N_262, B => \PIPEA1[11]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_567\);
    
    \VDBi[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_627\, CLR => 
        \un10_hwres\, Q => \VDBi[6]_net_1\);
    
    \VDBi_71[18]\ : MUX2H
      port map(A => \VDBi_60[18]_net_1\, B => \REG[427]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[18]_net_1\);
    
    \VDBi_23_m[4]\ : AND2
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[4]_net_1\, Y
         => \VDBi_23_m_i[4]\);
    
    \REG_1[451]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_416\, CLR => 
        \un10_hwres_24\, Q => \REG[451]\);
    
    REG_1_446 : MUX2H
      port map(A => VDB_in(23), B => \REG[505]\, S => N_3170_i_0, 
        Y => \REG_1_446\);
    
    un776_regmap_23 : NOR3
      port map(A => \REGMAP[19]_net_1\, B => \REGMAP[20]_net_1\, 
        C => \un776_regmap_23_0\, Y => \un776_regmap_23\);
    
    \PIPEA1_9_0[29]\ : OR2FT
      port map(A => N_85_0, B => DPR(29), Y => \PIPEA1_9[29]\);
    
    \PIPEA_7_r[18]\ : AND2
      port map(A => N_85_1, B => N_527, Y => \PIPEA_7[18]\);
    
    \VDBi_53_0_iv_1[9]\ : AO21TTF
      port map(A => \REGMAP_i_i[23]\, B => \REG[242]\, C => 
        \REG_1_m[194]_net_1\, Y => \VDBi_53_0_iv_1_i[9]\);
    
    REG_1_463 : MUX2H
      port map(A => VDB_in_0(8), B => \REG[56]\, S => N_3234_i, Y
         => \REG_1_463\);
    
    END_PK_1_0_i_a2_0_a2_0 : NAND2
      port map(A => \EVREAD_DS\, B => \STATE2[1]_net_1\, Y => 
        N_85_0);
    
    PIPEB_47 : MUX2H
      port map(A => \PIPEB[27]_net_1\, B => N_2637, S => N_1996_3, 
        Y => \PIPEB_47\);
    
    \VDBi_66[5]\ : MUX2H
      port map(A => \VDBi_60[5]_net_1\, B => N_2022, S => N_2033, 
        Y => \VDBi_66[5]_net_1\);
    
    REG_1_357_e_0 : OR2FT
      port map(A => \REGMAP_0[29]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_2976_i_0);
    
    \VDBi_92_0_iv_0_0_m2[10]\ : MUX2H
      port map(A => N_490, B => N_2062, S => \N_441\, Y => N_503);
    
    un1_TCNT_1_I_37 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_2_0[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_2_0[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_3_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_1_0[0]\);
    
    \VDBi_66_0[6]\ : MUX2H
      port map(A => \REG[399]\, B => \REG[383]\, S => 
        \REGMAP[29]_net_1\, Y => N_2023);
    
    PIPEA_616 : MUX2H
      port map(A => \PIPEA_7[27]\, B => \PIPEA[27]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_616\);
    
    REG_1_435 : MUX2H
      port map(A => VDB_in_0(12), B => \REG[494]\, S => 
        N_3170_i_1, Y => \REG_1_435\);
    
    REG_1_297 : MUX2H
      port map(A => VDB_in(19), B => \REG[284]\, S => N_2880_i, Y
         => \REG_1_297\);
    
    \VDBi_71[30]\ : MUX2H
      port map(A => \VDBi_60[30]_net_1\, B => \REG[439]\, S => 
        \REGMAP_0[31]_net_1\, Y => \VDBi_71[30]_net_1\);
    
    \LB_i_6_r[23]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_0, C => N_2205, 
        Y => \LB_i_6[23]\);
    
    END_PK_1_0_i_a2_0_a2 : NAND2
      port map(A => \EVREAD_DS\, B => \STATE2[1]_net_1\, Y => 
        N_85);
    
    N_1897 : AO21TTF
      port map(A => N_2565, B => \WRITES\, C => \N_1897_1\, Y => 
        \N_1897\);
    
    \VDBi[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_640\, CLR => 
        \un10_hwres_34\, Q => \VDBi[19]_net_1\);
    
    \REG_i[289]\ : INV
      port map(A => \REG[289]\, Y => REG_i_0_284);
    
    \REG_1[293]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_306\, CLR => 
        \un10_hwres_16\, Q => \REG[293]\);
    
    \FBOUT_m[0]\ : NAND2
      port map(A => FBOUT(0), B => \STATE1[2]_net_1\, Y => 
        \FBOUT_m[0]_net_1\);
    
    \REGMAP_0[24]\ : DFF
      port map(CLK => CLK_c_c, D => \un81_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[24]_net_1\);
    
    \REG3[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_124\, CLR => 
        \un10_hwres_5\, Q => \REG[11]\);
    
    \REG_i[288]\ : INV
      port map(A => \REG[288]\, Y => REG_i_0_283);
    
    OR_RDATA_185 : MUX2H
      port map(A => N_21, B => \OR_RDATA[3]_net_1\, S => N_1832, 
        Y => \OR_RDATA_185\);
    
    \VDBi[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_641\, CLR => 
        \un10_hwres_34\, Q => \VDBi[20]_net_1\);
    
    un5_noe16ri_0_0_a2_0_1 : NOR2FT
      port map(A => \MBLTCYC\, B => \ADACKCYC\, Y => NOEAD_c_1);
    
    \VDBi_92_0_iv_0_0[10]\ : OAI21FTT
      port map(A => N_503, B => N_2613_1, C => 
        \VDBi_92_0_iv_0_0_1[10]_net_1\, Y => \VDBi_92[10]\);
    
    \REG_1_m[162]\ : NAND2
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[162]\, Y => 
        \REG_1_m[162]_net_1\);
    
    VDBi_9_sqmuxa_i_3 : INV
      port map(A => \REGMAP[12]_net_1\, Y => \REGMAP_i_0[12]\);
    
    \REG_1_m[256]\ : NAND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[256]\, Y => 
        \REG_1_m[256]_net_1\);
    
    REG_1_218 : MUX2H
      port map(A => VDB_in(9), B => \REG[178]\, S => N_2720_i_0, 
        Y => \REG_1_218\);
    
    \LB_i_6_1[18]\ : MUX2H
      port map(A => VDB_in(18), B => \LB_DOUT[18]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2200);
    
    LB_i_516 : MUX2H
      port map(A => \LB_i[4]_net_1\, B => \LB_i_6[4]_net_1\, S
         => N_2570, Y => \LB_i_516\);
    
    \LB_i[21]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_533\, CLR => 
        HWRES_c_15, Q => \LB_i[21]_net_1\);
    
    \VDBi_18[24]\ : NAND2
      port map(A => \REG[72]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[24]_net_1\);
    
    CLOSEDTK : DFFC
      port map(CLK => \DS_i_a2\, D => \VCC\, CLR => \TST_c_c[3]\, 
        Q => \CLOSEDTK\);
    
    \VDBi_16_1_a2_1[4]\ : NAND2
      port map(A => N_2512, B => \REG[4]\, Y => N_2471);
    
    \REG_i[505]\ : INV
      port map(A => \REG[505]\, Y => \REG_i[505]_net_1\);
    
    REG_1_439 : MUX2H
      port map(A => VDB_in(16), B => \REG[498]\, S => N_3170_i_1, 
        Y => \REG_1_439\);
    
    \PIPEB[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_24\, CLR => CLEAR_28, 
        Q => \PIPEB[4]_net_1\);
    
    \PIPEA_7_r[14]\ : AND2
      port map(A => N_85_1, B => N_523, Y => \PIPEA_7[14]\);
    
    \VDBi_92_0_iv[8]\ : OAI21FTT
      port map(A => \VDBi_77[8]_net_1\, B => \N_2613_0\, C => 
        \VDBi_92_0_iv_1[8]_net_1\, Y => \VDBi_92[8]\);
    
    REG_1_369 : MUX2H
      port map(A => VDB_in_0(11), B => \REG[404]\, S => 
        N_3008_i_0, Y => \REG_1_369\);
    
    LB_ADDR_548 : MUX2H
      port map(A => \LB_ADDR[5]_net_1\, B => \VAS[5]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_548\);
    
    \VDBi_92_0_iv[20]\ : OAI21FTT
      port map(A => \VDBi_71[20]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[20]_net_1\, Y => \VDBi_92[20]\);
    
    \PULSE_42_f0_i[0]\ : OA21TTF
      port map(A => N_2419, B => \PULSE[0]\, C => 
        \STATE1[7]_net_1\, Y => N_2392);
    
    \REG_1[415]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_380\, CLR => 
        \un10_hwres_21\, Q => \REG[415]\);
    
    \PIPEB_4_i[1]\ : AND2
      port map(A => DPR(1), B => N_616, Y => N_2615);
    
    \LB_DOUT[29]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_177\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[29]_net_1\);
    
    \REG_1[249]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_262\, CLR => 
        \un10_hwres_14\, Q => \REG[249]\);
    
    un1_STATE2_12_0_o2_2_i_a2 : AND3
      port map(A => \PIPEB[30]_net_1\, B => 
        un1_STATE2_12_0_o2_2_i_a2_0_i, C => \PIPEB_i_i[28]\, Y
         => N_652);
    
    un1_LBUSTMO_1_I_6 : NOR2FT
      port map(A => \LBUSTMO[2]_net_1\, B => N_66_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\);
    
    REG3_118 : MUX2H
      port map(A => \REG[5]\, B => VDB_in(5), S => REG1_0_sqmuxa, 
        Y => \REG3_118\);
    
    PIPEB_39 : MUX2H
      port map(A => \PIPEB[19]_net_1\, B => N_2631, S => N_1996_4, 
        Y => \PIPEB_39\);
    
    VDBi_638 : MUX2H
      port map(A => \VDBi_92[17]\, B => \VDBi[17]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_638\);
    
    un1_WDOGRES_0_sqmuxa_0_a2_0_i : AND2
      port map(A => \WDOG[1]_net_1\, B => \WDOG[2]_net_1\, Y => 
        \un1_WDOGRES_0_sqmuxa_0_a2_0_i\);
    
    \LB_s[26]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_105\, CLR => 
        HWRES_c_18, Q => \LB_s[26]_net_1\);
    
    \VDBi_53_0_iv_2[8]\ : AO21TTF
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[193]\, C => 
        \REG_1_m[177]_net_1\, Y => \VDBi_53_0_iv_2_i[8]\);
    
    \REGMAP[14]\ : DFF
      port map(CLK => CLK_c_c, D => \un87_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[14]_net_1\);
    
    \LB_i[15]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_527\, CLR => 
        HWRES_c_14, Q => \LB_i[15]_net_1\);
    
    \VDBi_66[15]\ : MUX2H
      port map(A => \VDBi_60[15]_net_1\, B => N_2032, S => 
        N_2033_0, Y => \VDBi_66[15]_net_1\);
    
    un10_hwres_17 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_1, Y => 
        \un10_hwres_17\);
    
    un43_reg_ads_0_a3_0_a2_0 : OR2
      port map(A => N_666, B => N_662, Y => N_681_i);
    
    \VDBi_66_0[12]\ : MUX2H
      port map(A => \REG[405]\, B => \REG[389]\, S => 
        \REGMAP_0[29]_net_1\, Y => N_2029);
    
    \PIPEA1_9_i[23]\ : AND2
      port map(A => DPR(23), B => N_85_3, Y => N_286);
    
    un10_hwres_1 : OR2
      port map(A => HWRES_c_0_6_0, B => \WDOGTO\, Y => 
        \un10_hwres_1\);
    
    \PIPEB_4_i[3]\ : AND2
      port map(A => DPR(3), B => N_616, Y => N_2617);
    
    VAS_60 : MUX2H
      port map(A => \VAS[9]_net_1\, B => VAD_in_8, S => 
        \TST_c_0[1]\, Y => \VAS_60\);
    
    \REG_1[419]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_384\, SET => 
        \un10_hwres_22\, Q => \REG[419]\);
    
    \LB_DOUT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_152\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[4]_net_1\);
    
    un10_hwres_13 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_13\);
    
    \REG_1[385]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_350\, SET => 
        \un10_hwres_19\, Q => \NSELCLK_c\);
    
    \REG_1[153]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_193\, CLR => 
        \un10_hwres_8_0\, Q => \REG[153]\);
    
    \FBOUT_m[2]\ : NAND2
      port map(A => FBOUT(2), B => \STATE1[2]_net_1\, Y => 
        \FBOUT_m[2]_net_1\);
    
    REG_1_142 : MUX2H
      port map(A => \REG[134]\, B => VDB_in(13), S => 
        REG_0_sqmuxa_0, Y => \REG_1_142\);
    
    \VDBi_71_d[2]\ : MUX2H
      port map(A => N_2019, B => \REG[411]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71_d[2]_net_1\);
    
    \REG_1_m[249]\ : AND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[249]\, Y => 
        \REG_1_m_i[249]\);
    
    \VDBi_53_0_iv_2[15]\ : AOI21TTF
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[184]\, C => 
        \REG_1_m[168]_net_1\, Y => \VDBi_53_0_iv_2[15]_net_1\);
    
    \LB_i_6_r[30]\ : AND3
      port map(A => N_2572_0, B => LB_i_6_sn_N_2_0, C => N_2212, 
        Y => \LB_i_6[30]\);
    
    REG_1_144 : MUX2H
      port map(A => \REG[136]\, B => VDB_in(15), S => 
        REG_0_sqmuxa_0, Y => \REG_1_144\);
    
    un10_hwres_30 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_0, Y => 
        \un10_hwres_30\);
    
    \LB_ADDR[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_548\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[5]_net_1\);
    
    \PIPEB_4_i[27]\ : AND2
      port map(A => DPR(27), B => N_616_0, Y => N_2637);
    
    \PULSE_1[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_242\, CLR => 
        \un10_hwres_4\, Q => \PULSE[7]\);
    
    un10_hwres_7_0 : OR2
      port map(A => HWRES_c_0_0, B => WDOGTO_0, Y => 
        \un10_hwres_7_0\);
    
    \LB_i[28]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_540\, CLR => 
        HWRES_c_16, Q => \LB_i[28]_net_1\);
    
    \PIPEA1_9_i[3]\ : AND2
      port map(A => DPR(3), B => N_85, Y => N_246);
    
    \REG_88_0[83]\ : MUX2H
      port map(A => VDB_in_0(2), B => \REG[83]\, S => N_20, Y => 
        N_2154);
    
    un1_WDOGRES_0_sqmuxa_0_a2_0_a2 : OR3FFT
      port map(A => \STATE1[10]_net_1\, B => N_436, C => 
        \TST_c_0[2]\, Y => N_2431);
    
    \REG_1[86]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_493\, CLR => 
        \un10_hwres_31\, Q => \REG[86]\);
    
    REG_1_268 : MUX2H
      port map(A => VDB_in(6), B => \REG[255]\, S => N_2816_i_0, 
        Y => \REG_1_268\);
    
    \LB_i_6_1[11]\ : MUX2H
      port map(A => VDB_in_0(11), B => \LB_DOUT[11]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2193);
    
    \REG_1[160]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_200\, CLR => 
        \un10_hwres_9\, Q => \REG[160]\);
    
    \PIPEA_7_i_m2[18]\ : MUX2H
      port map(A => DPR(18), B => \PIPEA1[18]_net_1\, S => 
        N_1996_1, Y => N_527);
    
    un2_vsel_1_i : OAI21TTF
      port map(A => \un2_vsel_1_i_a2_0\, B => N_237, C => 
        \TST_c_0[0]\, Y => N_2385);
    
    PIPEB_41 : MUX2H
      port map(A => \PIPEB[21]_net_1\, B => N_2633, S => N_1996_3, 
        Y => \PIPEB_41\);
    
    \REGMAP[2]\ : DFF
      port map(CLK => CLK_c_c, D => \un13_reg_ads_0_a2_0_a2\, Q
         => \REGMAP[2]_net_1\);
    
    PIPEA_601 : MUX2H
      port map(A => \PIPEA_7[12]\, B => \PIPEA[12]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_601\);
    
    \LB_i_6_r[17]\ : AND3
      port map(A => N_2572_2, B => LB_i_6_sn_N_2_1, C => N_2199, 
        Y => \LB_i_6[17]\);
    
    un10_hwres_0 : OR2
      port map(A => HWRES_c_0_6_0, B => \WDOGTO\, Y => 
        \un10_hwres_0\);
    
    \REG3[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_118\, CLR => 
        \un10_hwres_6_0\, Q => \REG[5]\);
    
    END_PK_555 : MUX2H
      port map(A => \END_PK\, B => N_85, S => N_44, Y => 
        \END_PK_555\);
    
    VDBi_9_sqmuxa_1 : NOR3FFT
      port map(A => \REGMAP_i_0[12]\, B => \VDBi_9_sqmuxa_i_0\, C
         => \REGMAP_0[16]_net_1\, Y => \VDBi_9_sqmuxa_1\);
    
    REG_1_392 : MUX2H
      port map(A => VDB_in(18), B => \REG[427]\, S => N_3072_i_1, 
        Y => \REG_1_392\);
    
    \OR_RDATA[1]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_183\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[1]_net_1\);
    
    WDOG_3_I_1 : AND2
      port map(A => \WDOG[0]_net_1\, B => TICK(2), Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    LB_s_100 : MUX2H
      port map(A => LB_in(21), B => \LB_s[21]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_100\);
    
    un10_hwres_18 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_1, Y => 
        \un10_hwres_18\);
    
    \TCNT_10_0_a2[1]\ : AND2
      port map(A => N_2397, B => I_31_1, Y => \TCNT_10[1]\);
    
    \VDBi_53_0_iv_3[1]\ : AO21TTF
      port map(A => \REGMAP[18]_net_1\, B => \REG[154]\, C => 
        \REG_1_m[122]_net_1\, Y => \VDBi_53_0_iv_3_i[1]\);
    
    REG_1_498 : MUX2H
      port map(A => \REG[91]\, B => VDB_in_0(2), S => N_2416_i, Y
         => \REG_1_498\);
    
    \VDBi_92_0_iv_0_a2_4[21]\ : NAND2
      port map(A => N_793, B => \REG[503]\, Y => N_589);
    
    \VDBi_16_1_a2_1[8]\ : NAND2
      port map(A => N_2512, B => \REG[8]\, Y => N_2483);
    
    LB_i_543 : MUX2H
      port map(A => \LB_i[31]_net_1\, B => \LB_i_6[31]\, S => 
        N_2570_0, Y => \LB_i_543\);
    
    REG_1_504 : MUX2H
      port map(A => \REG[97]\, B => VDB_in_0(8), S => N_2416_i, Y
         => \REG_1_504\);
    
    \STATE2_ns_0_0_o2_i[3]\ : INV
      port map(A => \TST_c[2]\, Y => \TST_c_i_0[2]\);
    
    \LB_i_6_1[9]\ : MUX2H
      port map(A => VDB_in_0(9), B => \LB_DOUT[9]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2191);
    
    WDOGRES_71 : MUX2H
      port map(A => \WDOGRES\, B => un1_WDOGRES_0_sqmuxa, S => 
        N_1698, Y => \WDOGRES_71\);
    
    VDBi_633 : MUX2H
      port map(A => \VDBi_92[12]\, B => \VDBi[12]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_633\);
    
    REG_1_396 : MUX2H
      port map(A => VDB_in(22), B => \REG[431]\, S => N_3072_i_0, 
        Y => \REG_1_396\);
    
    PULSE_0_sqmuxa_1_0_a2_0_i2_0_a2_0_a2_2 : OR2FT
      port map(A => \STATE1_0[8]_net_1\, B => \WRITES_0\, Y => 
        PULSE_0_sqmuxa_1_2);
    
    \LB_DOUT[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_165\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[17]_net_1\);
    
    \VDBi_60[5]\ : MUX2H
      port map(A => \VDBi_60_d[5]_net_1\, B => \VDBi_55[5]_net_1\, 
        S => \VDBi_60_s[5]_net_1\, Y => \VDBi_60[5]_net_1\);
    
    \LB_i[13]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_525\, CLR => 
        HWRES_c_14, Q => \LB_i[13]_net_1\);
    
    \REG_1[76]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_483\, CLR => 
        \un10_hwres_30\, Q => \REG[76]\);
    
    \PIPEA1_9_i[17]\ : AND2
      port map(A => DPR(17), B => N_85_4, Y => N_274);
    
    \VDBi_92_iv[0]\ : OR3
      port map(A => \VDBi_80_m_i_i[0]\, B => \VDBi_92_iv_1_i[0]\, 
        C => \LB_s_m_i[0]\, Y => \VDBi_92[0]\);
    
    \REG_1[392]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_357\, CLR => 
        \un10_hwres_20\, Q => \REG[392]\);
    
    un1_NRDMEBi_2_sqmuxa_2_i_a2 : AND2
      port map(A => N_472_i_0, B => \STATE2[2]_net_1\, Y => 
        N_2499_i);
    
    REG_1_357_e : OR2FT
      port map(A => \REGMAP_0[29]_net_1\, B => PULSE_0_sqmuxa_1, 
        Y => N_2976_i);
    
    \PIPEB_4_i[12]\ : AND2
      port map(A => DPR(12), B => N_616_1, Y => N_2626);
    
    \OR_RDATA_5_i_o2_3[0]\ : OR2
      port map(A => N_66_0, B => \STATE5_0[2]_net_1\, Y => 
        N_2572_3);
    
    \REG_1[498]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_439\, SET => 
        \un10_hwres_26\, Q => \REG[498]\);
    
    un94_reg_ads_0_a3_0_a2_1 : NOR2FT
      port map(A => \WRITES_0\, B => N_671, Y => N_685);
    
    \STATE1[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[4]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1[6]_net_1\);
    
    un1_STATE1_34_0_0 : OA21
      port map(A => \STATE1[2]_net_1\, B => 
        un1_STATE1_34_0_a2_1_1_i, C => N_2542, Y => 
        \un1_STATE1_34_0_0\);
    
    \LB_s[21]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_100\, CLR => 
        HWRES_c_18, Q => \LB_s[21]_net_1\);
    
    LB_i_537 : MUX2H
      port map(A => \LB_i[25]_net_1\, B => \LB_i_6[25]\, S => 
        N_2570_0, Y => \LB_i_537\);
    
    \VDBi_71_i_m2[10]\ : MUX2H
      port map(A => \VDBi_66[10]_net_1\, B => \REG[419]\, S => 
        \REGMAP[31]_net_1\, Y => N_490);
    
    \PIPEB_4_i[25]\ : AND2
      port map(A => DPR(25), B => N_616_0, Y => N_229);
    
    \PIPEA_7_i_m2[8]\ : MUX2H
      port map(A => DPR(8), B => \PIPEA1[8]_net_1\, S => N_1996_2, 
        Y => N_517);
    
    \REG_1_m[251]\ : NAND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[251]\, Y => 
        \REG_1_m[251]_net_1\);
    
    \REG_1[172]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_212\, CLR => 
        \un10_hwres_10\, Q => \REG[172]\);
    
    STATE1_tr12_7_0_o2_1 : OR2
      port map(A => \TCNT_i_i[4]\, B => \TCNT[5]_net_1\, Y => 
        STATE1_tr12_7_0_o2_1_i);
    
    \PIPEA_7_i_m2[3]\ : MUX2H
      port map(A => DPR(3), B => \PIPEA1[3]_net_1\, S => N_1996_2, 
        Y => N_512);
    
    un1_anycyc_i_0_o2_i_a2_1 : OR2
      port map(A => \SINGCYC_0\, B => \BLTCYC_0\, Y => N_2507_1);
    
    \REG_1[405]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_370\, CLR => 
        \un10_hwres_21\, Q => \REG[405]\);
    
    \REG_1[396]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_361\, CLR => 
        \un10_hwres_20\, Q => \REG[396]\);
    
    LB_i_6_sn_m1_1 : XOR2FT
      port map(A => \STATE5[1]_net_1\, B => \STATE5_0[0]_net_1\, 
        Y => LB_i_6_sn_N_2_1);
    
    LB_i_530 : MUX2H
      port map(A => \LB_i[18]_net_1\, B => \LB_i_6[18]\, S => 
        N_2570_1, Y => \LB_i_530\);
    
    \REG_m[105]\ : NAND2
      port map(A => \REGMAP[12]_net_1\, B => REG_104, Y => 
        \REG_m[105]_net_1\);
    
    \PIPEB[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_33\, CLR => CLEAR_26, 
        Q => \PIPEB[13]_net_1\);
    
    \REG_1[174]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_214\, CLR => 
        \un10_hwres_10\, Q => \REG[174]\);
    
    PIPEA1_577 : MUX2H
      port map(A => N_282, B => \PIPEA1[21]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_577\);
    
    \VDBi_60_d[5]\ : MUX2H
      port map(A => REG_333, B => L1A_c_c, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60_d[5]_net_1\);
    
    REG_1_486_e_1 : OR2FT
      port map(A => N_2409, B => un1_STATE1_15, Y => N_3234_i_1);
    
    \PIPEA1[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_576\, CLR => CLEAR_21, 
        Q => \PIPEA1[20]_net_1\);
    
    \STATE1_ns_1_iv_0_0[5]\ : OAI21TTF
      port map(A => \SINGCYC\, B => 
        \STATE1_ns_1_iv_0_0_a2_0_0[5]_net_1\, C => N_572_i, Y => 
        \STATE1_ns[5]\);
    
    \VDBi_66[10]\ : MUX2H
      port map(A => \VDBi_60[10]_net_1\, B => N_2027, S => 
        N_2033_0, Y => \VDBi_66[10]_net_1\);
    
    \STATE5_ns_i_0[2]\ : OA21FTT
      port map(A => N_2599_1, B => \LB_REQ_sync\, C => 
        \STATE5_ns_i_0_0_i[2]\, Y => \STATE5_ns_i_0[2]_net_1\);
    
    \VDBi_77_0[13]\ : MUX2H
      port map(A => REG_469, B => \REG[454]\, S => 
        \REGMAP_i_i[33]\, Y => N_2065);
    
    \VDBi_71_i_m2[12]\ : MUX2H
      port map(A => \VDBi_66[12]_net_1\, B => \REG[421]\, S => 
        \REGMAP[31]_net_1\, Y => N_495);
    
    \REG_1[290]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_303\, CLR => 
        \un10_hwres_16\, Q => \REG[290]\);
    
    WDOGTOi_2 : DFFC
      port map(CLK => CLK_c_c, D => \un12_wdog_0_a3\, CLR => 
        un15_hwres_i, Q => WDOGTO_2);
    
    \REG_1[176]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_216\, CLR => 
        \un10_hwres_10\, Q => \REG[176]\);
    
    un1_TCNT_1_I_42 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_3[0]\, B => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_4[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_1_0[0]\);
    
    REG_1_400 : MUX2H
      port map(A => VDB_in(26), B => \REG[435]\, S => N_3072_i_0, 
        Y => \REG_1_400\);
    
    un8_d32_0_a3_0_a2 : AND3FFT
      port map(A => N_656, B => \LWORDS\, C => \VAS[12]_net_1\, Y
         => \un8_d32_0_a3_0_a2\);
    
    REG_1_255 : MUX2H
      port map(A => VDB_in(9), B => \REG[242]\, S => N_2784_i_0, 
        Y => \REG_1_255\);
    
    \VDBi_53_0_iv_3[2]\ : AO21TTF
      port map(A => \REGMAP[16]_net_1\, B => \REG[123]\, C => 
        \VDBi_53_0_iv_2[2]_net_1\, Y => \VDBi_53_0_iv_3_i[2]\);
    
    \REG_1[246]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_259\, SET => 
        \un10_hwres_14\, Q => \REG[246]\);
    
    \LB_i_6_r[25]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_0, C => N_2207, 
        Y => \LB_i_6[25]\);
    
    \STATE2[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE2_ns_i[5]\, CLR => 
        CLEAR_28, Q => \STATE2[0]_net_1\);
    
    PIPEA1_584 : MUX2H
      port map(A => \PIPEA1_9[28]\, B => \PIPEA1[28]_net_1\, S
         => un1_STATE2_13_4_0, Y => \PIPEA1_584\);
    
    \un5_noe16ri_0_0\ : AO21
      port map(A => N_566_1, B => N_436, C => \NOEAD_c_0\, Y => 
        un5_noe16ri_0_0);
    
    REG_1_275 : MUX2H
      port map(A => VDB_in(13), B => \REG[262]\, S => 
        N_2816_i_0_0, Y => \REG_1_275\);
    
    \REG_1[90]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_497\, CLR => 
        \un10_hwres_31\, Q => \REG[90]\);
    
    \REG_1[409]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_374\, CLR => 
        \un10_hwres_21\, Q => \REG[409]\);
    
    REG_1_261_e : OR2FT
      port map(A => \REGMAP_i_i_0[23]\, B => PULSE_0_sqmuxa_1, Y
         => N_2784_i);
    
    \VADm[29]\ : NOR2FT
      port map(A => \PIPEA[29]_net_1\, B => N_2507_0, Y => 
        VADm(29));
    
    REG_1_305 : MUX2H
      port map(A => VDB_in(27), B => \REG[292]\, S => N_2880_i_0, 
        Y => \REG_1_305\);
    
    \VDBi_80[4]\ : MUX2H
      port map(A => \VDBi_77[4]_net_1\, B => REG_476, S => 
        \REGMAP[35]_net_1\, Y => \VDBi_80[4]_net_1\);
    
    \PIPEA_7_r[0]\ : AND2
      port map(A => N_85_3, B => N_509, Y => \PIPEA_7[0]\);
    
    REG_1_sqmuxa_5_i : NAND2
      port map(A => \REGMAP[10]_net_1\, B => \STATE1[8]_net_1\, Y
         => N_20);
    
    \PIPEA[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_612\, CLR => CLEAR_24, 
        Q => \PIPEA[23]_net_1\);
    
    REG_1_130 : MUX2H
      port map(A => \REG[122]\, B => VDB_in(1), S => REG_0_sqmuxa, 
        Y => \REG_1_130\);
    
    \PIPEA1[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_565\, CLR => CLEAR_23, 
        Q => \PIPEA1[9]_net_1\);
    
    un4_asb_NE_0 : OR2
      port map(A => \un4_asb_2\, B => \un4_asb_3\, Y => 
        \un4_asb_NE_0\);
    
    REG_1_416 : MUX2H
      port map(A => VDB_in_0(10), B => \REG[451]\, S => 
        N_3104_i_0, Y => \REG_1_416\);
    
    \REG_1_m[165]\ : NAND2
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[165]\, Y => 
        \REG_1_m[165]_net_1\);
    
    \VADm[23]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[23]_net_1\, Y => 
        VADm(23));
    
    un1_STATE1_34_0 : AO21TTF
      port map(A => N_2535, B => \STATE1[9]_net_1\, C => 
        \un1_STATE1_34_0_0\, Y => un1_STATE1_34);
    
    REG_1_380 : MUX2H
      port map(A => VDB_in_0(6), B => \REG[415]\, S => N_3072_i, 
        Y => \REG_1_380\);
    
    \VDBi_92_0_iv_1[23]\ : AOI21TTF
      port map(A => \LB_s[23]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[23]_net_1\, Y => 
        \VDBi_92_0_iv_1[23]_net_1\);
    
    un1_TCNT_1_I_36 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_1_2[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\);
    
    REG_1_251 : MUX2H
      port map(A => VDB_in(5), B => \REG[238]\, S => N_2784_i, Y
         => \REG_1_251\);
    
    \STATE2_ns_o2_0_0_a2[0]\ : AND2
      port map(A => \REGMAP[0]_net_1\, B => N_436, Y => N_622);
    
    \PIPEA_7_i_m2[10]\ : MUX2H
      port map(A => DPR(10), B => \PIPEA1[10]_net_1\, S => 
        N_1996_1, Y => N_519);
    
    REG_1_271 : MUX2H
      port map(A => VDB_in(9), B => \REG[258]\, S => N_2816_i_0_0, 
        Y => \REG_1_271\);
    
    \VDBi_66_0[9]\ : MUX2H
      port map(A => \REG[402]\, B => \REG[386]\, S => 
        \REGMAP[29]_net_1\, Y => N_2026);
    
    \VDBi_23_m[13]\ : AND2
      port map(A => \VDBi_9_sqmuxa_0\, B => \VDBi_23[13]_net_1\, 
        Y => \VDBi_23_m_i[13]\);
    
    \LB_s[28]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_107\, CLR => 
        HWRES_c_18, Q => \LB_s[28]_net_1\);
    
    un1_STATE1_32_0_o2_0 : OR2FT
      port map(A => \MBLTCYC\, B => N_2507_1, Y => N_2413);
    
    \VDBi_18[28]\ : NAND2
      port map(A => \REG[76]\, B => \TST_c_0[5]\, Y => 
        \VDBi_18[28]_net_1\);
    
    \VDBi_77[4]\ : MUX2H
      port map(A => \VDBi_77_d[4]_net_1\, B => \VDBi_60[4]_net_1\, 
        S => \VDBi_77_s[3]_net_1\, Y => \VDBi_77[4]_net_1\);
    
    REG_1_348 : MUX2H
      port map(A => VDB_in_0(6), B => \REG[383]\, S => N_2976_i, 
        Y => \REG_1_348\);
    
    VDBi_635 : MUX2H
      port map(A => \VDBi_92[14]\, B => \VDBi[14]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_635\);
    
    OR_RDATA_186 : MUX2H
      port map(A => N_2567, B => \OR_RDATA[4]_net_1\, S => N_1832, 
        Y => \OR_RDATA_186\);
    
    REG_1_24_16 : AO21FTT
      port map(A => \WDOGCLEAR\, B => \REG[24]\, C => 
        \un12_wdog_0_a3\, Y => \REG_1_24_16\);
    
    un74_reg_ads_0_a2_0_a2 : OR2FT
      port map(A => \VAS[5]_net_1\, B => N_662, Y => N_198);
    
    PIPEA1_560 : MUX2H
      port map(A => N_248, B => \PIPEA1[4]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_560\);
    
    VDBi_637 : MUX2H
      port map(A => \VDBi_92[16]\, B => \VDBi[16]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_637\);
    
    \VDBi_71[20]\ : MUX2H
      port map(A => \VDBi_60[20]_net_1\, B => \REG[429]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[20]_net_1\);
    
    N_28_i_i_1 : NAND2
      port map(A => N_425, B => N_479, Y => N_2613_1);
    
    un1_STATE2_6_0_a2_0_o2 : OR2
      port map(A => \END_PK\, B => \EVREAD_DS\, Y => N_428);
    
    PURGED : DFFS
      port map(CLK => CLK_c_c, D => \PURGED_14\, SET => 
        N_2371_i_0, Q => \PURGED\);
    
    \LB_i_6_1[29]\ : MUX2H
      port map(A => VDB_in(29), B => \LB_DOUT[29]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2211);
    
    LB_s_103 : MUX2H
      port map(A => LB_in(24), B => \LB_s[24]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_103\);
    
    \TCNT_10_0_a2_1[6]\ : OR3
      port map(A => N_2565, B => N_2455_1, C => 
        \REGMAP[15]_net_1\, Y => N_2455);
    
    \REG_1[435]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_400\, CLR => 
        \un10_hwres_23\, Q => \REG[435]\);
    
    \REG_1[69]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_476\, CLR => 
        \un10_hwres_29\, Q => \REG[69]\);
    
    \VDBm[17]\ : MUX2H
      port map(A => N_2313, B => \VDBi[17]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_17);
    
    \REG_1[265]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_278\, CLR => 
        \un10_hwres_15\, Q => \REG[265]\);
    
    \PIPEA1_9_i[12]\ : AND2
      port map(A => DPR(12), B => N_85_4, Y => N_264);
    
    SINGCYC : DFFC
      port map(CLK => CLK_c_c, D => \SINGCYC_147\, CLR => 
        HWRES_c_21_0, Q => \SINGCYC\);
    
    \VDBm_0[9]\ : MUX2H
      port map(A => \PIPEB[9]_net_1\, B => \PIPEA[9]_net_1\, S
         => \BLTCYC_2\, Y => N_2305);
    
    PIPEA_607 : MUX2H
      port map(A => \PIPEA_7[18]\, B => \PIPEA[18]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_607\);
    
    \FBOUT_m[6]\ : NAND2
      port map(A => FBOUT(6), B => \STATE1[2]_net_1\, Y => 
        \FBOUT_m[6]_net_1\);
    
    \VADm[6]\ : NOR2FT
      port map(A => \PIPEA[6]_net_1\, B => N_2507_0, Y => VADm(6));
    
    un1_STATE1_28_i_a2_1 : NOR3FFT
      port map(A => \STATE1_i_0[8]\, B => 
        \un1_STATE1_28_i_a2_1_0\, C => N_1898, Y => N_2428_i);
    
    \STATE1[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[8]\, CLR => 
        \un10_hwres_32\, Q => \STATE1[2]_net_1\);
    
    \PIPEB[30]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEB_50\, SET => CLEAR_28, 
        Q => \PIPEB[30]_net_1\);
    
    VAS_59 : MUX2H
      port map(A => \VAS[8]_net_1\, B => VAD_in_7, S => 
        \TST_c_0[1]\, Y => \VAS_59\);
    
    CYCSF1_17 : MUX2H
      port map(A => \TST_c_i_0[0]\, B => \CYCSF1\, S => N_2423, Y
         => \CYCSF1_17\);
    
    un10_hwres_29 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_0, Y => 
        \un10_hwres_29\);
    
    REG_1_466 : MUX2H
      port map(A => VDB_in_0(11), B => \REG[59]\, S => N_3234_i_1, 
        Y => \REG_1_466\);
    
    \LB_i_6_1[8]\ : MUX2H
      port map(A => VDB_in_0(8), B => \LB_DOUT[8]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2190);
    
    un1_STATE1_17_0_i : INV
      port map(A => \STATE1[5]_net_1\, Y => \STATE1_i_0[5]\);
    
    \PIPEA_7_i_m2[16]\ : MUX2H
      port map(A => DPR(16), B => \PIPEA1[16]_net_1\, S => 
        N_1996_1, Y => N_525);
    
    un12_wdog_0_a3 : AND3FFT
      port map(A => un12_wdog_0_a3_0_i, B => un12_wdog_0_a3_1_i, 
        C => \un1_WDOGRES_0_sqmuxa_0_a2_0_i\, Y => 
        \un12_wdog_0_a3\);
    
    \REG_1[284]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_297\, CLR => 
        \un10_hwres_16\, Q => \REG[284]\);
    
    \REG_1[439]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_404\, CLR => 
        \un10_hwres_23\, Q => \REG[439]\);
    
    \REG_1[282]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_295\, CLR => 
        \un10_hwres_15\, Q => \REG[282]\);
    
    \REG_1_m[190]\ : NAND2
      port map(A => \REGMAP[20]_net_1\, B => \REG[190]\, Y => 
        \REG_1_m[190]_net_1\);
    
    \LB_i_6_1[4]\ : MUX2H
      port map(A => VDB_in_0(4), B => \LB_DOUT[4]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2186);
    
    \VDBm[27]\ : MUX2H
      port map(A => N_2323, B => \VDBi[27]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_27);
    
    \VDBm[5]\ : MUX2H
      port map(A => N_2301, B => \VDBi[5]_net_1\, S => \SINGCYC\, 
        Y => VDBm_5);
    
    REG_1_394 : MUX2H
      port map(A => VDB_in(20), B => \REG[429]\, S => N_3072_i_1, 
        Y => \REG_1_394\);
    
    \LB_s[12]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_91\, CLR => HWRES_c_17, 
        Q => \LB_s[12]_net_1\);
    
    \REG_i[284]\ : INV
      port map(A => \REG[284]\, Y => REG_i_0_279);
    
    \REG_1[261]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_274\, CLR => 
        \un10_hwres_15\, Q => \REG[261]\);
    
    \REG_1[253]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_266\, CLR => 
        \un10_hwres_14\, Q => \REG[253]\);
    
    \REG_1[444]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_409\, CLR => 
        \un10_hwres_24\, Q => \REG[444]\);
    
    \REG_1_m[196]\ : NAND2
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[196]\, Y => 
        \REG_1_m[196]_net_1\);
    
    \PIPEB[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_20\, CLR => CLEAR_26, 
        Q => \PIPEB[0]_net_1\);
    
    \REG_1[508]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_449\, SET => 
        \un10_hwres_27\, Q => \REG[508]\);
    
    \VDBi_53_0_iv_3[5]\ : AO21TTF
      port map(A => \REGMAP[16]_net_1\, B => \REG_0[126]\, C => 
        \VDBi_53_0_iv_2[5]_net_1\, Y => \VDBi_53_0_iv_3_i[5]\);
    
    WDOG_3_I_23 : XOR2
      port map(A => \WDOG[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => \WDOG_3[3]\);
    
    REG_1_497 : MUX2H
      port map(A => \REG[90]\, B => VDB_in_0(1), S => N_2416_i, Y
         => \REG_1_497\);
    
    un1_STATE2_16_0_0_1 : NAND3FTT
      port map(A => un1_STATE2_16_0_0_0_i, B => N_79, C => N_580, 
        Y => un1_STATE2_16_0);
    
    \LB_s[10]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_89\, CLR => HWRES_c_17, 
        Q => \LB_s[10]_net_1\);
    
    un114_reg_ads_0_a3_0_a2_0 : NOR2
      port map(A => N_664, B => \VAS[3]_net_1\, Y => N_674);
    
    LB_ADDR_550 : MUX2H
      port map(A => \LB_ADDR[7]_net_1\, B => \VAS[7]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_550\);
    
    un78_reg_ads_0_a2_i_o2 : AND2
      port map(A => \VAS[3]_net_1\, B => \VAS[4]_net_1\, Y => 
        N_463);
    
    \VDBi_53_0_iv[1]\ : AO21TTF
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[1]_net_1\, C
         => \VDBi_53_0_iv_6[1]_net_1\, Y => \VDBi_53[1]\);
    
    un1_LBUSTMO_1_I_12 : XOR2FT
      port map(A => N_66, B => \LBUSTMO_i_0_i[3]\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\);
    
    \VDBi_23[28]\ : MUX2H
      port map(A => \VDBi_18[28]_net_1\, B => \REG_i[510]_net_1\, 
        S => \REGMAP_0[13]_net_1\, Y => \VDBi_23[28]_net_1\);
    
    un1_STATE5_18_i_0 : NAND2
      port map(A => N_1837, B => N_2608, Y => N_1832);
    
    \REG_i[399]\ : INV
      port map(A => \REG[399]\, Y => REG_i_0_394);
    
    \REG_1[378]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_343\, CLR => 
        \un10_hwres_18\, Q => \REG[378]\);
    
    \REG_1[257]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_270\, CLR => 
        \un10_hwres_14\, Q => \REG[257]\);
    
    \REG_1[394]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_359\, CLR => 
        \un10_hwres_20\, Q => \REG[394]\);
    
    \LB_i[16]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_528\, CLR => 
        HWRES_c_14, Q => \LB_i[16]_net_1\);
    
    \LB_i[3]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_515\, CLR => 
        HWRES_c_16, Q => \LB_i[3]_net_1\);
    
    \LB_DOUT[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_163\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[15]_net_1\);
    
    \VDBi_92_0_iv[19]\ : OAI21FTT
      port map(A => \VDBi_71[19]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[19]_net_1\, Y => \VDBi_92[19]\);
    
    REG_1_327 : MUX2H
      port map(A => VDB_in(17), B => \REG[362]\, S => N_2944_i, Y
         => \REG_1_327\);
    
    un10_hwres_11 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_11\);
    
    REG_1_421 : MUX2H
      port map(A => VDB_in_0(15), B => \REG[456]\, S => 
        N_3104_i_0, Y => \REG_1_421\);
    
    \VDBi_92_0_iv_0_a2_11[21]\ : NOR2FT
      port map(A => \REGMAP_0[13]_net_1\, B => N_680, Y => N_793);
    
    \STATE5_ns_i_0_0[2]\ : OA21FTT
      port map(A => N_1861, B => \STATE5_0[2]_net_1\, C => 
        N_2593_i, Y => \STATE5_ns_i_0_0_i[2]\);
    
    \VDBi_53_0_iv_5[0]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[0]\, B => \REG_1_m_i[233]\, 
        C => \REG_1_m_i[249]\, Y => \VDBi_53_0_iv_5_i[0]\);
    
    \REG_1[497]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_438\, CLR => 
        \un10_hwres_26\, Q => \REG[497]\);
    
    REG_1_381 : MUX2H
      port map(A => VDB_in_0(7), B => \REG[416]\, S => N_3072_i, 
        Y => \REG_1_381\);
    
    \REG_1[19]\ : DFFC
      port map(CLK => ALICLK_c, D => \REG_1_19_70\, CLR => 
        HWRES_c_21, Q => \REG[19]\);
    
    \VDBi_71_s[1]\ : OR2FT
      port map(A => \VDBi_66_s[1]_net_1\, B => 
        \REGMAP_0[31]_net_1\, Y => \VDBi_71_s[1]_net_1\);
    
    \PIPEA1[29]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEA1_585\, SET => CLEAR_22, 
        Q => \PIPEA1[29]_net_1\);
    
    REG_1_492 : MUX2H
      port map(A => \REG_88[85]_net_1\, B => \REG[85]\, S => 
        un1_STATE1_15, Y => \REG_1_492\);
    
    LB_i_535 : MUX2H
      port map(A => \LB_i[23]_net_1\, B => \LB_i_6[23]\, S => 
        N_2570_0, Y => \LB_i_535\);
    
    \VDBi_92_0_iv_0[13]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[13]_net_1\, C
         => \PIPEA_m[13]_net_1\, Y => \VDBi_92_0_iv_0[13]_net_1\);
    
    \VDBi_16_1_a2_0[11]\ : AND2
      port map(A => N_2512_0, B => \REG[11]\, Y => N_2489_i);
    
    N_77_i_i_o2_1_0 : NAND2
      port map(A => \PIPEA[30]_net_1\, B => \PIPEA_i_0_i[28]\, Y
         => \N_77_i_i_o2_1_0\);
    
    \LB_DOUT[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_168\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[20]_net_1\);
    
    \VDBi_77[13]\ : MUX2H
      port map(A => \VDBi_71[13]_net_1\, B => N_2065, S => 
        N_441_0, Y => \VDBi_77[13]_net_1\);
    
    \STATE1_ns_1_iv_0_a2_0[3]\ : OAI21
      port map(A => N_2533, B => \WRITES_1\, C => 
        \STATE1_0[8]_net_1\, Y => N_2545);
    
    \REG_i[511]\ : INV
      port map(A => \REG[511]\, Y => \REG_i[511]_net_1\);
    
    \PIPEB[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_36\, CLR => CLEAR_26, 
        Q => \PIPEB[16]_net_1\);
    
    REG_1_350 : MUX2H
      port map(A => VDB_in_0(8), B => \NSELCLK_c\, S => 
        N_2976_i_0, Y => \REG_1_350\);
    
    \VDBi_92_0_iv[13]\ : OAI21FTT
      port map(A => \VDBi_77[13]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[13]_net_1\, Y => \VDBi_92[13]\);
    
    \LB_i_6_1[20]\ : MUX2H
      port map(A => VDB_in(20), B => \LB_DOUT[20]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2202);
    
    REG_1_370 : MUX2H
      port map(A => VDB_in_0(12), B => \REG[405]\, S => 
        N_3008_i_0, Y => \REG_1_370\);
    
    \VDBm_0[5]\ : MUX2H
      port map(A => \PIPEB[5]_net_1\, B => \PIPEA[5]_net_1\, S
         => \BLTCYC\, Y => N_2301);
    
    \REGMAP[31]\ : DFF
      port map(CLK => CLK_c_c, D => \un111_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[31]_net_1\);
    
    DSS : DFFS
      port map(CLK => CLK_c_c, D => \DSSF1\, SET => HWRES_c_13, Q
         => \TST_c[2]\);
    
    \VDBi_23[20]\ : MUX2H
      port map(A => \VDBi_18[20]_net_1\, B => \REG_i[502]_net_1\, 
        S => \REGMAP_1[13]_net_1\, Y => \VDBi_23[20]_net_1\);
    
    \VDBi_55[2]\ : MUX2H
      port map(A => \VDBi_53[2]\, B => SPULSE2_c_c, S => 
        \REGMAP[26]_net_1\, Y => \VDBi_55[2]_net_1\);
    
    REG_1_249 : MUX2H
      port map(A => VDB_in(3), B => \REG[236]\, S => N_2784_i, Y
         => \REG_1_249\);
    
    \REG_1[100]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_507\, CLR => 
        \un10_hwres_7\, Q => \REG[100]\);
    
    \VDBi_92_0_iv[28]\ : OAI21FTT
      port map(A => \VDBi_71[28]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[28]_net_1\, Y => \VDBi_92[28]\);
    
    \VDBi_77_0[3]\ : MUX2H
      port map(A => REG_459, B => \REG[444]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_2055);
    
    \VDBi_60[18]\ : MUX2H
      port map(A => \VDBi_55[18]_net_1\, B => LBSP_in_18, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[18]_net_1\);
    
    RAMAD_VME_6 : MUX2H
      port map(A => \VAS[3]_net_1\, B => \RAMAD_VME[2]_net_1\, S
         => \TCNT_0_sqmuxa_i_s\, Y => \RAMAD_VME_6\);
    
    REG_1_235 : MUX2H
      port map(A => VDB_in(10), B => \REG[195]\, S => N_2752_i_0, 
        Y => \REG_1_235\);
    
    \REG_1[492]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_433\, SET => 
        \un10_hwres_26\, Q => \REG[492]\);
    
    \REG_m[113]\ : NAND2
      port map(A => \REGMAP[12]_net_1\, B => REG_112, Y => 
        \REG_m[113]_net_1\);
    
    WDOG_3_I_31 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \WDOG[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    \VDBi_92_0_iv_0[31]\ : OR3
      port map(A => \VDBi_92_0_iv_0_4_i[31]\, B => 
        \VDBi_92_0_iv_0_2_i[31]\, C => \VDBi_92_0_iv_0_1_i[31]\, 
        Y => \VDBi_92[31]\);
    
    un1_STATE1_34_0_0_0 : AO21TTF
      port map(A => N_2535, B => \STATE1_0[9]_net_1\, C => 
        \un1_STATE1_34_0_0\, Y => \un1_STATE1_34_0\);
    
    \REG_1[67]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_474\, CLR => 
        \un10_hwres_29\, Q => \REG[67]\);
    
    \PIPEB_4_i[24]\ : AND2
      port map(A => DPR(24), B => N_616_0, Y => N_2635);
    
    \PIPEA[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_615\, CLR => CLEAR_24, 
        Q => \PIPEA[26]_net_1\);
    
    \VDBi_71_s_0[1]\ : NOR2
      port map(A => \REGMAP[27]_net_1\, B => \VDBi_71_s[1]_net_1\, 
        Y => \VDBi_71_s_0[1]_net_1\);
    
    VDBi_641 : MUX2H
      port map(A => \VDBi_92[20]\, B => \VDBi[20]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_641\);
    
    \VDBi_23_m[11]\ : AND2
      port map(A => \VDBi_9_sqmuxa_0\, B => \VDBi_23[11]_net_1\, 
        Y => \VDBi_23_m_i[11]\);
    
    \REG_88_0[84]\ : MUX2H
      port map(A => VDB_in_0(3), B => \REG[84]\, S => N_20, Y => 
        N_2155);
    
    \VDBi_92_iv_1[1]\ : AOI21TTF
      port map(A => N_457_i_0, B => \PIPEA[1]_net_1\, C => 
        \VDBi_92_iv_0[1]_net_1\, Y => \VDBi_92_iv_1[1]_net_1\);
    
    \VADm[12]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[12]_net_1\, Y => VADm(12));
    
    LB_ADDR_549 : MUX2H
      port map(A => \LB_ADDR[6]_net_1\, B => \VAS[6]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_549\);
    
    \REG_i[512]\ : INV
      port map(A => \REG[512]\, Y => \REG_i[512]_net_1\);
    
    un17_reg_ads_0_a3_0_a2_1 : OR2FT
      port map(A => \VAS[3]_net_1\, B => N_694, Y => 
        un17_reg_ads_1);
    
    \STATE2[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE2_ns[3]\, CLR => 
        CLEAR_28, Q => \STATE2[2]_net_1\);
    
    REG_1_231 : MUX2H
      port map(A => VDB_in(6), B => \REG[191]\, S => N_2752_i, Y
         => \REG_1_231\);
    
    \REG_1[423]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_388\, CLR => 
        \un10_hwres_22\, Q => \REG[423]\);
    
    \REG_i[498]\ : INV
      port map(A => \REG[498]\, Y => \REG_i[498]_net_1\);
    
    \REG_i[394]\ : INV
      port map(A => \REG[394]\, Y => REG_i_0_389);
    
    REG_1_195 : MUX2H
      port map(A => VDB_in(2), B => \REG[155]\, S => N_2688_i, Y
         => \REG_1_195\);
    
    REG_1_510 : MUX2H
      port map(A => \REG[103]\, B => VDB_in_0(14), S => N_2416_i, 
        Y => \REG_1_510\);
    
    un1_EVREAD_DS_1_sqmuxa_1_0 : OR2FT
      port map(A => N_426, B => N_86, Y => 
        un1_EVREAD_DS_1_sqmuxa_1);
    
    \REG_i[292]\ : INV
      port map(A => \REG[292]\, Y => REG_i_0_287);
    
    \VDBi[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_625\, CLR => 
        \un10_hwres_35\, Q => \VDBi[4]_net_1\);
    
    REG_1_204 : MUX2H
      port map(A => VDB_in(11), B => \REG[164]\, S => N_2688_i_0, 
        Y => \REG_1_204\);
    
    un1_TCNT_1_I_39 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_1_1[0]\, B => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_2_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    REG_1_202 : MUX2H
      port map(A => VDB_in(9), B => \REG[162]\, S => N_2688_i_0, 
        Y => \REG_1_202\);
    
    \VDBi_92_iv_1[3]\ : AOI21TTF
      port map(A => N_457_i_0, B => \PIPEA[3]_net_1\, C => 
        \VDBi_92_iv_0[3]_net_1\, Y => \VDBi_92_iv_1[3]_net_1\);
    
    \REG_1[178]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_218\, CLR => 
        \un10_hwres_11\, Q => \REG[178]\);
    
    \VDBi_23[6]\ : MUX2H
      port map(A => N_491, B => \REG[488]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23[6]_net_1\);
    
    \PIPEA_7_r[4]\ : AND2
      port map(A => N_85_2, B => N_513, Y => \PIPEA_7[4]\);
    
    un1_STATE1_17_0_o2_i_o2 : NOR2
      port map(A => \STATE1[4]_net_1\, B => \STATE1[6]_net_1\, Y
         => N_462);
    
    \VDBi_18[19]\ : AND2
      port map(A => \REG[67]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[19]_net_1\);
    
    \VDBi_53_0_iv_3[4]\ : AO21TTF
      port map(A => \REGMAP[16]_net_1\, B => \REG_0[125]\, C => 
        \VDBi_53_0_iv_2[4]_net_1\, Y => \VDBi_53_0_iv_3_i[4]\);
    
    un1_noe16wi_i_s_0 : OR2FT
      port map(A => N_436, B => \WRITES_1\, Y => \NOE16W_c\);
    
    REG3_120 : MUX2H
      port map(A => \REG[7]\, B => VDB_in(7), S => REG1_0_sqmuxa, 
        Y => \REG3_120\);
    
    \TCNT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[5]\, CLR => 
        \un10_hwres_33\, Q => \TCNT[5]_net_1\);
    
    \LB_i_6_1[6]\ : MUX2H
      port map(A => VDB_in_0(6), B => \LB_DOUT[6]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2188);
    
    \REG_1_m[261]\ : NAND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[261]\, Y => 
        \REG_1_m[261]_net_1\);
    
    \RAMAD_VME[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_10\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[6]_net_1\);
    
    \REG_88_0[85]\ : MUX2H
      port map(A => VDB_in_0(4), B => \REG[85]\, S => N_20, Y => 
        N_2156);
    
    END_PK_1_0_i_a2_0_a2_3 : NAND2
      port map(A => \EVREAD_DS\, B => \STATE2[1]_net_1\, Y => 
        N_85_3);
    
    \VDBi_92_0_iv_0[23]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[23]_net_1\, C
         => \PIPEA_m[23]_net_1\, Y => \VDBi_92_0_iv_0[23]_net_1\);
    
    \LB_i[11]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_523\, CLR => 
        HWRES_c_14, Q => \LB_i[11]_net_1\);
    
    \VDBi_55[16]\ : NOR2
      port map(A => \REGMAP[26]_net_1\, B => \VDBi_23[16]_net_1\, 
        Y => \VDBi_55[16]_net_1\);
    
    nLBRD_146 : MUX2H
      port map(A => \NLBRD_c\, B => N_1837, S => N_2569, Y => 
        \nLBRD_146\);
    
    REG3_114 : MUX2H
      port map(A => \REG[1]\, B => VDB_in(1), S => REG1_0_sqmuxa, 
        Y => \REG3_114\);
    
    RAMAD_VME_4 : MUX2H
      port map(A => \VAS[1]_net_1\, B => \RAMAD_VME[0]_net_1\, S
         => \TCNT_0_sqmuxa_i_s\, Y => \RAMAD_VME_4\);
    
    \REG_1[195]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_235\, CLR => 
        \un10_hwres_12\, Q => \REG[195]\);
    
    \REG_1[360]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_325\, CLR => 
        \un10_hwres_17\, Q => \REG[360]\);
    
    PIPEA1_570 : MUX2H
      port map(A => N_268, B => \PIPEA1[14]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_570\);
    
    \VDBi_80_m_0[0]\ : MUX2H
      port map(A => d_m7, B => \VDBi_66[0]_net_1\, S => 
        \VDBi_80_m_0_m4_0_a2\, Y => \VDBi_80_m_i_i[0]\);
    
    \REGMAP_1[8]\ : DFF
      port map(CLK => CLK_c_c, D => \un37_reg_ads_0_a2_4_a2\, Q
         => \TST_c_1[5]\);
    
    \OR_RDATA_5_i_o2_2[0]\ : OR2
      port map(A => N_66_0, B => \STATE5_0[2]_net_1\, Y => 
        N_2572_2);
    
    LB_s_95 : MUX2H
      port map(A => LB_in(16), B => \LB_s[16]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_95\);
    
    \PULSE_1[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_241\, CLR => 
        \un10_hwres_4\, Q => \PULSE[6]\);
    
    un1_EVREAD_DS_1_sqmuxa_1_0_a2_2_a2 : OA21TTF
      port map(A => N_440, B => N_665, C => N_725, Y => N_86);
    
    \VDBi[29]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_650\, CLR => 
        \un10_hwres_35\, Q => \VDBi[29]_net_1\);
    
    WRITES : DFFC
      port map(CLK => CLK_c_c, D => \WRITES_2\, CLR => HWRES_c_23, 
        Q => \WRITES\);
    
    PIPEA1_565 : MUX2H
      port map(A => N_258, B => \PIPEA1[9]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_565\);
    
    \LB_i_6_r[12]\ : AND3
      port map(A => N_2572_2, B => LB_i_6_sn_N_2_1, C => N_2194, 
        Y => \LB_i_6[12]\);
    
    \VDBi_77_0[11]\ : MUX2H
      port map(A => REG_467, B => \REG[452]\, S => 
        \REGMAP_i_i[33]\, Y => N_2063);
    
    un1_NRDMEBi_2_sqmuxa_2_i_a2_1 : NOR3
      port map(A => N_583, B => N_426, C => N_428, Y => N_7139_i);
    
    DSSF1_13 : MUX2H
      port map(A => DSSF1_2, B => \DSSF1\, S => N_2421, Y => 
        \DSSF1_13\);
    
    \VDBi_77_d[3]\ : MUX2H
      port map(A => \VDBi_71_d[3]_net_1\, B => N_2055, S => 
        \N_441\, Y => \VDBi_77_d[3]_net_1\);
    
    LB_i_539 : MUX2H
      port map(A => \LB_i[27]_net_1\, B => \LB_i_6[27]\, S => 
        N_2570_0, Y => \LB_i_539\);
    
    \VDBi_53_0_iv_5[12]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[12]\, B => 
        \VDBi_53_0_iv_0_i[12]\, C => \VDBi_53_0_iv_1_i[12]\, Y
         => \VDBi_53_0_iv_5_i[12]\);
    
    \STATE1_ns_1_iv_0_1[3]\ : AND3
      port map(A => N_2544, B => N_2545, C => N_2542, Y => 
        \STATE1_ns_1_iv_0_1[3]_net_1\);
    
    \REGMAP[21]\ : DFF
      port map(CLK => CLK_c_c, D => \un70_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[21]_net_1\);
    
    \VDBi_23[7]\ : MUX2H
      port map(A => \VDBi_16[7]\, B => \VDBi_23_d[7]_net_1\, S
         => \VDBi_23_s[7]_net_1\, Y => \VDBi_23[7]_net_1\);
    
    \RAMAD_VME[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_5\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[1]_net_1\);
    
    \PIPEA_m[28]\ : NAND2
      port map(A => N_457_i_0_0, B => \PIPEA_i_0_i[28]\, Y => 
        \PIPEA_m[28]_net_1\);
    
    \VDBi_53_0_iv_3[12]\ : AO21TTF
      port map(A => \REGMAP_0[16]_net_1\, B => \REG[133]\, C => 
        \VDBi_53_0_iv_2[12]_net_1\, Y => \VDBi_53_0_iv_3_i[12]\);
    
    \VDBi_60[15]\ : MUX2H
      port map(A => \VDBi_58[15]_net_1\, B => LBSP_in_15, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[15]_net_1\);
    
    \VDBi_92_0_iv_0_m2[12]\ : MUX2H
      port map(A => N_495, B => N_496, S => N_441_0, Y => N_502);
    
    \VDBi_92_iv_0[2]\ : AOI21TTF
      port map(A => \RAMDTS[2]_net_1\, B => \STATE1[1]_net_1\, C
         => \FBOUT_m[2]_net_1\, Y => \VDBi_92_iv_0[2]_net_1\);
    
    \REG_1[130]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_138\, CLR => 
        \un10_hwres_8\, Q => \REG[130]\);
    
    \REG_1[250]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_263\, CLR => 
        \un10_hwres_14\, Q => \REG[250]\);
    
    \VDBi_16_1_a2_2_0[1]\ : NOR2FT
      port map(A => \REGMAP[6]_net_1\, B => \REGMAP_0[2]_net_1\, 
        Y => N_2511_0);
    
    PIPEA_613 : MUX2H
      port map(A => \PIPEA_7[24]\, B => \PIPEA[24]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_613\);
    
    \VDBi_80[2]\ : MUX2H
      port map(A => \VDBi_71[2]_net_1\, B => \VDBi_80_d[2]_net_1\, 
        S => \VDBi_80_s[2]_net_1\, Y => \VDBi_80[2]_net_1\);
    
    nLBLAST : DFFS
      port map(CLK => ALICLK_c, D => \nLBLAST_112\, SET => 
        HWRES_c_23, Q => \NLBLAST_c\);
    
    \VDBi_92_0_iv_0_0_1[10]\ : AOI21TTF
      port map(A => \LB_s[10]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0_0_0[10]_net_1\, Y => 
        \VDBi_92_0_iv_0_0_1[10]_net_1\);
    
    \VDBi_23_m_i_0[12]\ : AND2
      port map(A => N_494, B => \VDBi_9_sqmuxa_0\, Y => N_412_i);
    
    \STATE1_0[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[8]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1_0[2]_net_1\);
    
    \STATE2_ns_0[0]\ : AO21
      port map(A => N_1756, B => \STATE2[5]_net_1\, C => N_1762, 
        Y => \STATE2_ns[0]\);
    
    REG_1_351 : MUX2H
      port map(A => VDB_in_0(9), B => \REG[386]\, S => N_2976_i_0, 
        Y => \REG_1_351\);
    
    un1_STATE2_12_0_0_o2 : OR2
      port map(A => \STATE2[0]_net_1\, B => \STATE2[5]_net_1\, Y
         => N_485);
    
    REG_1_371 : MUX2H
      port map(A => VDB_in_0(13), B => \REG[406]\, S => 
        N_3008_i_0, Y => \REG_1_371\);
    
    \REG_1[483]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_424\, CLR => 
        \un10_hwres_25\, Q => \REG[483]\);
    
    \VAS[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_66\, CLR => HWRES_c_22_0, 
        Q => \VAS[15]_net_1\);
    
    \RAMAD_VME[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_8\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[4]_net_1\);
    
    \VDBi_55[28]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[28]_net_1\, Y => \VDBi_55[28]_net_1\);
    
    \VDBi_92_0_iv_0_a2_0[12]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[12]_net_1\, Y => 
        N_599);
    
    \LB_i[27]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_539\, CLR => 
        HWRES_c_15, Q => \LB_i[27]_net_1\);
    
    \VDBi_66_0[4]\ : MUX2H
      port map(A => \REG[397]\, B => \REG[381]\, S => 
        \REGMAP[29]_net_1\, Y => N_2021);
    
    \VAS[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_54\, CLR => HWRES_c_22_0, 
        Q => \VAS[3]_net_1\);
    
    \REG_1[506]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_447\, SET => 
        \un10_hwres_27\, Q => \REG[506]\);
    
    \REG_1_m[122]\ : NAND2
      port map(A => \REGMAP[16]_net_1\, B => \REG[122]\, Y => 
        \REG_1_m[122]_net_1\);
    
    \LB_i[18]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_530\, CLR => 
        HWRES_c_15, Q => \LB_i[18]_net_1\);
    
    un1_TCNT_1_I_24 : XOR2
      port map(A => \TCNT_i_i[4]\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[4]\);
    
    \VDBi_80_d[2]\ : MUX2H
      port map(A => N_2054, B => REG_474, S => \REGMAP[35]_net_1\, 
        Y => \VDBi_80_d[2]_net_1\);
    
    END_PK_1_0_i_a2_0_a2_1 : NAND2
      port map(A => \EVREAD_DS\, B => \STATE2[1]_net_1\, Y => 
        N_85_1);
    
    \VDBi_55[5]\ : OA21TTF
      port map(A => \VDBi_23_m_i[5]\, B => \VDBi_53_0_iv_5_i[5]\, 
        C => \REGMAP[26]_net_1\, Y => \VDBi_55[5]_net_1\);
    
    LB_REQ : DFFC
      port map(CLK => CLK_c_c, D => \LB_REQ_67\, CLR => 
        \un10_hwres_3\, Q => \LB_REQ\);
    
    \WDOG_i[5]\ : AO21
      port map(A => \WDOGRES\, B => WDOGRES1_i, C => HWRES_c_1, Y
         => un15_hwres_i);
    
    un105_reg_ads_0_a3_0_a2_1_0 : OR2
      port map(A => N_672, B => N_671, Y => un105_reg_ads_1_0);
    
    \PIPEB_4_i[2]\ : AND2
      port map(A => DPR(2), B => N_616, Y => N_2616);
    
    \STATE5_ns_0_0_a2[1]\ : NAND3
      port map(A => N_2606_i_i, B => \STATE5[2]_net_1\, C => 
        \REQUESTER\, Y => N_2595);
    
    PIPEA1_561 : MUX2H
      port map(A => N_250, B => \PIPEA1[5]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_561\);
    
    \REG_i[502]\ : INV
      port map(A => \REG[502]\, Y => \REG_i[502]_net_1\);
    
    REG_1_246 : MUX2H
      port map(A => VDB_in(0), B => \REG[233]\, S => N_2784_i, Y
         => \REG_1_246\);
    
    VDBi_622 : MUX2H
      port map(A => \VDBi_92[1]\, B => \VDBi[1]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_622\);
    
    \STATE1_0[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[3]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1_0[7]_net_1\);
    
    \OR_RDATA_5_i_o2_i[0]\ : INV
      port map(A => \STATE5[2]_net_1\, Y => \STATE5_i_0[2]\);
    
    \STATE1[0]\ : DFFC
      port map(CLK => CLK_c_c, D => N_43, CLR => \un10_hwres_32\, 
        Q => \STATE1[0]_net_1\);
    
    REG_1_368 : MUX2H
      port map(A => VDB_in_0(10), B => \REG[403]\, S => 
        N_3008_i_0, Y => \REG_1_368\);
    
    \REGMAP_0[31]\ : DFF
      port map(CLK => CLK_c_c, D => \un111_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[31]_net_1\);
    
    PIPEA1_556 : MUX2H
      port map(A => N_238, B => \PIPEA1[0]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_556\);
    
    un1_STATE5_18_i_0_a2 : OR2FT
      port map(A => \STATE5_0[2]_net_1\, B => \REQUESTER\, Y => 
        N_2608);
    
    \VDBi_23_i_0_m2[12]\ : MUX2H
      port map(A => N_497, B => \REG[494]\, S => 
        \REGMAP_1[13]_net_1\, Y => N_494);
    
    \LB_i_6_0[7]\ : MUX2H
      port map(A => OR_RADDR(5), B => \LB_ADDR[7]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2177);
    
    un94_reg_ads_0_a3_0_a2_0 : NOR2FT
      port map(A => \VAS[3]_net_1\, B => N_664, Y => N_682);
    
    REG_1_383 : MUX2H
      port map(A => VDB_in_0(9), B => \REG[418]\, S => N_3072_i, 
        Y => \REG_1_383\);
    
    \VDBi_16_1_a2_0[6]\ : AND2
      port map(A => N_2511, B => REG_37, Y => N_2476_i);
    
    \VDBi[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_623\, CLR => 
        \un10_hwres_35\, Q => \VDBi[2]_net_1\);
    
    \STATE1[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[9]\, CLR => 
        \un10_hwres_32\, Q => \STATE1[1]_net_1\);
    
    \REG_1[389]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_354\, CLR => 
        \un10_hwres_19\, Q => \REG[389]\);
    
    \REG_1_m[198]\ : NAND2
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[198]\, Y => 
        \REG_1_m[198]_net_1\);
    
    \VDBm_0[31]\ : MUX2H
      port map(A => \PIPEB[31]_net_1\, B => \PIPEA[31]_net_1\, S
         => \BLTCYC_0\, Y => N_2327);
    
    \PIPEB[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_37\, CLR => CLEAR_26, 
        Q => \PIPEB[17]_net_1\);
    
    \STATE2_ns_0_0_a2[4]\ : OR2FT
      port map(A => \STATE2[1]_net_1\, B => \TST_c_0[2]\, Y => 
        N_580);
    
    \PIPEB_4_i[5]\ : AND2
      port map(A => DPR(5), B => N_616, Y => N_2619);
    
    LB_DOUT_165 : MUX2H
      port map(A => VDB_in(17), B => \LB_DOUT[17]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_165\);
    
    \VADm[28]\ : NOR2FT
      port map(A => \PIPEA_i_0_i[28]\, B => N_2507_0, Y => 
        VADm(28));
    
    REG_1_330 : MUX2H
      port map(A => VDB_in(20), B => \REG[365]\, S => N_2944_i, Y
         => \REG_1_330\);
    
    un776_regmap_25 : NAND3
      port map(A => \un776_regmap_23\, B => \VDBi_9_sqmuxa_i_1\, 
        C => \VDBi_9_sqmuxa_i_0\, Y => un776_regmap_25_i);
    
    \VDBi_53_0_iv_5[13]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[13]\, B => 
        \VDBi_53_0_iv_0_i[13]\, C => \VDBi_53_0_iv_1_i[13]\, Y
         => \VDBi_53_0_iv_5_i[13]\);
    
    \PIPEB_4_i[31]\ : AND2
      port map(A => N_616_0, B => DPR(31), Y => N_236);
    
    un98_reg_ads_0_a3_0_a2_1 : OR2
      port map(A => N_672, B => N_666, Y => un98_reg_ads_1);
    
    \VDBi_16_1_a2_1[5]\ : NAND2
      port map(A => N_2512, B => \REG[5]\, Y => N_2474);
    
    \VDBi_53_0_iv_3[13]\ : AO21TTF
      port map(A => \REGMAP_0[16]_net_1\, B => \REG[134]\, C => 
        \VDBi_53_0_iv_2[13]_net_1\, Y => \VDBi_53_0_iv_3_i[13]\);
    
    \LB_i_6[7]\ : MUX2H
      port map(A => N_2177, B => N_2189, S => LB_i_6_sn_N_2, Y
         => N_2223);
    
    \VDBi_60[24]\ : MUX2H
      port map(A => \VDBi_55[24]_net_1\, B => LBSP_in_24, S => 
        \REGMAP_0[28]_net_1\, Y => \VDBi_60[24]_net_1\);
    
    VAS_61 : MUX2H
      port map(A => \VAS[10]_net_1\, B => VAD_in_9, S => 
        \TST_c_0[1]\, Y => \VAS_61\);
    
    \VDBi_71_d[6]\ : MUX2H
      port map(A => \VDBi_66_d[6]_net_1\, B => \REG[415]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71_d[6]_net_1\);
    
    \REG_88_0[81]\ : MUX2H
      port map(A => VDB_in_0(0), B => \REG[81]\, S => N_20, Y => 
        N_2152);
    
    \VDBi_92_0_iv_0_0_2[21]\ : AO21TTF
      port map(A => N_792, B => LBSP_in_21, C => 
        \VDBi_92_0_iv_0_0_0[21]_net_1\, Y => 
        \VDBi_92_0_iv_0_0_2_i[21]\);
    
    \VDBm[14]\ : MUX2H
      port map(A => N_2310, B => \VDBi[14]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_14);
    
    REG_1_487_e : NOR3FFT
      port map(A => \REGMAP[9]_net_1\, B => \STATE1_0[8]_net_1\, 
        C => un1_STATE1_15, Y => N_3236_i);
    
    REG_1_490 : MUX2H
      port map(A => \REG_88[83]_net_1\, B => \REG[83]\, S => 
        un1_STATE1_15, Y => \REG_1_490\);
    
    N_2522_i_i_o2 : AND3
      port map(A => N_425, B => \STATE1[9]_net_1\, C => 
        \REGMAP[0]_net_1\, Y => N_457_i_0);
    
    \REG_1[179]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_219\, CLR => 
        \un10_hwres_11\, Q => \REG[179]\);
    
    \REG_1[361]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_326\, CLR => 
        \un10_hwres_17\, Q => \REG[361]\);
    
    \PIPEA[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_616\, CLR => CLEAR_25, 
        Q => \PIPEA[27]_net_1\);
    
    \PIPEA1[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_566\, CLR => CLEAR_20, 
        Q => \PIPEA1[10]_net_1\);
    
    REG_1_395 : MUX2H
      port map(A => VDB_in(21), B => \REG[430]\, S => N_3072_i_0, 
        Y => \REG_1_395\);
    
    \PIPEB_4_i[13]\ : AND2
      port map(A => DPR(13), B => N_616_1, Y => N_2627);
    
    \LB_s[3]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_82\, CLR => HWRES_c_19, 
        Q => \LB_s[3]_net_1\);
    
    un1_TCNT_1_I_33 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[5]\, B => 
        \DWACT_ADD_CI_0_g_array_12_1_0[0]\, Y => I_33_1);
    
    \RAMDTS[4]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(4), CLR => HWRES_c_21, 
        Q => \RAMDTS[4]_net_1\);
    
    LB_DOUT_164 : MUX2H
      port map(A => VDB_in(16), B => \LB_DOUT[16]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_164\);
    
    \VDBi_60[10]\ : MUX2H
      port map(A => \VDBi_58[10]_net_1\, B => LOS_c_c, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60[10]_net_1\);
    
    \PIPEA_7_i_m2[7]\ : MUX2H
      port map(A => DPR(7), B => \PIPEA1[7]_net_1\, S => N_1996_2, 
        Y => N_516);
    
    \VDBm[24]\ : MUX2H
      port map(A => N_2320, B => \VDBi[24]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_24);
    
    \LB_i[6]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_518\, CLR => 
        HWRES_c_16, Q => \LB_i[6]_net_1\);
    
    \VADm[2]\ : NOR2FT
      port map(A => \PIPEA[2]_net_1\, B => N_2507_0, Y => VADm(2));
    
    LB_DOUT_151 : MUX2H
      port map(A => VDB_in(3), B => \LB_DOUT[3]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_151\);
    
    \VDBi_71[23]\ : MUX2H
      port map(A => \VDBi_60[23]_net_1\, B => \REG[432]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[23]_net_1\);
    
    \REG_1[490]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_431\, SET => 
        \un10_hwres_26\, Q => \REG[490]\);
    
    \VDBi_92_0_iv_0_1[25]\ : AO21TTF
      port map(A => N_457_i_0_0, B => \PIPEA[25]_net_1\, C => 
        N_608, Y => \VDBi_92_0_iv_0_1_i[25]\);
    
    LB_i_523 : MUX2H
      port map(A => \LB_i[11]_net_1\, B => \LB_i_6[11]_net_1\, S
         => N_2570_1, Y => \LB_i_523\);
    
    REG_1_219 : MUX2H
      port map(A => VDB_in(10), B => \REG[179]\, S => N_2720_i_0, 
        Y => \REG_1_219\);
    
    \LB_i_6_0[3]\ : MUX2H
      port map(A => OR_RADDR(1), B => \LB_ADDR[3]_net_1\, S => 
        \STATE5[0]_net_1\, Y => N_2173);
    
    \WDOG[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \WDOG_3[4]\, CLR => 
        un15_hwres_i, Q => \WDOG_i_0_i[4]\);
    
    LB_DOUT_163 : MUX2H
      port map(A => VDB_in(15), B => \LB_DOUT[15]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_163\);
    
    \VDBi_16_r[4]\ : OA21TTF
      port map(A => \VDBi_16_1_0_i[4]\, B => N_2470_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[4]\);
    
    REG_1_486_e : OR2FT
      port map(A => N_2409, B => un1_STATE1_15, Y => N_3234_i);
    
    \REG_1[395]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_360\, CLR => 
        \un10_hwres_20\, Q => \REG[395]\);
    
    FWIMG2LOAD_111 : MUX2H
      port map(A => FWIMG2LOAD_net_1, B => VDB_in(0), S => 
        FWIMG2LOAD_0_sqmuxa, Y => \FWIMG2LOAD_111\);
    
    \REG_1[288]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_301\, CLR => 
        \un10_hwres_16\, Q => \REG[288]\);
    
    REG_1_454_e : OR2FT
      port map(A => \REGMAP_0[13]_net_1\, B => PULSE_0_sqmuxa_1, 
        Y => N_3170_i);
    
    PIPEA_589 : MUX2H
      port map(A => \PIPEA_7[0]\, B => \PIPEA[0]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_589\);
    
    REG1_1_sqmuxa : AND2
      port map(A => REG1_0_sqmuxa_1, B => NLBCLR_c, Y => 
        \REG1_1_sqmuxa\);
    
    \LB_i_6_0[9]\ : AND2
      port map(A => \LB_ADDR[9]_net_1\, B => \STATE5_3[0]_net_1\, 
        Y => N_2179);
    
    VDBi_80_m_0_m4_0_a2_1 : OR3
      port map(A => \REGMAP[32]_net_1\, B => \REGMAP[35]_net_1\, 
        C => \REGMAP_0[31]_net_1\, Y => VDBi_80_m_0_m4_0_a2_1_i);
    
    LB_i_538 : MUX2H
      port map(A => \LB_i[26]_net_1\, B => \LB_i_6[26]\, S => 
        N_2570_0, Y => \LB_i_538\);
    
    \LB_s[1]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_80\, CLR => HWRES_c_18, 
        Q => \LB_s[1]_net_1\);
    
    un1_STATE5_10_i_a2 : OR2
      port map(A => N_2573, B => \STATE5[2]_net_1\, Y => N_2603);
    
    \REG3[514]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_514_180\, CLR => 
        \un10_hwres_6_0\, Q => \RUN_c\);
    
    REG_1_403 : MUX2H
      port map(A => VDB_in(29), B => \REG[438]\, S => N_3072_i_0, 
        Y => \REG_1_403\);
    
    \VDBi_53_0_iv[0]\ : AO21TTF
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[0]_net_1\, C
         => \VDBi_53_0_iv_6[0]_net_1\, Y => \VDBi_53[0]\);
    
    \VDBi_23_m[9]\ : AND2
      port map(A => \VDBi_9_sqmuxa_0\, B => \VDBi_23[9]_net_1\, Y
         => \VDBi_23_m_i[9]\);
    
    \VDBi_16_r[7]\ : OA21TTF
      port map(A => \VDBi_16_1_0_i[7]\, B => N_2479_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[7]\);
    
    LB_i_534 : MUX2H
      port map(A => \LB_i[22]_net_1\, B => \LB_i_6[22]\, S => 
        N_2570_0, Y => \LB_i_534\);
    
    \LB_ADDR[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_553\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[10]_net_1\);
    
    \PIPEA1[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_581\, CLR => CLEAR_22, 
        Q => \PIPEA1[25]_net_1\);
    
    \LB_i_6_1[19]\ : MUX2H
      port map(A => VDB_in(19), B => \LB_DOUT[19]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2201);
    
    LB_i_540 : MUX2H
      port map(A => \LB_i[28]_net_1\, B => \LB_i_6[28]\, S => 
        N_2570_0, Y => \LB_i_540\);
    
    \PIPEA_7_i_m2[28]\ : MUX2H
      port map(A => DPR(28), B => \PIPEA1[28]_net_1\, S => 
        N_1996_0, Y => N_537);
    
    \REG_1[445]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_410\, CLR => 
        \un10_hwres_24\, Q => \REG[445]\);
    
    \LB_s[27]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_106\, CLR => 
        HWRES_c_18, Q => \LB_s[27]_net_1\);
    
    \LB_i_6_r[6]\ : AND2
      port map(A => N_2222, B => N_2572_3, Y => \LB_i_6[6]_net_1\);
    
    REG_1_444 : MUX2H
      port map(A => VDB_in(21), B => \REG[503]\, S => N_3170_i_0, 
        Y => \REG_1_444\);
    
    \VDBi_92_iv_0[0]\ : AOI21TTF
      port map(A => \RAMDTS[0]_net_1\, B => \STATE1[1]_net_1\, C
         => \FBOUT_m[0]_net_1\, Y => \VDBi_92_iv_0[0]_net_1\);
    
    \REG_1_0[125]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_133\, CLR => 
        \un10_hwres_7_0\, Q => \REG_0[125]\);
    
    \VDBi_92_0_iv_0_0[31]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[31]_net_1\, C
         => N_610, Y => \VDBi_92_0_iv_0_0[31]_net_1\);
    
    \REG_1[235]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_248\, SET => 
        \un10_hwres_13\, Q => \REG[235]\);
    
    PIPEB_33 : MUX2H
      port map(A => \PIPEB[13]_net_1\, B => N_2627, S => N_1996_4, 
        Y => \PIPEB_33\);
    
    VAS_57 : MUX2H
      port map(A => \VAS[6]_net_1\, B => VAD_in_5, S => 
        \TST_c[1]\, Y => \VAS_57\);
    
    PIPEA1_575 : MUX2H
      port map(A => N_278, B => \PIPEA1[19]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_575\);
    
    \PIPEA1_9_0[28]\ : OR2FT
      port map(A => N_85_0, B => DPR(28), Y => \PIPEA1_9[28]\);
    
    REG_1_141 : MUX2H
      port map(A => \REG[133]\, B => VDB_in(12), S => 
        REG_0_sqmuxa_0, Y => \REG_1_141\);
    
    un29_reg_ads_0_a2_0_a2_1 : NOR2FT
      port map(A => \LWORDS\, B => N_659, Y => N_660);
    
    \VDBi_18[8]\ : MUX2H
      port map(A => \VDBi_16[8]\, B => \REG[56]\, S => \TST_c[5]\, 
        Y => \VDBi_18[8]_net_1\);
    
    REG_1_223 : MUX2H
      port map(A => VDB_in(14), B => \REG[183]\, S => N_2720_i_0, 
        Y => \REG_1_223\);
    
    \VDBi[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_637\, CLR => 
        \un10_hwres_34\, Q => \VDBi[16]_net_1\);
    
    N_1897_0 : OA21
      port map(A => \STATE1_0[8]_net_1\, B => \WRITES_1\, C => 
        \REGMAP[10]_net_1\, Y => \N_1897_0\);
    
    WDOGRES : DFFC
      port map(CLK => CLK_c_c, D => \WDOGRES_71\, CLR => 
        \un10_hwres\, Q => \WDOGRES\);
    
    REG_1_387 : MUX2H
      port map(A => VDB_in_0(13), B => \REG[422]\, S => 
        N_3072_i_1, Y => \REG_1_387\);
    
    \VDBi_55[27]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[27]_net_1\, Y => \VDBi_55[27]_net_1\);
    
    un1_STATE1_32_0_2 : NOR3FTT
      port map(A => \un1_STATE1_32_0_1\, B => \STATE1[10]_net_1\, 
        C => N_479, Y => \un1_STATE1_32_0_2\);
    
    REG_1_481 : MUX2H
      port map(A => VDB_in(26), B => \REG[74]\, S => N_3234_i_0, 
        Y => \REG_1_481\);
    
    \REG_i[506]\ : INV
      port map(A => \REG[506]\, Y => \REG_i[506]_net_1\);
    
    REG_1_309 : MUX2H
      port map(A => VDB_in(31), B => \REG[296]\, S => N_2880_i_0, 
        Y => \REG_1_309\);
    
    \REG3[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_126\, CLR => 
        \un10_hwres_6\, Q => \REG[13]\);
    
    LB_s_105 : MUX2H
      port map(A => LB_in(26), B => \LB_s[26]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_105\);
    
    \REG_1[449]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_414\, CLR => 
        \un10_hwres_24\, Q => \REG[449]\);
    
    \REG_i[396]\ : INV
      port map(A => \REG[396]\, Y => REG_i_0_391);
    
    \PIPEA1_9_i[24]\ : AND2
      port map(A => DPR(24), B => N_85_3, Y => N_288);
    
    LB_DOUT_158 : MUX2H
      port map(A => VDB_in(10), B => \LB_DOUT[10]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_158\);
    
    REG_1_269 : MUX2H
      port map(A => VDB_in(7), B => \REG[256]\, S => N_2816_i_0, 
        Y => \REG_1_269\);
    
    \PIPEA_7_r[22]\ : AND2
      port map(A => N_85_1, B => N_531, Y => \PIPEA_7[22]\);
    
    REG_1_227 : MUX2H
      port map(A => VDB_in(2), B => \REG[187]\, S => N_2752_i, Y
         => \REG_1_227\);
    
    \REG_1[452]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_417\, CLR => 
        \un10_hwres_25\, Q => \REG[452]\);
    
    \VADm[27]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[27]_net_1\, Y => 
        VADm(27));
    
    REG_1_331 : MUX2H
      port map(A => VDB_in(21), B => \REG[366]\, S => N_2944_i, Y
         => \REG_1_331\);
    
    PIPEB_36 : MUX2H
      port map(A => \PIPEB[16]_net_1\, B => N_186, S => N_1996_4, 
        Y => \PIPEB_36\);
    
    \VDBm_0[19]\ : MUX2H
      port map(A => \PIPEB[19]_net_1\, B => \PIPEA[19]_net_1\, S
         => \BLTCYC_1\, Y => N_2315);
    
    un105_reg_ads_0_a3_0_a2_1 : OR2FT
      port map(A => \VAS[4]_net_1\, B => \VAS[3]_net_1\, Y => 
        N_667);
    
    \VDBi_92_0_iv_0_2[25]\ : AO21TTF
      port map(A => N_792, B => LBSP_in_25, C => 
        \VDBi_92_0_iv_0_0[25]_net_1\, Y => 
        \VDBi_92_0_iv_0_2_i[25]\);
    
    un87_reg_ads_0_a3_0_a2_1 : OR2FT
      port map(A => \VAS[1]_net_1\, B => \VAS[4]_net_1\, Y => 
        N_678);
    
    REG_1_353 : MUX2H
      port map(A => VDB_in_0(11), B => \REG[388]\, S => 
        N_2976_i_0, Y => \REG_1_353\);
    
    \VDBm_0[23]\ : MUX2H
      port map(A => \PIPEB[23]_net_1\, B => \PIPEA[23]_net_1\, S
         => \BLTCYC_1\, Y => N_2319);
    
    \VDBi_71[26]\ : MUX2H
      port map(A => \VDBi_60[26]_net_1\, B => \REG[435]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[26]_net_1\);
    
    \REG_88_0[87]\ : MUX2H
      port map(A => VDB_in_0(6), B => \REG[87]\, S => N_20, Y => 
        N_2158);
    
    VAS_53 : MUX2H
      port map(A => \VAS[2]_net_1\, B => VAD_in_1, S => 
        \TST_c[1]\, Y => \VAS_53\);
    
    REG_1_373 : MUX2H
      port map(A => VDB_in_0(15), B => \REG[408]\, S => 
        N_3008_i_0, Y => \REG_1_373\);
    
    LB_ADDR_546 : MUX2H
      port map(A => \LB_ADDR[3]_net_1\, B => \VAS[3]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_546\);
    
    un1_STATE1_34_0_a2_1_1 : OR3
      port map(A => \STATE1_0[7]_net_1\, B => \STATE1_0[1]_net_1\, 
        C => \STATE1[9]_net_1\, Y => un1_STATE1_34_0_a2_1_1_i);
    
    \REG3[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_114\, CLR => 
        \un10_hwres_6\, Q => \REG[1]\);
    
    \VDBi_92_iv_1[4]\ : AOI21TTF
      port map(A => N_457_i_0, B => \PIPEA[4]_net_1\, C => 
        \VDBi_92_iv_0[4]_net_1\, Y => \VDBi_92_iv_1[4]_net_1\);
    
    \VADm[25]\ : NOR2FT
      port map(A => \PIPEA[25]_net_1\, B => N_2507_0, Y => 
        VADm(25));
    
    \REG_1[426]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_391\, CLR => 
        \un10_hwres_22\, Q => \REG[426]\);
    
    un11_asbs_i_a2 : NOR2
      port map(A => N_230, B => \TST_c[0]\, Y => N_2423);
    
    \VDBi_16_1_a2[13]\ : AND2
      port map(A => N_2511_0, B => REG_44, Y => N_2492_i);
    
    \VDBm_0[24]\ : MUX2H
      port map(A => \PIPEB[24]_net_1\, B => \PIPEA[24]_net_1\, S
         => \BLTCYC_1\, Y => N_2320);
    
    PIPEA1_571 : MUX2H
      port map(A => N_270, B => \PIPEA1[15]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_571\);
    
    \VADm[19]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[19]_net_1\, Y => 
        VADm(19));
    
    un10_hwres_19 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_1, Y => 
        \un10_hwres_19\);
    
    \PIPEA[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_603\, CLR => CLEAR_23, 
        Q => \PIPEA[14]_net_1\);
    
    un61_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_683_i, B => N_689_i, Y => 
        \un61_reg_ads_0_a3_0_a2\);
    
    REG3_116 : MUX2H
      port map(A => \REG[3]\, B => VDB_in(3), S => REG1_0_sqmuxa, 
        Y => \REG3_116\);
    
    \VDBi_53_0_iv_5[14]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[14]\, B => 
        \VDBi_53_0_iv_0_i[14]\, C => \VDBi_53_0_iv_1_i[14]\, Y
         => \VDBi_53_0_iv_5_i[14]\);
    
    un70_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_684_i, B => N_791, Y => 
        \un70_reg_ads_0_a3_0_a2\);
    
    \VDBi_58[3]\ : MUX2H
      port map(A => \VDBi_55[3]_net_1\, B => L2A_c_c, S => 
        \REGMAP[27]_net_1\, Y => \VDBi_58[3]_net_1\);
    
    \VDBi_53_0_iv_3[14]\ : AO21TTF
      port map(A => \REGMAP_0[16]_net_1\, B => \REG[135]\, C => 
        \VDBi_53_0_iv_2[14]_net_1\, Y => \VDBi_53_0_iv_3_i[14]\);
    
    \VDBi_16_1_a3_2_0[0]\ : NOR2FT
      port map(A => \REG_c[0]\, B => \REGMAP[14]_net_1\, Y => 
        \VDBi_16_1_a3_2_0[0]_net_1\);
    
    \REG3[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_113\, CLR => 
        \un10_hwres_5\, Q => \REG_c[0]\);
    
    REG_1_208 : MUX2H
      port map(A => VDB_in(15), B => \REG[168]\, S => N_2688_i_0, 
        Y => \REG_1_208\);
    
    \VADm[13]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[13]_net_1\, Y => VADm(13));
    
    \REG_i[504]\ : INV
      port map(A => \REG[504]\, Y => \REG_i[504]_net_1\);
    
    \REG_1[171]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_211\, CLR => 
        \un10_hwres_10\, Q => \REG[171]\);
    
    \VDBi_18_i_m2[6]\ : MUX2H
      port map(A => \VDBi_16[6]\, B => \REG[54]\, S => \TST_c[5]\, 
        Y => N_491);
    
    \VAS[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_65\, CLR => HWRES_c_22, 
        Q => \VAS[14]_net_1\);
    
    un1_STATE2_16_0_0 : NAND3FTT
      port map(A => un1_STATE2_16_0_0_0_i, B => N_79, C => N_580, 
        Y => un1_STATE2_16);
    
    \REG_1_m[199]\ : NAND2
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[199]\, Y => 
        \REG_1_m[199]_net_1\);
    
    \PIPEB_4_i[6]\ : AND2
      port map(A => DPR(6), B => N_616, Y => N_2620);
    
    \REG_1[155]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_195\, CLR => 
        \un10_hwres_9\, Q => \REG[155]\);
    
    \LB_i_6_1[10]\ : MUX2H
      port map(A => VDB_in_0(10), B => \LB_DOUT[10]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2192);
    
    DSSF1_2_0 : OR2FT
      port map(A => N_230, B => \TST_c_0[0]\, Y => DSSF1_2);
    
    \PIPEB_4_i[0]\ : AND2
      port map(A => DPR(0), B => N_616, Y => N_2614);
    
    un1_STATE1_28_i_0 : OA21FTF
      port map(A => \STATE1[10]_net_1\, B => N_231, C => N_2428_i, 
        Y => \un1_STATE1_28_i_0\);
    
    \REG_i[509]\ : INV
      port map(A => \REG[509]\, Y => \REG_i[509]_net_1\);
    
    \VDBi_58[9]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[9]\, B => \VDBi_23_m_i[9]\, 
        C => \VDBi_58_0[9]\, Y => \VDBi_58[9]_net_1\);
    
    un1_TCNT_1_I_35 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_0[0]\, B => 
        \DWACT_ADD_CI_0_TMP_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\);
    
    un117_reg_ads_0_a3_0_a2_0 : OR2FT
      port map(A => \VAS[2]_net_1\, B => \VAS[5]_net_1\, Y => 
        N_666);
    
    \PIPEA[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_593\, CLR => CLEAR_25, 
        Q => \PIPEA[4]_net_1\);
    
    \PIPEA1[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_575\, CLR => CLEAR_21, 
        Q => \PIPEA1[19]_net_1\);
    
    REG_1_216 : MUX2H
      port map(A => VDB_in(7), B => \REG[176]\, S => N_2720_i, Y
         => \REG_1_216\);
    
    \REG_1[48]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_455\, CLR => 
        \un10_hwres_26\, Q => \REG[48]\);
    
    \VAS[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_56\, CLR => HWRES_c_22_0, 
        Q => \VAS[5]_net_1\);
    
    PULSE_0_sqmuxa_1_0_a2_0_i2_0_a2_0_a2_0 : OR2FT
      port map(A => \STATE1_0[8]_net_1\, B => \WRITES_0\, Y => 
        PULSE_0_sqmuxa_1_0);
    
    LB_s_85 : MUX2H
      port map(A => LB_in(6), B => \LB_s[6]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_85\);
    
    DSSF1_2_0_a2 : NAND2
      port map(A => DS0B_c, B => DS1B_c, Y => N_230);
    
    \STATE1_1[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[8]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1_1[2]_net_1\);
    
    \PIPEA_7_i_m2[20]\ : MUX2H
      port map(A => DPR(20), B => \PIPEA1[20]_net_1\, S => 
        N_1996_1, Y => N_529);
    
    un776_regmap_9 : OR3FTT
      port map(A => \un776_regmap_4\, B => \REGMAP[1]_net_1\, C
         => \REGMAP[6]_net_1\, Y => un776_regmap_9_i);
    
    ASBS : DFFS
      port map(CLK => CLK_c_c, D => \ASBSF1\, SET => HWRES_c_13, 
        Q => \TST_c[0]\);
    
    \VDBi_71[6]\ : MUX2H
      port map(A => \VDBi_58[6]_net_1\, B => \VDBi_71_d[6]_net_1\, 
        S => \VDBi_71_s[1]_net_1\, Y => \VDBi_71[6]_net_1\);
    
    un1_STATE5_15_i_a2_1 : NOR2
      port map(A => N_65, B => N_66, Y => N_2606_i_i);
    
    un10_hwres_7 : OR2
      port map(A => HWRES_c_0_6, B => WDOGTO_2, Y => 
        \un10_hwres_7\);
    
    \REG_1[363]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_328\, CLR => 
        \un10_hwres_17\, Q => \REG[363]\);
    
    \PIPEA1[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_582\, CLR => CLEAR_22, 
        Q => \PIPEA1[26]_net_1\);
    
    LB_ADDR_0_sqmuxa_1 : NOR2FT
      port map(A => \STATE1_0[9]_net_1\, B => N_2535, Y => 
        \LB_ADDR_0_sqmuxa_1\);
    
    \VDBi_53_0_iv_0[4]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_140, C => 
        \REG_1_m[253]_net_1\, Y => \VDBi_53_0_iv_0_i[4]\);
    
    \VDBi_53_0_iv_6[8]\ : OR3
      port map(A => \VDBi_53_0_iv_5_i[8]\, B => 
        \VDBi_53_0_iv_2_i[8]\, C => \VDBi_53_0_iv_0_i[8]\, Y => 
        \VDBi_53_0_iv_6_i[8]\);
    
    \VDBi_66_d[1]\ : MUX2H
      port map(A => LBSP_in_1, B => N_2018, S => N_2033, Y => 
        \VDBi_66_d[1]_net_1\);
    
    VAS_64 : MUX2H
      port map(A => \VAS[13]_net_1\, B => VAD_in_12, S => 
        \TST_c_0[1]\, Y => \VAS_64\);
    
    \OR_RDATA_5_i[8]\ : AND2
      port map(A => N_2572, B => LB_in(8), Y => N_31);
    
    \VDBi_71_i_m2[7]\ : MUX2H
      port map(A => \VDBi_60[7]_net_1\, B => 
        \VDBi_71_i_m2_d[7]_net_1\, S => \VDBi_71_s[4]_net_1\, Y
         => N_492);
    
    \LB_DOUT[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_159\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[11]_net_1\);
    
    \RAMDTS[0]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(0), CLR => HWRES_c_20, 
        Q => \RAMDTS[0]_net_1\);
    
    \REG_i[266]\ : INV
      port map(A => \REG[266]\, Y => REG_i_0_261);
    
    \VDBi_16_1_a2_0[2]\ : AND2
      port map(A => N_2511, B => REG_33, Y => N_2464_i);
    
    un1_STATE5_15_i_a2 : NOR2
      port map(A => \STATE5_0[0]_net_1\, B => \STATE5_0[2]_net_1\, 
        Y => N_2601_i);
    
    \VADm[30]\ : NOR2FT
      port map(A => \PIPEA[30]_net_1\, B => N_2507_1, Y => 
        VADm(30));
    
    \VDBi_18[22]\ : NAND2
      port map(A => \REG[70]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[22]_net_1\);
    
    \VDBi_53_0_iv_5[10]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[10]\, B => 
        \VDBi_53_0_iv_0_i[10]\, C => \VDBi_53_0_iv_1_i[10]\, Y
         => \VDBi_53_0_iv_5_i[10]\);
    
    \PIPEB[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_44\, CLR => CLEAR_27, 
        Q => \PIPEB[24]_net_1\);
    
    \PIPEA1_9_i[8]\ : AND2
      port map(A => DPR(8), B => N_85, Y => N_256);
    
    \REG_1[486]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_427\, SET => 
        \un10_hwres_25\, Q => \REG[486]\);
    
    REG_1_294 : MUX2H
      port map(A => VDB_in(16), B => \REG[281]\, S => N_2880_i, Y
         => \REG_1_294\);
    
    \VDBi_53_0_iv_1[2]\ : AO21TTF
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[235]\, C => 
        \REG_1_m[187]_net_1\, Y => \VDBi_53_0_iv_1_i[2]\);
    
    \STATE5_ns_0_0_a2_1[0]\ : NOR2FT
      port map(A => \STATE5_0[0]_net_1\, B => \STATE5[1]_net_1\, 
        Y => N_2599_1);
    
    \REG_1[122]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_130\, CLR => 
        \un10_hwres_7_0\, Q => \REG[122]\);
    
    \VDBi_53_0_iv_3[10]\ : AO21TTF
      port map(A => \REGMAP_0[16]_net_1\, B => \REG[131]\, C => 
        \VDBi_53_0_iv_2[10]_net_1\, Y => \VDBi_53_0_iv_3_i[10]\);
    
    \TCNT[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[6]\, CLR => 
        \un10_hwres_33\, Q => \TCNT_i_i[6]\);
    
    LB_i_513 : MUX2H
      port map(A => \LB_i[1]_net_1\, B => \LB_i_6[1]_net_1\, S
         => N_2570, Y => \LB_i_513\);
    
    \VDBi_55[24]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[24]_net_1\, Y => \VDBi_55[24]_net_1\);
    
    un74_reg_ads_0_a3 : AND3FTT
      port map(A => N_198, B => \un74_reg_ads_0_a3_1\, C => N_463, 
        Y => \un74_reg_ads_0_a3\);
    
    REG_1_428 : MUX2H
      port map(A => VDB_in_0(5), B => \REG[487]\, S => N_3170_i, 
        Y => \REG_1_428\);
    
    OR_RDATA_190 : MUX2H
      port map(A => N_31, B => \OR_RDATA[8]_net_1\, S => N_1832, 
        Y => \OR_RDATA_190\);
    
    un1_STATE5_14_i_0_a2 : NAND2
      port map(A => N_65, B => \STATE5[2]_net_1\, Y => N_2592);
    
    \VDBi_92_0_iv_1[20]\ : AOI21TTF
      port map(A => \LB_s[20]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[20]_net_1\, Y => 
        \VDBi_92_0_iv_1[20]_net_1\);
    
    \VDBi_71[22]\ : MUX2H
      port map(A => \VDBi_60[22]_net_1\, B => \REG[431]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[22]_net_1\);
    
    \REG_1[124]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_132\, CLR => 
        \un10_hwres_7_0\, Q => REG_123);
    
    REG_1_357 : MUX2H
      port map(A => VDB_in_0(15), B => \REG[392]\, S => 
        N_2976_i_0, Y => \REG_1_357\);
    
    REG_1_377 : MUX2H
      port map(A => VDB_in_0(3), B => \REG[412]\, S => N_3072_i, 
        Y => \REG_1_377\);
    
    \PIPEA_7_s[29]\ : OR2FT
      port map(A => N_85_0, B => N_538, Y => \PIPEA_7[29]\);
    
    un117_reg_ads_0_a3_0_a2_2 : OR2FT
      port map(A => \VAS[1]_net_1\, B => N_667, Y => N_684_i);
    
    REG_1_451 : MUX2H
      port map(A => VDB_in(28), B => \REG[510]\, S => N_3170_i_0, 
        Y => \REG_1_451\);
    
    un1_STATE2_13_i_0_a2_1 : NAND2FT
      port map(A => \STATE2[1]_net_1\, B => N_472_i_0, Y => N_676);
    
    \TCNT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[4]\, CLR => 
        \un10_hwres_33\, Q => \TCNT_i_i[4]\);
    
    \VDBi_60[27]\ : MUX2H
      port map(A => \VDBi_55[27]_net_1\, B => LBSP_in_27, S => 
        \REGMAP_0[28]_net_1\, Y => \VDBi_60[27]_net_1\);
    
    REG_1_326 : MUX2H
      port map(A => VDB_in(16), B => \REG[361]\, S => N_2944_i, Y
         => \REG_1_326\);
    
    \VDBi_60[4]\ : MUX2H
      port map(A => \VDBi_58[4]_net_1\, B => L0_c_c, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60[4]_net_1\);
    
    \VDBi_23[29]\ : MUX2H
      port map(A => \VDBi_18[29]_net_1\, B => \REG_i[511]_net_1\, 
        S => \REGMAP_0[13]_net_1\, Y => \VDBi_23[29]_net_1\);
    
    \STATE1_ns_0_iv_0_a2_0_2[9]\ : OR3FTT
      port map(A => \REGMAP[15]_net_1\, B => N_486, C => N_1898, 
        Y => \STATE1_ns_0_iv_0_a2_0_1[9]_net_1\);
    
    REG_1_471 : MUX2H
      port map(A => VDB_in(16), B => \REG[64]\, S => N_3234_i_1, 
        Y => \REG_1_471\);
    
    \REG_1[126]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_134\, CLR => 
        \un10_hwres_8\, Q => REG_125);
    
    VDBi_631 : MUX2H
      port map(A => \VDBi_92[10]\, B => \VDBi[10]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_631\);
    
    un10_hwres_35 : OR2
      port map(A => HWRES_c_0_3, B => WDOGTO_0, Y => 
        \un10_hwres_35\);
    
    \VDBi_71[17]\ : MUX2H
      port map(A => \VDBi_60[17]_net_1\, B => \REG[426]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[17]_net_1\);
    
    \REGMAP_1[13]\ : DFF
      port map(CLK => CLK_c_c, D => \un84_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_1[13]_net_1\);
    
    REG_1_266 : MUX2H
      port map(A => VDB_in(4), B => \REG[253]\, S => N_2816_i_0, 
        Y => \REG_1_266\);
    
    \REG_1[294]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_307\, CLR => 
        \un10_hwres_16\, Q => \REG[294]\);
    
    \PIPEA_7_i_m2[26]\ : MUX2H
      port map(A => DPR(26), B => \PIPEA1[26]_net_1\, S => 
        N_1996_0, Y => N_535);
    
    \REG_1_0[126]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_134\, CLR => 
        \un10_hwres_8_0\, Q => \REG_0[126]\);
    
    \REG_1[292]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_305\, CLR => 
        \un10_hwres_16\, Q => \REG[292]\);
    
    REG_1_220 : MUX2H
      port map(A => VDB_in(11), B => \REG[180]\, S => N_2720_i_0, 
        Y => \REG_1_220\);
    
    \PIPEA1[30]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEA1_586\, SET => CLEAR_22, 
        Q => \PIPEA1[30]_net_1\);
    
    un1_TCNT_1_I_7 : AND2
      port map(A => \TCNT_i_i[4]\, B => N_83, Y => 
        \DWACT_ADD_CI_0_g_array_0_4[0]\);
    
    TCNT_0_sqmuxa_i_s : OR3FFT
      port map(A => \REGMAP[15]_net_1\, B => \WRITES_1\, C => 
        N_1898, Y => \TCNT_0_sqmuxa_i_s\);
    
    un29_reg_ads_0_a2_0_a2 : NOR2
      port map(A => N_683_i, B => un33_reg_ads_1, Y => 
        \un29_reg_ads_0_a2_0_a2\);
    
    \REG_i[294]\ : INV
      port map(A => \REG[294]\, Y => REG_i_0_289);
    
    VDBi_9_sqmuxa_0 : AND3
      port map(A => \un776_regmap_23\, B => \VDBi_9_sqmuxa_1\, C
         => \VDBi_9_sqmuxa_i_1\, Y => \VDBi_9_sqmuxa_0\);
    
    \VDBi_16_s[2]\ : OR3
      port map(A => N_2464_i, B => \VDBi_16_1_0_i[2]\, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[2]\);
    
    \VDBi_16_1_a2_0[7]\ : AND2
      port map(A => N_2511, B => REG_38, Y => N_2479_i);
    
    un78_reg_ads_0_a3_0_a2_0 : OR2
      port map(A => N_198, B => \VAS[2]_net_1\, Y => N_689_i);
    
    \VDBi_92_0_iv_0_a2_2[10]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[10]_net_1\, Y => 
        N_624);
    
    \REG_1_m[194]\ : NAND2
      port map(A => \REGMAP_0[20]_net_1\, B => \REG[194]\, Y => 
        \REG_1_m[194]_net_1\);
    
    PULSE_0_sqmuxa_1_0_a2_0_i2_0_a2_0_a2_1 : OR2FT
      port map(A => \STATE1_0[8]_net_1\, B => \WRITES_0\, Y => 
        PULSE_0_sqmuxa_1_1);
    
    \REG_1_m[254]\ : NAND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[254]\, Y => 
        \REG_1_m[254]_net_1\);
    
    LB_ACK_1_sqmuxa_i_0 : NOR3FFT
      port map(A => \STATE5_0[0]_net_1\, B => \LB_REQ_sync\, C
         => \STATE5_i_0[2]\, Y => \LB_ACK_1_sqmuxa_i_0\);
    
    un1_LBUSTMO_1_I_11 : XOR2FT
      port map(A => N_66, B => \LBUSTMO[2]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_1[0]\);
    
    \LB_i[29]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_541\, CLR => 
        HWRES_c_16, Q => \LB_i[29]_net_1\);
    
    un776_regmap_23_0 : OR2
      port map(A => \REGMAP[21]_net_1\, B => \REGMAP[22]_net_1\, 
        Y => \un776_regmap_23_0\);
    
    un94_reg_ads_0_a3_0_a2 : AND3
      port map(A => N_688, B => N_685, C => N_682, Y => 
        \un94_reg_ads_0_a3_0_a2\);
    
    \VDBi_66_s[1]\ : NOR2
      port map(A => N_2033, B => \REGMAP[28]_net_1\, Y => 
        \VDBi_66_s[1]_net_1\);
    
    un1_REG_0_sqmuxa_i_o2_i : INV
      port map(A => \STATE5[0]_net_1\, Y => \STATE5_i_0[0]\);
    
    \STATE2_ns_o2_0_0_1[0]\ : NOR3FTT
      port map(A => EVRDY_c, B => \EFS\, C => N_622, Y => 
        N_1756_1);
    
    \VDBi_92_0_iv[15]\ : OAI21FTT
      port map(A => \VDBi_77[15]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[15]_net_1\, Y => \VDBi_92[15]\);
    
    \VDBi_92_iv_1[6]\ : AOI21TTF
      port map(A => N_457_i_0, B => \PIPEA[6]_net_1\, C => 
        \VDBi_92_iv_0[6]_net_1\, Y => \VDBi_92_iv_1[6]_net_1\);
    
    \VDBi_92_0_iv_1[27]\ : AOI21TTF
      port map(A => \LB_s[27]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[27]_net_1\, Y => 
        \VDBi_92_0_iv_1[27]_net_1\);
    
    un1_TCNT_1_I_10 : AND2
      port map(A => \TCNT_i_i[6]\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_6[0]\);
    
    REG_1_414 : MUX2H
      port map(A => VDB_in_0(8), B => \REG[449]\, S => N_3104_i_0, 
        Y => \REG_1_414\);
    
    PIPEA_600 : MUX2H
      port map(A => \PIPEA_7[11]\, B => \PIPEA[11]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_600\);
    
    \REG_1[53]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_460\, CLR => 
        \un10_hwres_28\, Q => \REG[53]\);
    
    un7_ronly_0_a3_0_a2_0 : OR3
      port map(A => \un7_ronly_0_a3_0_a2_0_0\, B => 
        \VAS[9]_net_1\, C => \VAS[10]_net_1\, Y => N_658);
    
    \PIPEA_7_r[11]\ : AND2
      port map(A => N_85_2, B => N_520, Y => \PIPEA_7[11]\);
    
    \REG_1[509]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_450\, CLR => 
        \un10_hwres_27\, Q => \REG[509]\);
    
    \PIPEA_7_r[8]\ : AND2
      port map(A => N_85_2, B => N_517, Y => \PIPEA_7[8]\);
    
    \REGMAP[32]\ : DFF
      port map(CLK => CLK_c_c, D => \un117_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[32]_net_1\);
    
    REG_1_333 : MUX2H
      port map(A => VDB_in(23), B => \REG[368]\, S => N_2944_i_0, 
        Y => \REG_1_333\);
    
    \LB_i_6_r[3]\ : AND2
      port map(A => N_2219, B => N_2572_3, Y => \LB_i_6[3]_net_1\);
    
    un1_LB_DOUT_0_sqmuxa_0 : NAND3FFT
      port map(A => un1_LB_DOUT_0_sqmuxa_0_1_i, B => N_2430, C
         => LB_DOUT_0_sqmuxa_0, Y => un1_LB_DOUT_0_sqmuxa);
    
    un3_clear_i_a3 : OR2FT
      port map(A => EVRDY_c, B => CLEAR_0, Y => N_2371_i_0);
    
    LB_DOUT_162 : MUX2H
      port map(A => VDB_in(14), B => \LB_DOUT[14]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_162\);
    
    \PIPEB[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_51\, CLR => CLEAR_28, 
        Q => \PIPEB[31]_net_1\);
    
    \REG_1[65]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_472\, CLR => 
        \un10_hwres_29\, Q => \REG[65]\);
    
    \REG_1[182]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_222\, CLR => 
        \un10_hwres_11\, Q => \REG[182]\);
    
    \REG_1[367]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_332\, CLR => 
        \un10_hwres_17\, Q => \REG[367]\);
    
    \VAS[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_60\, CLR => HWRES_c_23, 
        Q => \VAS[9]_net_1\);
    
    \LB_s[5]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_84\, CLR => HWRES_c_19, 
        Q => \LB_s[5]_net_1\);
    
    \PIPEA1_9_i[26]\ : AND2
      port map(A => DPR(26), B => N_85_3, Y => N_292);
    
    VDBi_624 : MUX2H
      port map(A => \VDBi_92[3]\, B => \VDBi[3]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_624\);
    
    \LB_i_6[6]\ : MUX2H
      port map(A => N_2176, B => N_2188, S => LB_i_6_sn_N_2, Y
         => N_2222);
    
    \REG_1[184]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_224\, CLR => 
        \un10_hwres_11\, Q => \REG[184]\);
    
    \LB_i_6[1]\ : MUX2H
      port map(A => N_2171, B => N_2183, S => LB_i_6_sn_N_2, Y
         => N_2217);
    
    VDBi_629 : MUX2H
      port map(A => \VDBi_92[8]\, B => \VDBi[8]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_629\);
    
    \REG_1[450]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_415\, CLR => 
        \un10_hwres_24\, Q => \REG[450]\);
    
    LB_DOUT_171 : MUX2H
      port map(A => VDB_in(23), B => \LB_DOUT[23]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_171\);
    
    un10_hwres : OR2
      port map(A => HWRES_c_0, B => \WDOGTO\, Y => \un10_hwres\);
    
    \VDBi[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_639\, CLR => 
        \un10_hwres_34\, Q => \VDBi[18]_net_1\);
    
    \LB_i_6_r[24]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_0, C => N_2206, 
        Y => \LB_i_6[24]\);
    
    LB_ADDR_552 : MUX2H
      port map(A => \LB_ADDR[9]_net_1\, B => \VAS[9]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_552\);
    
    \VDBi_16_r[5]\ : OA21TTF
      port map(A => \VDBi_16_1_0_i[5]\, B => N_2473_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[5]\);
    
    PIPEA1_564 : MUX2H
      port map(A => N_256, B => \PIPEA1[8]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_564\);
    
    \REG_1[186]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_226\, CLR => 
        \un10_hwres_11\, Q => \REG[186]\);
    
    \LB_i[24]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_536\, CLR => 
        HWRES_c_15, Q => \LB_i[24]_net_1\);
    
    \VDBi_92_iv_0[4]\ : AOI21TTF
      port map(A => \RAMDTS[4]_net_1\, B => \STATE1[1]_net_1\, C
         => \FBOUT_m[4]_net_1\, Y => \VDBi_92_iv_0[4]_net_1\);
    
    un776_regmap_17 : NOR3FTT
      port map(A => \un776_regmap_13\, B => \REGMAP[35]_net_1\, C
         => un776_regmap_9_i, Y => \un776_regmap_17\);
    
    \REG_1[54]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_461\, CLR => 
        \un10_hwres_28\, Q => \REG[54]\);
    
    LB_s_102 : MUX2H
      port map(A => LB_in(23), B => \LB_s[23]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_102\);
    
    \VDBi_53_0_iv_5[9]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[9]\, B => 
        \VDBi_53_0_iv_0_i[9]\, C => \VDBi_53_0_iv_1_i[9]\, Y => 
        \VDBi_53_0_iv_5_i[9]\);
    
    un108_reg_ads_0_a3_0_a2_0 : OR2
      port map(A => \VAS[5]_net_1\, B => \VAS[2]_net_1\, Y => 
        N_671);
    
    \LB_i[17]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_529\, CLR => 
        HWRES_c_15, Q => \LB_i[17]_net_1\);
    
    REG_1_406 : MUX2H
      port map(A => VDB_in_0(0), B => \REG[441]\, S => N_3104_i, 
        Y => \REG_1_406\);
    
    un1_noe16wi_i_s_0_o2 : OR2
      port map(A => \MBLTCYC\, B => N_2507_1, Y => N_436);
    
    PIPEA_609 : MUX2H
      port map(A => \PIPEA_7[20]\, B => \PIPEA[20]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_609\);
    
    un5_noe16ri_0_0_a2_0_0 : NOR2FT
      port map(A => \MBLTCYC\, B => \ADACKCYC\, Y => \NOEAD_c_0\);
    
    un1_STATE5_14_i_0_o2 : AND2
      port map(A => un2_nlbrdy_i_0, B => nLBRDY_c, Y => N_65);
    
    \REG_1_m[188]\ : NAND2
      port map(A => \REGMAP[20]_net_1\, B => \REG[188]\, Y => 
        \REG_1_m[188]_net_1\);
    
    \REGMAP[27]\ : DFF
      port map(CLK => CLK_c_c, D => \un98_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[27]_net_1\);
    
    WDOG_3_I_22 : XOR2
      port map(A => \WDOG[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => \WDOG_3[2]\);
    
    \REG_1[60]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_467\, CLR => 
        \un10_hwres_29\, Q => \REG[60]\);
    
    \REG_1[82]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_489\, CLR => 
        \un10_hwres_31\, Q => \REG[82]\);
    
    \REGMAP[0]\ : DFF
      port map(CLK => CLK_c_c, D => \un2_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[0]_net_1\);
    
    REG_1_464 : MUX2H
      port map(A => VDB_in_0(9), B => \REG[57]\, S => N_3234_i, Y
         => \REG_1_464\);
    
    \VDBi_92_0_iv_1[24]\ : AOI21TTF
      port map(A => \LB_s[24]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[24]_net_1\, Y => 
        \VDBi_92_0_iv_1[24]_net_1\);
    
    REG_1_505 : MUX2H
      port map(A => \REG[98]\, B => VDB_in_0(9), S => N_2416_i, Y
         => \REG_1_505\);
    
    \LB_s[15]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_94\, CLR => HWRES_c_17, 
        Q => \LB_s[15]_net_1\);
    
    \VDBi_92_0_iv_1[30]\ : AOI21TTF
      port map(A => \LB_s[30]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[30]_net_1\, Y => 
        \VDBi_92_0_iv_1[30]_net_1\);
    
    \VDBi_53_0_iv_0[3]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_139, C => 
        \REG_1_m[252]_net_1\, Y => \VDBi_53_0_iv_0_i[3]\);
    
    \PIPEB[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_28\, CLR => CLEAR_28, 
        Q => \PIPEB[8]_net_1\);
    
    \STATE1_ns_0_iv_0[8]\ : AO21TTF
      port map(A => N_2531, B => \STATE1_0[2]_net_1\, C => N_2550, 
        Y => \STATE1_ns[8]\);
    
    \VDBi_23[4]\ : MUX2H
      port map(A => \VDBi_16[4]\, B => \VDBi_23_d[4]_net_1\, S
         => \VDBi_23_s[7]_net_1\, Y => \VDBi_23[4]_net_1\);
    
    \REGMAP[22]\ : DFF
      port map(CLK => CLK_c_c, D => \un74_reg_ads_0_a3\, Q => 
        \REGMAP[22]_net_1\);
    
    \STATE1[10]\ : DFFS
      port map(CLK => CLK_c_c, D => \STATE1_ns[0]\, SET => 
        \un10_hwres_32\, Q => \STATE1[10]_net_1\);
    
    \PIPEB[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_27\, CLR => CLEAR_28, 
        Q => \PIPEB[7]_net_1\);
    
    un10_hwres_34 : OR2
      port map(A => HWRES_c_0_3, B => WDOGTO_0, Y => 
        \un10_hwres_34\);
    
    \VDBi_92_0_iv_0_a2_2[25]\ : NAND2
      port map(A => N_793, B => \REG[507]\, Y => N_605);
    
    \PULSE_42_f0_i_o2[0]\ : AND2
      port map(A => \REGMAP_i_0_i[3]\, B => \STATE1[8]_net_1\, Y
         => N_2419);
    
    REG_1_445 : MUX2H
      port map(A => VDB_in(22), B => \REG[504]\, S => N_3170_i_0, 
        Y => \REG_1_445\);
    
    LB_DOUT_178 : MUX2H
      port map(A => VDB_in(30), B => \LB_DOUT[30]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_178\);
    
    \STATE5_ns_0_0_a2_0[0]\ : OR3FFT
      port map(A => \LB_REQ_sync\, B => N_2607, C => 
        \OR_RREQ_sync\, Y => N_2600);
    
    \VDBi_58[4]\ : MUX2H
      port map(A => \VDBi_55[4]_net_1\, B => REG_332, S => 
        \REGMAP[27]_net_1\, Y => \VDBi_58[4]_net_1\);
    
    \OR_RDATA[7]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_189\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[7]_net_1\);
    
    \LB_DOUT[30]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_178\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[30]_net_1\);
    
    \PIPEA_7_r[10]\ : AND2
      port map(A => N_85_2, B => N_519, Y => \PIPEA_7[10]\);
    
    \VDBi_23[0]\ : MUX2H
      port map(A => \VDBi_21[0]_net_1\, B => \REG[482]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23[0]_net_1\);
    
    \REG_1[163]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_203\, CLR => 
        \un10_hwres_9\, Q => \REG[163]\);
    
    \LB_s[29]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_108\, CLR => 
        HWRES_c_18, Q => \LB_s[29]_net_1\);
    
    \REG_1[72]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_479\, CLR => 
        \un10_hwres_30\, Q => \REG[72]\);
    
    \LB_i_6_1[23]\ : MUX2H
      port map(A => VDB_in(23), B => \LB_DOUT[23]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2205);
    
    \REG_1[177]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_217\, CLR => 
        \un10_hwres_10\, Q => \REG[177]\);
    
    \VDBi_55[1]\ : MUX2H
      port map(A => \VDBi_53[1]\, B => SPULSE1_c_c, S => 
        \REGMAP[26]_net_1\, Y => \VDBi_55[1]_net_1\);
    
    \REG_1[81]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_488\, CLR => 
        \un10_hwres_30\, Q => \REG[81]\);
    
    \VDBi_92_0_iv_1[13]\ : AOI21TTF
      port map(A => \LB_s[13]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[13]_net_1\, Y => 
        \VDBi_92_0_iv_1[13]_net_1\);
    
    \VDBi_92_0_iv_0_0_0[10]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[10]_net_1\, C
         => N_624, Y => \VDBi_92_0_iv_0_0_0[10]_net_1\);
    
    LB_i_531 : MUX2H
      port map(A => \LB_i[19]_net_1\, B => \LB_i_6[19]\, S => 
        N_2570_1, Y => \LB_i_531\);
    
    REG_1_427 : MUX2H
      port map(A => VDB_in_0(4), B => \REG[486]\, S => N_3170_i, 
        Y => \REG_1_427\);
    
    un10_hwres_6_0 : OR2
      port map(A => HWRES_c_0_6_0, B => WDOGTO_2, Y => 
        \un10_hwres_6_0\);
    
    REG_1_337 : MUX2H
      port map(A => VDB_in(27), B => \REG[372]\, S => N_2944_i_0, 
        Y => \REG_1_337\);
    
    \VDBm[13]\ : MUX2H
      port map(A => N_2309, B => \VDBi[13]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_13);
    
    \REGMAP[28]\ : DFF
      port map(CLK => CLK_c_c, D => \un102_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[28]_net_1\);
    
    \VDBi_92_0_iv_0[17]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[17]_net_1\, C
         => \PIPEA_m[17]_net_1\, Y => \VDBi_92_0_iv_0[17]_net_1\);
    
    \VDBi_92_0_iv_0[9]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[9]_net_1\, C
         => \PIPEA_m[9]_net_1\, Y => \VDBi_92_0_iv_0[9]_net_1\);
    
    REG_1_431 : MUX2H
      port map(A => VDB_in_0(8), B => \REG[490]\, S => N_3170_i, 
        Y => \REG_1_431\);
    
    \REGMAP[34]\ : DFF
      port map(CLK => CLK_c_c, D => \un120_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[34]_net_1\);
    
    un84_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_724, B => un84_reg_ads_1, Y => 
        \un84_reg_ads_0_a3_0_a2\);
    
    REG_1_449 : MUX2H
      port map(A => VDB_in(26), B => \REG[508]\, S => N_3170_i_0, 
        Y => \REG_1_449\);
    
    \STATE1_ns_1_iv_0_0_a2[5]\ : OA21FTT
      port map(A => N_462, B => N_480, C => \TST_c_0[2]\, Y => 
        N_572_i);
    
    \PIPEB[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_32\, CLR => CLEAR_26, 
        Q => \PIPEB[12]_net_1\);
    
    REG_1_493 : MUX2H
      port map(A => \REG_88[86]_net_1\, B => \REG[86]\, S => 
        un1_STATE1_15, Y => \REG_1_493\);
    
    VDBi_640 : MUX2H
      port map(A => \VDBi_92[19]\, B => \VDBi[19]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_640\);
    
    \VDBi_16_1_a2_0[15]\ : AND2
      port map(A => N_2512_0, B => \REG[15]\, Y => N_2497_i);
    
    PULSE_1_245 : MUX2H
      port map(A => \PULSE_42[10]\, B => \PULSE[10]\, S => 
        un1_STATE1_17, Y => \PULSE_1_245\);
    
    un1_LBUSTMO_1_I_27 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_1_0[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\);
    
    un1_STATE1_5_i_a2_i_o2 : NOR2
      port map(A => \STATE1[7]_net_1\, B => \STATE1[10]_net_1\, Y
         => N_2410);
    
    un1_STATE2_13_i_0_a2_1_0 : NOR3FFT
      port map(A => DPR(28), B => DPR(30), C => 
        \un1_STATE2_13_i_0_a2_1_0_0\, Y => N_583);
    
    \LB_DOUT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_153\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[5]_net_1\);
    
    \STATE2[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE2[0]_net_1\, CLR => 
        CLEAR, Q => \STATE2[4]_net_1\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \REG_1[245]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_258\, SET => 
        \un10_hwres_13\, Q => \REG[245]\);
    
    LB_ACK : DFFC
      port map(CLK => ALICLK_c, D => \LB_ACK_1_sqmuxa_i_0\, CLR
         => HWRES_c_14, Q => \LB_ACK\);
    
    \VDBi_16_r[14]\ : OA21TTF
      port map(A => N_2495_i, B => N_2494_i, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[14]\);
    
    un1_TCNT_1_I_17 : XOR2
      port map(A => \TCNT_i_i[4]\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_3[0]\);
    
    \VDBm[23]\ : MUX2H
      port map(A => N_2319, B => \VDBi[23]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_23);
    
    \PIPEA[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_599\, CLR => CLEAR_23, 
        Q => \PIPEA[10]_net_1\);
    
    un5_noe16ri_0_0_0 : AO21
      port map(A => N_566_1, B => N_436, C => \NOEAD_c_0_0\, Y
         => un5_noe16ri_0);
    
    REG_1_422 : MUX2H
      port map(A => \REG[481]\, B => VDB_in_0(0), S => 
        FWIMG2LOAD_0_sqmuxa, Y => \REG_1_422\);
    
    \VDBm_0[12]\ : MUX2H
      port map(A => \PIPEB[12]_net_1\, B => \PIPEA[12]_net_1\, S
         => \BLTCYC_2\, Y => N_2308);
    
    \VDBi_92_0_iv_0[20]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[20]_net_1\, C
         => \PIPEA_m[20]_net_1\, Y => \VDBi_92_0_iv_0[20]_net_1\);
    
    un10_hwres_4 : OR2
      port map(A => HWRES_c_0_6, B => \WDOGTO\, Y => 
        \un10_hwres_4\);
    
    LB_s_99 : MUX2H
      port map(A => LB_in(20), B => \LB_s[20]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_99\);
    
    \REG_1[493]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_434\, CLR => 
        \un10_hwres_26\, Q => \REG[493]\);
    
    \REG_1_m[156]\ : NAND2
      port map(A => \REGMAP[18]_net_1\, B => \REG[156]\, Y => 
        \REG_1_m[156]_net_1\);
    
    \PIPEA[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_611\, CLR => CLEAR_24, 
        Q => \PIPEA[22]_net_1\);
    
    \LB_s[13]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_92\, CLR => HWRES_c_17, 
        Q => \LB_s[13]_net_1\);
    
    \PIPEA1[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_571\, CLR => CLEAR_21, 
        Q => \PIPEA1[15]_net_1\);
    
    \VDBi_60[19]\ : MUX2H
      port map(A => \VDBi_55[19]_net_1\, B => LBSP_in_19, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[19]_net_1\);
    
    \REG_1[71]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_478\, CLR => 
        \un10_hwres_30\, Q => \REG[71]\);
    
    PIPEA_599 : MUX2H
      port map(A => \PIPEA_7[10]\, B => \PIPEA[10]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_599\);
    
    un102_reg_ads_0_a3_0_a2 : NOR2FT
      port map(A => N_674, B => un111_reg_ads_1, Y => 
        \un102_reg_ads_0_a3_0_a2\);
    
    \LB_i_6_1[31]\ : MUX2H
      port map(A => VDB_in(31), B => \LB_DOUT[31]_net_1\, S => 
        \STATE5_0[0]_net_1\, Y => N_2213);
    
    \REG_1[411]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_376\, CLR => 
        \un10_hwres_21\, Q => \REG[411]\);
    
    \REG_1[388]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_353\, CLR => 
        \un10_hwres_19\, Q => \REG[388]\);
    
    \VDBi_23[23]\ : MUX2H
      port map(A => \VDBi_18[23]_net_1\, B => \REG_i[505]_net_1\, 
        S => \REGMAP_1[13]_net_1\, Y => \VDBi_23[23]_net_1\);
    
    \LB_s[24]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_103\, CLR => 
        HWRES_c_18, Q => \LB_s[24]_net_1\);
    
    REG3_127 : MUX2H
      port map(A => \REG[14]\, B => VDB_in(14), S => 
        REG1_0_sqmuxa_0, Y => \REG3_127\);
    
    REG_1_399 : MUX2H
      port map(A => VDB_in(25), B => \REG[434]\, S => N_3072_i_0, 
        Y => \REG_1_399\);
    
    \REG_1[241]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_254\, SET => 
        \un10_hwres_13\, Q => \REG[241]\);
    
    \REG_1_m[234]\ : AND2
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[234]\, Y => 
        \REG_1_m_i[234]\);
    
    \REG_1[128]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_136\, CLR => 
        \un10_hwres_8\, Q => \REG[128]\);
    
    PULSE_1_73 : MUX2H
      port map(A => \PULSE[1]\, B => N_2389, S => N_2454, Y => 
        \PULSE_1_73\);
    
    \VDBi_16_s[1]\ : OR3
      port map(A => N_2461_i, B => \VDBi_16_1_0_i[1]\, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[1]\);
    
    LB_ADDR_551 : MUX2H
      port map(A => \LB_ADDR[8]_net_1\, B => \VAS[8]_net_1\, S
         => LB_ADDR_0_sqmuxa_2, Y => \LB_ADDR_551\);
    
    STATE1_tr12_7_0_o2 : OR3
      port map(A => STATE1_tr12_7_0_o2_4_i, B => 
        STATE1_tr12_7_0_o2_0_i, C => STATE1_tr12_7_0_o2_1_i, Y
         => N_2531);
    
    \VDBi_92_0_iv_0_4[25]\ : AO21TTF
      port map(A => N_790, B => \REG[73]\, C => N_605, Y => 
        \VDBi_92_0_iv_0_4_i[25]\);
    
    PIPEB_24 : MUX2H
      port map(A => \PIPEB[4]_net_1\, B => N_2618, S => N_1996, Y
         => \PIPEB_24\);
    
    \LB_i_6_r[26]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_0, C => N_2208, 
        Y => \LB_i_6[26]\);
    
    \LB_i_6_r[18]\ : AND3
      port map(A => N_2572_2, B => LB_i_6_sn_N_2_1, C => N_2200, 
        Y => \LB_i_6[18]\);
    
    \VADm[18]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[18]_net_1\, Y => 
        VADm(18));
    
    PIPEA1_569 : MUX2H
      port map(A => N_266, B => \PIPEA1[13]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_569\);
    
    PIPEA_597 : MUX2H
      port map(A => \PIPEA_7[8]\, B => \PIPEA[8]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_597\);
    
    \VDBi_16_1_a2_0[5]\ : AND2
      port map(A => N_2511, B => REG_36, Y => N_2473_i);
    
    un1_STATE2_13_i_0 : AO21TTF
      port map(A => N_1762, B => \un1_STATE2_13_i_0_a2_0_0\, C
         => N_581, Y => N_44);
    
    \VDBi[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_624\, CLR => 
        \un10_hwres_35\, Q => \VDBi[3]_net_1\);
    
    \REG_1[399]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_364\, CLR => 
        \un10_hwres_20\, Q => \REG[399]\);
    
    \VDBi_92_0_iv_0[14]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[14]_net_1\, C
         => \PIPEA_m[14]_net_1\, Y => \VDBi_92_0_iv_0[14]_net_1\);
    
    OR_RDATA_183 : MUX2H
      port map(A => N_17, B => \OR_RDATA[1]_net_1\, S => N_1832, 
        Y => \OR_RDATA_183\);
    
    \REG_1[88]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_495\, CLR => 
        \un10_hwres_31\, Q => \REG[88]\);
    
    \VDBi_92_0_iv_0[27]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[27]_net_1\, C
         => \PIPEA_m[27]_net_1\, Y => \VDBi_92_0_iv_0[27]_net_1\);
    
    \VDBi_92_0_iv_0_a2_2[21]\ : NAND2
      port map(A => N_723, B => \REG[430]\, Y => N_587);
    
    \VDBi_16_1_a2_3_0[1]\ : NOR2FT
      port map(A => \REGMAP[1]_net_1\, B => \REGMAP[6]_net_1\, Y
         => \VDBi_16_1_a2_3_0[1]_net_1\);
    
    un5_noe16ri_0_0_a2_0 : NOR2FT
      port map(A => \MBLTCYC\, B => \ADACKCYC\, Y => NOEAD_c);
    
    REG_1_133 : MUX2H
      port map(A => \REG_0[125]\, B => VDB_in(4), S => 
        REG_0_sqmuxa, Y => \REG_1_133\);
    
    un1_TCNT_1_I_44 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1_0[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_2_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\);
    
    \REGMAP[24]\ : DFF
      port map(CLK => CLK_c_c, D => \un81_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[24]_net_1\);
    
    \LB_s[7]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_86\, CLR => HWRES_c_19, 
        Q => \LB_s[7]_net_1\);
    
    VDBi_652 : MUX2H
      port map(A => \VDBi_92[31]\, B => \VDBi[31]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_652\);
    
    N_77_i_i_o2_1 : NOR3
      port map(A => \N_77_i_i_o2_1_0\, B => \PIPEA[29]_net_1\, C
         => \PIPEA[31]_net_1\, Y => N_440);
    
    \LB_DOUT[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_154\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[6]_net_1\);
    
    \VDBi_60[2]\ : MUX2H
      port map(A => \VDBi_60_d[2]_net_1\, B => \VDBi_55[2]_net_1\, 
        S => \VDBi_60_s[5]_net_1\, Y => \VDBi_60[2]_net_1\);
    
    PIPEA1_574 : MUX2H
      port map(A => N_276, B => \PIPEA1[18]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_574\);
    
    \REGMAP[7]\ : DFF
      port map(CLK => CLK_c_c, D => \un33_reg_ads_0_a2_0_a2\, Q
         => \REGMAP[7]_net_1\);
    
    \VDBi[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_647\, CLR => 
        \un10_hwres_35\, Q => \VDBi[26]_net_1\);
    
    LB_i_527 : MUX2H
      port map(A => \LB_i[15]_net_1\, B => \LB_i_6[15]\, S => 
        N_2570_1, Y => \LB_i_527\);
    
    \PIPEB[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_40\, CLR => CLEAR_27, 
        Q => \PIPEB[20]_net_1\);
    
    \PIPEA_7_i_m2[2]\ : MUX2H
      port map(A => DPR(2), B => \PIPEA1[2]_net_1\, S => N_1996_2, 
        Y => N_511);
    
    \PIPEA_7_r[23]\ : AND2
      port map(A => N_85_1, B => N_532, Y => \PIPEA_7[23]\);
    
    un13_reg_ads_0_a2_0_a2_1 : OR2
      port map(A => N_678, B => \VAS[3]_net_1\, Y => 
        un13_reg_ads_1);
    
    LB_i_520 : MUX2H
      port map(A => \LB_i[8]_net_1\, B => \LB_i_6[8]_net_1\, S
         => N_2570, Y => \LB_i_520\);
    
    \PIPEA_7_i_m2[19]\ : MUX2H
      port map(A => DPR(19), B => \PIPEA1[19]_net_1\, S => 
        N_1996_1, Y => N_528);
    
    un74_reg_ads_0_a3_i : INV
      port map(A => \VAS[2]_net_1\, Y => \VAS_i_0[2]\);
    
    \STATE1_0[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[1]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1_0[9]_net_1\);
    
    LB_WRITE : DFFC
      port map(CLK => CLK_c_c, D => \LB_WRITE_68\, CLR => 
        \un10_hwres_3\, Q => \LB_WRITE\);
    
    REG_1_298 : MUX2H
      port map(A => VDB_in(20), B => \REG[285]\, S => N_2880_i, Y
         => \REG_1_298\);
    
    \RAMDTS[7]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(7), CLR => HWRES_c_21, 
        Q => \RAMDTS[7]_net_1\);
    
    \REGMAP_0[7]\ : DFF
      port map(CLK => CLK_c_c, D => \un33_reg_ads_0_a2_0_a2\, Q
         => \REGMAP_0[7]_net_1\);
    
    \STATE1_ns_0_iv_0[2]\ : OAI21TTF
      port map(A => \LB_ACK_sync\, B => LB_DOUT_0_sqmuxa_0, C => 
        \STATE1[0]_net_1\, Y => \STATE1_ns[2]\);
    
    \VDBi_23[3]\ : MUX2H
      port map(A => \VDBi_18[3]_net_1\, B => \REG[485]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23[3]_net_1\);
    
    PIPEA_612 : MUX2H
      port map(A => \PIPEA_7[23]\, B => \PIPEA[23]_net_1\, S => 
        un1_STATE2_16_0, Y => \PIPEA_612\);
    
    \VDBi_77[14]\ : MUX2H
      port map(A => \VDBi_71[14]_net_1\, B => N_2066, S => 
        N_441_0, Y => \VDBi_77[14]_net_1\);
    
    \REG_1_m[264]\ : NAND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[264]\, Y => 
        \REG_1_m[264]_net_1\);
    
    REG_1_421_e : OR2FT
      port map(A => \REGMAP_i_i_0[33]\, B => PULSE_0_sqmuxa_1, Y
         => N_3104_i);
    
    \REG_1_m[189]\ : NAND2
      port map(A => \REGMAP[20]_net_1\, B => \REG[189]\, Y => 
        \REG_1_m[189]_net_1\);
    
    \REG_1[254]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_267\, CLR => 
        \un10_hwres_14\, Q => \REG[254]\);
    
    \STATE5_ns_0_0_a2_1[1]\ : OR2FT
      port map(A => N_2597_1, B => \STATE5_0[0]_net_1\, Y => 
        N_2597);
    
    REG_1_382 : MUX2H
      port map(A => VDB_in_0(8), B => \REG[417]\, S => N_3072_i, 
        Y => \REG_1_382\);
    
    \PIPEB[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_38\, CLR => CLEAR_26, 
        Q => \PIPEB[18]_net_1\);
    
    \REG_i[265]\ : INV
      port map(A => \REG[265]\, Y => REG_i_0_260);
    
    \REG_1[252]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_265\, CLR => 
        \un10_hwres_14\, Q => \REG[252]\);
    
    un1_LBUSTMO_1_I_15 : XOR2FT
      port map(A => N_66, B => \LBUSTMO[2]_net_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[2]\);
    
    \VDBi_92_0_iv[11]\ : OAI21FTT
      port map(A => \VDBi_77[11]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[11]_net_1\, Y => \VDBi_92[11]\);
    
    \PIPEA_m[14]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[14]_net_1\, Y => 
        \PIPEA_m[14]_net_1\);
    
    \REG_1[78]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_485\, CLR => 
        \un10_hwres_30\, Q => \REG[78]\);
    
    \STATE5_ns_0_0_0[0]\ : AO21TTF
      port map(A => \LB_REQ_sync\, B => N_2599_1, C => N_2600, Y
         => \STATE5_ns_0_0_0_i[0]\);
    
    un7_noe32ri_0_0_a2_0 : AND2
      port map(A => N_436, B => N_566_1, Y => 
        \un7_noe32ri_0_0_a2_0\);
    
    PIPEB_28 : MUX2H
      port map(A => \PIPEB[8]_net_1\, B => N_2622, S => N_1996, Y
         => \PIPEB_28\);
    
    REG_1_488 : MUX2H
      port map(A => \REG_88[81]_net_1\, B => \REG[81]\, S => 
        un1_STATE1_15, Y => \REG_1_488\);
    
    REG_1_253 : MUX2H
      port map(A => VDB_in(7), B => \REG[240]\, S => N_2784_i, Y
         => \REG_1_253\);
    
    STATE1_tr27_i_o4_0_o2 : NAND2
      port map(A => \LB_ACK_sync\, B => \REGMAP[36]_net_1\, Y => 
        N_425);
    
    un1_STATE2_13_i_0_a2_0_1 : NOR2
      port map(A => N_485, B => \STATE2[4]_net_1\, Y => N_582_1);
    
    REG_1_273 : MUX2H
      port map(A => VDB_in(11), B => \REG[260]\, S => 
        N_2816_i_0_0, Y => \REG_1_273\);
    
    \WDOG[0]\ : DFFC
      port map(CLK => CLK_c_c, D => 
        \DWACT_ADD_CI_0_partial_sum_1[0]\, CLR => un15_hwres_i, Q
         => \WDOG[0]_net_1\);
    
    \VDBi_53_0_iv_0[5]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_141, C => 
        \REG_1_m[254]_net_1\, Y => \VDBi_53_0_iv_0_i[5]\);
    
    \VDBi_92_iv_0[6]\ : AOI21TTF
      port map(A => \RAMDTS[6]_net_1\, B => \STATE1_0[1]_net_1\, 
        C => \FBOUT_m[6]_net_1\, Y => \VDBi_92_iv_0[6]_net_1\);
    
    \REG_1[188]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_228\, CLR => 
        \un10_hwres_11\, Q => \REG[188]\);
    
    STATE5_0_sqmuxa_0_a3_0_a2_0 : NAND2FT
      port map(A => N_2608, B => N_2606_i_i, Y => 
        STATE5_0_sqmuxa_0);
    
    STATE1_tr27_i_0 : OAI21FTT
      port map(A => \WRITES_1\, B => \STATE1_tr27_i_a2_0_0\, C
         => \STATE1_0[9]_net_1\, Y => \STATE1_tr27_i_0\);
    
    \PIPEA_7_i_m2[14]\ : MUX2H
      port map(A => DPR(14), B => \PIPEA1[14]_net_1\, S => 
        N_1996_1, Y => N_523);
    
    \LB_i_6_r[11]\ : AND2
      port map(A => N_2227, B => N_2572_2, Y => 
        \LB_i_6[11]_net_1\);
    
    REG_1_386 : MUX2H
      port map(A => VDB_in_0(12), B => \REG[421]\, S => 
        N_3072_i_1, Y => \REG_1_386\);
    
    \REG_1[49]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_456\, CLR => 
        \un10_hwres_27\, Q => \REG[49]\);
    
    \VDBm[2]\ : MUX2H
      port map(A => N_2298, B => \VDBi[2]_net_1\, S => \SINGCYC\, 
        Y => VDBm_2);
    
    \REG3[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_116\, CLR => 
        \un10_hwres_6_0\, Q => \REG[3]\);
    
    \VDBi_16_1_a2_0[9]\ : AND2
      port map(A => N_2512_0, B => \REG[9]\, Y => N_2485_i);
    
    \LB_ADDR[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_550\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[7]_net_1\);
    
    \VDBi[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_636\, CLR => 
        \un10_hwres_34\, Q => \VDBi[15]_net_1\);
    
    REG_1_257 : MUX2H
      port map(A => VDB_in(11), B => \REG[244]\, S => N_2784_i_0, 
        Y => \REG_1_257\);
    
    \VDBi_53_0_iv_3[7]\ : AO21TTF
      port map(A => \REGMAP[16]_net_1\, B => \REG[128]\, C => 
        \VDBi_53_0_iv_2[7]_net_1\, Y => \VDBi_53_0_iv_3_i[7]\);
    
    WDOG_3_I_34 : AND2
      port map(A => \WDOG[2]_net_1\, B => \WDOG[3]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    \PIPEA[28]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEA_617\, SET => CLEAR_25, 
        Q => \PIPEA_i_0_i[28]\);
    
    REG_1_277 : MUX2H
      port map(A => VDB_in(15), B => \REG[264]\, S => 
        N_2816_i_0_0, Y => \REG_1_277\);
    
    PURGED_14 : OA21
      port map(A => \EVREAD\, B => \PURGED\, C => un22_bltcyc, Y
         => \PURGED_14\);
    
    \VDBi_16_1_a2_0[12]\ : AND2
      port map(A => N_2512_0, B => \REG[12]\, Y => N_2491_i);
    
    \OR_RDATA_5_i[6]\ : AND2
      port map(A => N_2572, B => LB_in(6), Y => N_2568);
    
    \STATE1_ns_0_iv_0[6]\ : OAI21FTF
      port map(A => \STATE1[4]_net_1\, B => \TST_c_0[2]\, C => 
        N_2612, Y => \STATE1_ns[6]\);
    
    \VDBi_92_0_iv_0[24]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[24]_net_1\, C
         => \PIPEA_m[24]_net_1\, Y => \VDBi_92_0_iv_0[24]_net_1\);
    
    un54_reg_ads_0_a3_0_a2 : AND2
      port map(A => N_682, B => N_675, Y => 
        \un54_reg_ads_0_a3_0_a2\);
    
    \VDBi_23[11]\ : MUX2H
      port map(A => \VDBi_18[11]_net_1\, B => \REG[493]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23[11]_net_1\);
    
    REG_1_308 : MUX2H
      port map(A => VDB_in(30), B => \REG[295]\, S => N_2880_i_0, 
        Y => \REG_1_308\);
    
    \REG_1[401]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_366\, CLR => 
        \un10_hwres_20\, Q => \REG[401]\);
    
    \LB_DOUT[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_170\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[22]_net_1\);
    
    VDBi_628 : MUX2H
      port map(A => \VDBi_92[7]\, B => \VDBi[7]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_628\);
    
    \PIPEA1[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_578\, CLR => CLEAR_21, 
        Q => \PIPEA1[22]_net_1\);
    
    \PIPEA1[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_572\, CLR => CLEAR_21, 
        Q => \PIPEA1[16]_net_1\);
    
    un1_STATE1_20_1_i_0_a2_0_a2 : OR2
      port map(A => \STATE1[10]_net_1\, B => \STATE1[9]_net_1\, Y
         => N_1698);
    
    LB_s_109 : MUX2H
      port map(A => LB_in(30), B => \LB_s[30]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_109\);
    
    REG_1_140 : MUX2H
      port map(A => \REG[132]\, B => VDB_in(11), S => 
        REG_0_sqmuxa_0, Y => \REG_1_140\);
    
    \LB_i_6_1[25]\ : MUX2H
      port map(A => VDB_in(25), B => \LB_DOUT[25]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2207);
    
    \REG_1[289]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_302\, CLR => 
        \un10_hwres_16\, Q => \REG[289]\);
    
    \VDBi_71[19]\ : MUX2H
      port map(A => \VDBi_60[19]_net_1\, B => \REG[428]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[19]_net_1\);
    
    \VDBi_66_0[2]\ : MUX2H
      port map(A => \REG[395]\, B => \REG[379]\, S => 
        \REGMAP[29]_net_1\, Y => N_2019);
    
    \STATE5_ns_0_0[1]\ : NAND3FTT
      port map(A => \STATE5_ns_0_0_0_i[1]\, B => N_2595, C => 
        N_2596, Y => \STATE5_ns[1]\);
    
    \STATE2_ns_0_0_o2[3]\ : OR3FTT
      port map(A => \REGMAP[0]_net_1\, B => \ADACKCYC\, C => 
        \TST_c[2]\, Y => N_449);
    
    REG_1_415 : MUX2H
      port map(A => VDB_in_0(9), B => \REG[450]\, S => N_3104_i_0, 
        Y => \REG_1_415\);
    
    \STATE2_ns_0_0_0[3]\ : AOI21TTF
      port map(A => N_449, B => \STATE2[2]_net_1\, C => 
        \STATE2_i_0[3]\, Y => \STATE2_ns_0_0_0[3]_net_1\);
    
    \VDBi_53_0_iv_5[5]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[5]\, B => 
        \VDBi_53_0_iv_0_i[5]\, C => \VDBi_53_0_iv_1_i[5]\, Y => 
        \VDBi_53_0_iv_5_i[5]\);
    
    \VADm[17]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[17]_net_1\, Y => VADm(17));
    
    \VDBi_60[16]\ : MUX2H
      port map(A => \VDBi_55[16]_net_1\, B => LBSP_in_16, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[16]_net_1\);
    
    PIPEB_20 : MUX2H
      port map(A => \PIPEB[0]_net_1\, B => N_2614, S => N_1996, Y
         => \PIPEB_20\);
    
    \VDBi_77[9]\ : MUX2H
      port map(A => \VDBi_71[9]_net_1\, B => N_2061, S => \N_441\, 
        Y => \VDBi_77[9]_net_1\);
    
    \REG_1[129]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_137\, CLR => 
        \un10_hwres_8\, Q => \REG[129]\);
    
    \STATE2_i[4]\ : INV
      port map(A => \STATE2[4]_net_1\, Y => \STATE2_i[4]_net_1\);
    
    \VDBi_16_r[8]\ : OA21TTF
      port map(A => \VDBi_16_1_0_i[8]\, B => N_2482_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[8]\);
    
    \VDBi_60_d[0]\ : MUX2H
      port map(A => \VDBi_58_d[0]_net_1\, B => LBSP_in_0, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60_d[0]_net_1\);
    
    \STATE1_ns_1_iv_0_a2[3]\ : NAND2FT
      port map(A => N_2531, B => N_83_0, Y => N_2544);
    
    LB_nOE_15 : MUX2H
      port map(A => N_2573, B => LB_nOE_net_1, S => un1_STATE5_8, 
        Y => \LB_nOE_15\);
    
    \VDBi_60[30]\ : MUX2H
      port map(A => \VDBi_55[30]_net_1\, B => LBSP_in_30, S => 
        \REGMAP_0[28]_net_1\, Y => \VDBi_60[30]_net_1\);
    
    \REG_1[263]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_276\, CLR => 
        \un10_hwres_15\, Q => \REG[263]\);
    
    \REG_88[83]\ : NOR2FT
      port map(A => N_2154, B => N_2566, Y => \REG_88[83]_net_1\);
    
    \VDBi_16_1_a2_1[1]\ : NAND2
      port map(A => N_2512, B => \REG[1]\, Y => N_2462);
    
    \TCNT_10_r[5]\ : OA21FTT
      port map(A => \N_1897\, B => I_33_1, C => N_2523_0, Y => 
        \TCNT_10[5]\);
    
    \LB_s[16]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_95\, CLR => HWRES_c_17, 
        Q => \LB_s[16]_net_1\);
    
    \VDBi_71[1]\ : MUX2H
      port map(A => \VDBi_71_d_0[1]_net_1\, B => 
        \VDBi_55[1]_net_1\, S => \VDBi_71_s_0[1]_net_1\, Y => 
        \VDBi_71[1]_net_1\);
    
    \PIPEA[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_597\, CLR => CLEAR_25, 
        Q => \PIPEA[8]_net_1\);
    
    un33_reg_ads_0_a2_0_a2 : NOR2
      port map(A => N_684_i, B => un33_reg_ads_1, Y => 
        \un33_reg_ads_0_a2_0_a2\);
    
    \PIPEA_7_s[28]\ : OR2FT
      port map(A => N_85_0, B => N_537, Y => \PIPEA_7[28]\);
    
    \VDBm[3]\ : MUX2H
      port map(A => N_2299, B => \VDBi[3]_net_1\, S => \SINGCYC\, 
        Y => VDBm_3);
    
    STATE1_tr27_i : NOR3
      port map(A => N_2532, B => N_2561, C => \STATE1_tr27_i_0\, 
        Y => N_43);
    
    PIPEA_608 : MUX2H
      port map(A => \PIPEA_7[19]\, B => \PIPEA[19]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_608\);
    
    WDOGRES_i : INV
      port map(A => \WDOGRES\, Y => \WDOGRES_i\);
    
    \VADm[15]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[15]_net_1\, Y => VADm(15));
    
    REG_1_419 : MUX2H
      port map(A => VDB_in_0(13), B => \REG[454]\, S => 
        N_3104_i_0, Y => \REG_1_419\);
    
    LB_DOUT_166 : MUX2H
      port map(A => VDB_in(18), B => \LB_DOUT[18]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_166\);
    
    \PIPEB_4_i[21]\ : AND2
      port map(A => DPR(21), B => N_616_0, Y => N_2633);
    
    \REG_1_m[170]\ : NAND2
      port map(A => \REGMAP[19]_net_1\, B => \REG[170]\, Y => 
        \REG_1_m[170]_net_1\);
    
    un1_LB_DOUT_0_sqmuxa_0_a2 : NAND2
      port map(A => \STATE1[5]_net_1\, B => \TST_c[0]\, Y => 
        N_2429);
    
    \VDBi_55[29]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[29]_net_1\, Y => \VDBi_55[29]_net_1\);
    
    WDOGCLEAR_69 : MUX2H
      port map(A => \STATE1[8]_net_1\, B => \WDOGCLEAR\, S => 
        un1_STATE1_29, Y => \WDOGCLEAR_69\);
    
    \VDBi_92_iv_2[2]\ : AOI21TTF
      port map(A => \LB_s[2]_net_1\, B => N_7_i, C => 
        \VDBi_92_iv_1[2]_net_1\, Y => \VDBi_92_iv_2[2]_net_1\);
    
    un1_WDOGRES_0_sqmuxa_0_a2_0_3 : NAND3FFT
      port map(A => \WDOG_i_0_i[4]\, B => \WDOG[5]_net_1\, C => 
        \un1_WDOGRES_0_sqmuxa_0_a2_0_i\, Y => 
        un1_WDOGRES_0_sqmuxa_0_a2_0_3_i);
    
    \PIPEA1[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_556\, CLR => CLEAR_20, 
        Q => \PIPEA1[0]_net_1\);
    
    \LBUSTMO[1]\ : DFFS
      port map(CLK => ALICLK_c, D => \LBUSTMO_3[1]\, SET => 
        HWRES_c_13_0, Q => \LBUSTMO_i_0_i[1]\);
    
    PIPEB_25 : MUX2H
      port map(A => \PIPEB[5]_net_1\, B => N_2619, S => N_1996, Y
         => \PIPEB_25\);
    
    REG_1_420 : MUX2H
      port map(A => VDB_in_0(14), B => \REG[455]\, S => 
        N_3104_i_0, Y => \REG_1_420\);
    
    \VDBi_60[7]\ : MUX2H
      port map(A => \VDBi_58[7]_net_1\, B => L2A_c_c, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60[7]_net_1\);
    
    un1_TCNT_1_I_16 : XOR2
      port map(A => \TCNT_i_i[6]\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_5[0]\);
    
    VSEL_0_a2 : NOR2FT
      port map(A => N_2403, B => \TST_c_0[0]\, Y => \TST_c[1]\);
    
    \VDBi_66[11]\ : MUX2H
      port map(A => \VDBi_66_d[11]_net_1\, B => 
        \VDBi_58[11]_net_1\, S => \VDBi_66_s[1]_net_1\, Y => 
        \VDBi_66[11]_net_1\);
    
    \VDBi_16_1_1[0]\ : AO21TTF
      port map(A => N_2380_1, B => \VDBi_16_1_a3_1_0[0]_net_1\, C
         => \VDBi_16_1_0[0]_net_1\, Y => \VDBi_16_1_1_i[0]\);
    
    \REG_1_0[124]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_132\, CLR => 
        \un10_hwres_7_0\, Q => \REG_0[124]\);
    
    LB_s_93 : MUX2H
      port map(A => LB_in(14), B => \LB_s[14]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_93\);
    
    \PIPEA1[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_560\, CLR => CLEAR_22, 
        Q => \PIPEA1[4]_net_1\);
    
    \un7_noe32ri_0_0\ : OAI21FTF
      port map(A => \un7_noe32ri_0_0_a2_0\, B => \LWORDS\, C => 
        \NOEAD_c_0\, Y => un7_noe32ri_0_0);
    
    REG_1_325 : MUX2H
      port map(A => VDB_in_0(15), B => \REG[360]\, S => N_2944_i, 
        Y => \REG_1_325\);
    
    un1_anycyc_i_0_o2_i_a2_0 : OR2
      port map(A => \SINGCYC_0\, B => \BLTCYC_0\, Y => N_2507_0);
    
    \REG_1[103]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_510\, CLR => 
        \un10_hwres_7\, Q => \REG[103]\);
    
    \LB_i[19]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_531\, CLR => 
        HWRES_c_15, Q => \LB_i[19]_net_1\);
    
    VDBi_623 : MUX2H
      port map(A => \VDBi_92[2]\, B => \VDBi[2]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_623\);
    
    PIPEA1_579 : MUX2H
      port map(A => N_286, B => \PIPEA1[23]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_579\);
    
    \REGMAP[6]\ : DFF
      port map(CLK => CLK_c_c, D => \un29_reg_ads_0_a2_0_a2\, Q
         => \REGMAP[6]_net_1\);
    
    REG_1_208_e : OR2FT
      port map(A => \REGMAP_0[18]_net_1\, B => PULSE_0_sqmuxa_1_2, 
        Y => N_2688_i);
    
    \REG_1[431]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_396\, CLR => 
        \un10_hwres_23\, Q => \REG[431]\);
    
    \REG_1[170]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_210\, CLR => 
        \un10_hwres_10\, Q => \REG[170]\);
    
    \REG_1_m[158]\ : NAND2
      port map(A => \REGMAP[18]_net_1\, B => \REG[158]\, Y => 
        \REG_1_m[158]_net_1\);
    
    REG_1_465 : MUX2H
      port map(A => VDB_in_0(10), B => \REG[58]\, S => N_3234_i_1, 
        Y => \REG_1_465\);
    
    REG_1_sqmuxa_1_i_o2 : AND2
      port map(A => \TST_c_0[5]\, B => \STATE1_0[8]_net_1\, Y => 
        N_2409);
    
    REG_1_352 : MUX2H
      port map(A => VDB_in_0(10), B => \REG[387]\, S => 
        N_2976_i_0, Y => \REG_1_352\);
    
    WDOGTOi_0 : DFFC
      port map(CLK => CLK_c_c, D => \un12_wdog_0_a3\, CLR => 
        un15_hwres_i, Q => WDOGTO_0);
    
    \LB_i[30]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_542\, CLR => 
        HWRES_c_16, Q => \LB_i[30]_net_1\);
    
    un5_noe16ri_0_0_i : INV
      port map(A => \NOEAD_c_0\, Y => NOEAD_c_i_0);
    
    \PIPEB_4_i_a2_1[0]\ : NAND2
      port map(A => N_428, B => \STATE2_i_0[3]\, Y => N_616_1);
    
    \VDBi_16_r[3]\ : OA21TTF
      port map(A => \VDBi_16_1_0_i[3]\, B => N_2467_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[3]\);
    
    STATE1_tr27_i_a2_0_0 : OR2FT
      port map(A => \REGMAP[15]_net_1\, B => \REGMAP[36]_net_1\, 
        Y => \STATE1_tr27_i_a2_0_0\);
    
    \PIPEA1_9_i[10]\ : AND2
      port map(A => DPR(10), B => N_85_4, Y => N_260);
    
    REG_1_372 : MUX2H
      port map(A => VDB_in_0(14), B => \REG[407]\, S => 
        N_3008_i_0, Y => \REG_1_372\);
    
    REG_1_458 : MUX2H
      port map(A => VDB_in_0(3), B => \REG[51]\, S => N_3234_i, Y
         => \REG_1_458\);
    
    \VDBi_60_s[5]\ : NOR2
      port map(A => \REGMAP[27]_net_1\, B => \REGMAP[28]_net_1\, 
        Y => \VDBi_60_s[5]_net_1\);
    
    \TCNT_10_0_a2[6]\ : AND2
      port map(A => N_2397, B => I_27, Y => \TCNT_10[6]\);
    
    \OR_RDATA_5_i[1]\ : AND2
      port map(A => N_2572, B => LB_in(1), Y => N_17);
    
    un4_asb_3 : XOR2FT
      port map(A => GA_c(3), B => VAD_in_30, Y => \un4_asb_3\);
    
    \REG3_0[514]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_514_180\, CLR => 
        \un10_hwres_0\, Q => RUN_c_0);
    
    REG_1_478 : MUX2H
      port map(A => VDB_in(23), B => \REG[71]\, S => N_3234_i_0, 
        Y => \REG_1_478\);
    
    REG3_514_180 : MUX2H
      port map(A => \REG1_15[514]_net_1\, B => \RUN_c\, S => 
        \REG1_1_sqmuxa\, Y => \REG3_514_180\);
    
    \PIPEA_7_r[6]\ : AND2
      port map(A => N_85_2, B => N_515, Y => \PIPEA_7[6]\);
    
    \PIPEA[30]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEA_619\, SET => CLEAR_25, 
        Q => \PIPEA[30]_net_1\);
    
    \OR_RDATA_5_i[7]\ : AND2
      port map(A => N_2572, B => LB_in(7), Y => N_29);
    
    PIPEA_598 : MUX2H
      port map(A => \PIPEA_7[9]\, B => \PIPEA[9]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_598\);
    
    LB_i_525 : MUX2H
      port map(A => \LB_i[13]_net_1\, B => \LB_i_6[13]\, S => 
        N_2570_1, Y => \LB_i_525\);
    
    EVREAD_DS : DFFC
      port map(CLK => CLK_c_c, D => \EVREAD_DS_145\, CLR => 
        CLEAR_20, Q => \EVREAD_DS\);
    
    VDBi_646 : MUX2H
      port map(A => \VDBi_92[25]\, B => \VDBi[25]_net_1\, S => 
        \un1_STATE1_34_0\, Y => \VDBi_646\);
    
    \REG_1_m[160]\ : NAND2
      port map(A => \REGMAP[18]_net_1\, B => \REG[160]\, Y => 
        \REG_1_m[160]_net_1\);
    
    PIPEA1_557 : MUX2H
      port map(A => N_242, B => \PIPEA1[1]_net_1\, S => 
        un1_STATE2_13_4, Y => \PIPEA1_557\);
    
    \VDBi[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_633\, CLR => 
        \un10_hwres_33\, Q => \VDBi[12]_net_1\);
    
    \REG_1[189]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_229\, CLR => 
        \un10_hwres_11\, Q => \REG[189]\);
    
    REG_1_356 : MUX2H
      port map(A => VDB_in_0(14), B => \REG[391]\, S => 
        N_2976_i_0, Y => \REG_1_356\);
    
    \VDBi_53_0_iv_1[12]\ : AO21TTF
      port map(A => \REGMAP_i_i[23]\, B => \REG[245]\, C => 
        \REG_1_m[197]_net_1\, Y => \VDBi_53_0_iv_1_i[12]\);
    
    \STATE5_ns_i_0_a2_0[2]\ : OR3FFT
      port map(A => \STATE5[1]_net_1\, B => \STATE5_0[2]_net_1\, 
        C => \OR_RREQ_sync\, Y => N_2593_i);
    
    REG_1_376 : MUX2H
      port map(A => VDB_in_0(2), B => \REG[411]\, S => N_3072_i, 
        Y => \REG_1_376\);
    
    \VDBi_18[3]\ : MUX2H
      port map(A => \VDBi_16[3]\, B => \REG[51]\, S => \TST_c[5]\, 
        Y => \VDBi_18[3]_net_1\);
    
    REG_1_496 : MUX2H
      port map(A => \REG[89]\, B => VDB_in_0(0), S => N_2416_i, Y
         => \REG_1_496\);
    
    REG_1_469 : MUX2H
      port map(A => VDB_in_0(14), B => \REG[62]\, S => N_3234_i_1, 
        Y => \REG_1_469\);
    
    LB_i_517 : MUX2H
      port map(A => \LB_i[5]_net_1\, B => \LB_i_6[5]_net_1\, S
         => N_2570, Y => \LB_i_517\);
    
    un1_STATE2_13_i_0_o2_0 : OA21FTT
      port map(A => \TST_c_0[2]\, B => \END_PK\, C => 
        \STATE2[1]_net_1\, Y => N_450_i);
    
    \REG_1_m[253]\ : NAND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[253]\, Y => 
        \REG_1_m[253]_net_1\);
    
    \REG_1_m[166]\ : NAND2
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[166]\, Y => 
        \REG_1_m[166]_net_1\);
    
    \VDBi_23[2]\ : MUX2H
      port map(A => \VDBi_18[2]_net_1\, B => \REG[484]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23[2]_net_1\);
    
    REG_1_250 : MUX2H
      port map(A => VDB_in(4), B => \REG[237]\, S => N_2784_i, Y
         => \REG_1_250\);
    
    LB_DOUT_169 : MUX2H
      port map(A => VDB_in(21), B => \LB_DOUT[21]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_169\);
    
    REG_1_384 : MUX2H
      port map(A => VDB_in_0(10), B => \REG[419]\, S => 
        N_3072_i_1, Y => \REG_1_384\);
    
    \VDBi_77_0[2]\ : MUX2H
      port map(A => REG_458, B => \REG[443]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_2054);
    
    \PIPEA_7_i_m2[30]\ : MUX2H
      port map(A => DPR(30), B => \PIPEA1[30]_net_1\, S => 
        N_1996_0, Y => N_539);
    
    REG_1_270 : MUX2H
      port map(A => VDB_in(8), B => \REG[257]\, S => N_2816_i_0_0, 
        Y => \REG_1_270\);
    
    REG_1_209 : MUX2H
      port map(A => VDB_in(0), B => \REG[169]\, S => N_2720_i, Y
         => \REG_1_209\);
    
    VAS_52 : MUX2H
      port map(A => \VAS[1]_net_1\, B => VAD_in_0, S => 
        \TST_c[1]\, Y => \VAS_52\);
    
    un67_reg_ads_0_a3_0_a2 : NOR2FT
      port map(A => N_675, B => N_683_i, Y => 
        \un67_reg_ads_0_a3_0_a2\);
    
    \VDBi_23[27]\ : MUX2H
      port map(A => \VDBi_18[27]_net_1\, B => \REG_i[509]_net_1\, 
        S => \REGMAP_0[13]_net_1\, Y => \VDBi_23[27]_net_1\);
    
    LB_WRITE_68 : MUX2H
      port map(A => \LB_WRITE\, B => \STATE1[8]_net_1\, S => 
        N_2384, Y => \LB_WRITE_68\);
    
    \PIPEA_7_r[1]\ : AND2
      port map(A => N_85_3, B => N_510, Y => \PIPEA_7[1]\);
    
    REG_1_233 : MUX2H
      port map(A => VDB_in(8), B => \REG[193]\, S => N_2752_i_0, 
        Y => \REG_1_233\);
    
    \OR_RDATA[8]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_190\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[8]_net_1\);
    
    REG_1_487 : MUX2H
      port map(A => \REG[80]\, B => VDB_in_0(0), S => N_3236_i, Y
         => \REG_1_487\);
    
    \OR_RDATA[2]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_184\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[2]_net_1\);
    
    \LB_i[14]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_526\, CLR => 
        HWRES_c_14, Q => \LB_i[14]_net_1\);
    
    \REGMAP[3]\ : DFF
      port map(CLK => CLK_c_c, D => \un17_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_0_i[3]\);
    
    \PIPEA1[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_558\, CLR => CLEAR_22, 
        Q => \PIPEA1[2]_net_1\);
    
    \VDBi_92_0_iv_1[26]\ : AOI21TTF
      port map(A => \LB_s[26]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[26]_net_1\, Y => 
        \VDBi_92_0_iv_1[26]_net_1\);
    
    \REG_1[496]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_437\, SET => 
        \un10_hwres_26\, Q => \REG[496]\);
    
    \LB_i_6_r[27]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_0, C => N_2209, 
        Y => \LB_i_6[27]\);
    
    \REG_1[453]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_418\, CLR => 
        \un10_hwres_25\, Q => \REG[453]\);
    
    \LB_s[11]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_90\, CLR => HWRES_c_17, 
        Q => \LB_s[11]_net_1\);
    
    \VDBi_92_0_iv_0_a2_7[21]\ : NAND2
      port map(A => \LB_s[21]_net_1\, B => N_7_i_0, Y => N_592);
    
    \VDBi_55[23]\ : NOR2
      port map(A => \REGMAP_0[26]_net_1\, B => 
        \VDBi_23[23]_net_1\, Y => \VDBi_55[23]_net_1\);
    
    \LB_ADDR[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_552\, CLR => 
        \un10_hwres_1\, Q => \LB_ADDR[9]_net_1\);
    
    \REG_1[286]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_299\, CLR => 
        \un10_hwres_16\, Q => \REG[286]\);
    
    \VDBi_53_0_iv_0[12]\ : AO21TTF
      port map(A => \REGMAP[12]_net_1\, B => REG_116, C => 
        \REG_1_m[261]_net_1\, Y => \VDBi_53_0_iv_0_i[12]\);
    
    \VDBi_55[20]\ : NOR2
      port map(A => \REGMAP[26]_net_1\, B => \VDBi_23[20]_net_1\, 
        Y => \VDBi_55[20]_net_1\);
    
    REG_1_237 : MUX2H
      port map(A => VDB_in(12), B => \REG[197]\, S => N_2752_i_0, 
        Y => \REG_1_237\);
    
    \PIPEA_m[19]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[19]_net_1\, Y => 
        \PIPEA_m[19]_net_1\);
    
    \PIPEB_4_i[20]\ : AND2
      port map(A => DPR(20), B => N_616_1, Y => N_2632);
    
    LB_s_89 : MUX2H
      port map(A => LB_in(10), B => \LB_s[10]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_89\);
    
    un7_noe32ri_0_0_a2_1 : NOR2FT
      port map(A => \WRITES_0\, B => \DS_i_a2\, Y => N_566_1);
    
    \PULSE_1[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_74\, CLR => 
        \un10_hwres_4\, Q => \PULSE[2]\);
    
    \VDBi[28]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_649\, CLR => 
        \un10_hwres_35\, Q => \VDBi[28]_net_1\);
    
    LB_DOUT_160 : MUX2H
      port map(A => VDB_in(12), B => \LB_DOUT[12]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_160\);
    
    un29_reg_ads_0_a2_0_a2_0 : OR2FT
      port map(A => N_660, B => \VAS[6]_net_1\, Y => N_662);
    
    \VDBi[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_628\, CLR => 
        \un10_hwres\, Q => \VDBi[7]_net_1\);
    
    \VDBi_23[26]\ : MUX2H
      port map(A => \VDBi_18[26]_net_1\, B => \REG_i[508]_net_1\, 
        S => \REGMAP_0[13]_net_1\, Y => \VDBi_23[26]_net_1\);
    
    \TCNT_10_0_a2[3]\ : AND2
      port map(A => N_2397, B => I_30_2, Y => \TCNT_10[3]\);
    
    \VDBi_92_0_iv[26]\ : OAI21FTT
      port map(A => \VDBi_71[26]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[26]_net_1\, Y => \VDBi_92[26]\);
    
    OR_RDATA_182 : MUX2H
      port map(A => N_13, B => \OR_RDATA[0]_net_1\, S => N_1832, 
        Y => \OR_RDATA_182\);
    
    nLBASi_3 : MUX2H
      port map(A => LB_i_6_sn_N_2, B => \nLBAS_c\, S => 
        \STATE5[2]_net_1\, Y => \nLBASi_3\);
    
    \PIPEB_4_i[8]\ : AND2
      port map(A => DPR(8), B => N_616, Y => N_2622);
    
    \VDBi_92_0_iv_0_4[31]\ : AO21TTF
      port map(A => N_790, B => \REG[79]\, C => N_612, Y => 
        \VDBi_92_0_iv_0_4_i[31]\);
    
    \REG_1[362]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_327\, CLR => 
        \un10_hwres_17\, Q => \REG[362]\);
    
    \REG_1[133]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_141\, CLR => 
        \un10_hwres_8_0\, Q => \REG[133]\);
    
    REG3_115 : MUX2H
      port map(A => \REG[2]\, B => VDB_in(2), S => REG1_0_sqmuxa, 
        Y => \REG3_115\);
    
    \LB_DOUT[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_155\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[7]_net_1\);
    
    REG_1_482 : MUX2H
      port map(A => VDB_in(27), B => \REG[75]\, S => N_3234_i_0, 
        Y => \REG_1_482\);
    
    \LB_DOUT[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_162\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[14]_net_1\);
    
    \VDBi_71[24]\ : MUX2H
      port map(A => \VDBi_60[24]_net_1\, B => \REG[433]\, S => 
        \REGMAP_1[31]_net_1\, Y => \VDBi_71[24]_net_1\);
    
    \LB_i_6_1[0]\ : MUX2H
      port map(A => VDB_in_0(0), B => \LB_DOUT[0]_net_1\, S => 
        \STATE5[0]_net_1\, Y => N_2182);
    
    \REG_1[424]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_389\, CLR => 
        \un10_hwres_22\, Q => \REG[424]\);
    
    \LB_i_6_0[2]\ : MUX2H
      port map(A => OR_RADDR(0), B => \LB_ADDR[2]_net_1\, S => 
        \STATE5[0]_net_1\, Y => N_2172);
    
    \VDBi_55[18]\ : NOR2FT
      port map(A => \VDBi_23[18]_net_1\, B => 
        \REGMAP_0[26]_net_1\, Y => \VDBi_55[18]_net_1\);
    
    \LB_i_6_1[13]\ : MUX2H
      port map(A => VDB_in_0(13), B => \LB_DOUT[13]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2195);
    
    VDBi_625 : MUX2H
      port map(A => \VDBi_92[4]\, B => \VDBi[4]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_625\);
    
    WDOGTOi : DFFC
      port map(CLK => CLK_c_c, D => \un12_wdog_0_a3\, CLR => 
        un15_hwres_i, Q => \WDOGTO\);
    
    \VDBi_23[22]\ : MUX2H
      port map(A => \VDBi_18[22]_net_1\, B => \REG_i[504]_net_1\, 
        S => \REGMAP_1[13]_net_1\, Y => \VDBi_23[22]_net_1\);
    
    \REG_88_0[82]\ : MUX2H
      port map(A => VDB_in_0(1), B => \REG[82]\, S => N_20, Y => 
        N_2153);
    
    \REG_1[121]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_129\, SET => 
        \un10_hwres_7_0\, Q => \REG[121]\);
    
    RAMAD_VME_11 : MUX2H
      port map(A => \VAS[8]_net_1\, B => \RAMAD_VME[7]_net_1\, S
         => N_2523_0, Y => \RAMAD_VME_11\);
    
    \VDBi_92_0_iv_0_0_0[21]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[21]_net_1\, C
         => N_587, Y => \VDBi_92_0_iv_0_0_0[21]_net_1\);
    
    \REG_1[366]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_331\, CLR => 
        \un10_hwres_17\, Q => \REG[366]\);
    
    \REGMAP[16]\ : DFF
      port map(CLK => CLK_c_c, D => \un54_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[16]_net_1\);
    
    \PIPEA1_9_i[4]\ : AND2
      port map(A => DPR(4), B => N_85, Y => N_248);
    
    VDBi_627 : MUX2H
      port map(A => \VDBi_92[6]\, B => \VDBi[6]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_627\);
    
    VSEL_0_a2_0 : NOR2FT
      port map(A => N_2403, B => \TST_c_0[0]\, Y => \TST_c_0[1]\);
    
    un1_LBUSTMO_1_I_1 : NOR2FT
      port map(A => \LBUSTMO_i_0_i[0]\, B => N_66, Y => 
        \DWACT_ADD_CI_0_TMP_0[0]\);
    
    \STATE1_ns_0_iv_0_0_0[1]\ : OAI21FTT
      port map(A => N_479, B => \SINGCYC_0\, C => N_629, Y => 
        \STATE1_ns_0_iv_0_0_0_i[1]\);
    
    \REG_1[511]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_452\, CLR => 
        \un10_hwres_28\, Q => \REG[511]\);
    
    \VDBi_16_1_a2_0[4]\ : AND2
      port map(A => N_2511, B => REG_35, Y => N_2470_i);
    
    \VDBi_53_0_iv_1[13]\ : AO21TTF
      port map(A => \REGMAP_i_i[23]\, B => \REG[246]\, C => 
        \REG_1_m[198]_net_1\, Y => \VDBi_53_0_iv_1_i[13]\);
    
    CYCS1 : DFFC
      port map(CLK => CLK_c_c, D => \un7_cycs_0_a2\, CLR => 
        HWRES_c_13, Q => \CYCS1\);
    
    \REG_1[260]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_273\, CLR => 
        \un10_hwres_15\, Q => \REG[260]\);
    
    \VDBi_16_r[9]\ : OA21TTF
      port map(A => N_2485_i, B => N_2484_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[9]\);
    
    un1_STATE1_15_0 : NAND2
      port map(A => N_231, B => N_446, Y => un1_STATE1_15);
    
    REG_1_341_e : OR2FT
      port map(A => \REGMAP_0[28]_net_1\, B => PULSE_0_sqmuxa_1, 
        Y => N_2944_i);
    
    \PIPEA_7_i_m2[6]\ : MUX2H
      port map(A => DPR(6), B => \PIPEA1[6]_net_1\, S => N_1996_2, 
        Y => N_515);
    
    \REG_1[56]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_463\, CLR => 
        \un10_hwres_28\, Q => \REG[56]\);
    
    PIPEB_32 : MUX2H
      port map(A => \PIPEB[12]_net_1\, B => N_2626, S => N_1996_4, 
        Y => \PIPEB_32\);
    
    \REG3[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_120\, CLR => 
        \un10_hwres_6_0\, Q => \REG[7]\);
    
    \VDBi_92_0_iv_0[8]\ : AOI21TTF
      port map(A => \STATE1[2]_net_1\, B => \VDBi[8]_net_1\, C
         => \PIPEA_m[8]_net_1\, Y => \VDBi_92_0_iv_0[8]_net_1\);
    
    \REG_i[281]\ : INV
      port map(A => \REG[281]\, Y => REG_i_0_276);
    
    LB_i_529 : MUX2H
      port map(A => \LB_i[17]_net_1\, B => \LB_i_6[17]\, S => 
        N_2570_1, Y => \LB_i_529\);
    
    \LB_s[18]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_97\, CLR => HWRES_c_17, 
        Q => \LB_s[18]_net_1\);
    
    \VDBi_92_0_iv_0_0_1[21]\ : AO21TTF
      port map(A => N_457_i_0_0, B => \PIPEA[21]_net_1\, C => 
        N_592, Y => \VDBi_92_0_iv_0_0_1_i[21]\);
    
    REG_1_194 : MUX2H
      port map(A => VDB_in(1), B => \REG[154]\, S => N_2688_i, Y
         => \REG_1_194\);
    
    \VDBi_16_1_0[4]\ : AO21TTF
      port map(A => \REGMAP[2]_net_1\, B => REG_19, C => N_2471, 
        Y => \VDBi_16_1_0_i[4]\);
    
    \VDBi_16_1_a2_1[2]\ : OR3FFT
      port map(A => \REG[2]\, B => \VDBi_16_1_a2_3_0[1]_net_1\, C
         => \REGMAP_0[2]_net_1\, Y => N_2465);
    
    un74_reg_ads_0_a3_1 : NOR3FFT
      port map(A => \VAS_i_0[2]\, B => \WRITES_1\, C => 
        \VAS[1]_net_1\, Y => \un74_reg_ads_0_a3_1\);
    
    un776_regmap_14 : NOR3
      port map(A => \REGMAP_0[2]_net_1\, B => un776_regmap_7_i, C
         => un776_regmap_8_0_i, Y => \un776_regmap_14\);
    
    REG_1_196 : MUX2H
      port map(A => VDB_in(3), B => \REG[156]\, S => N_2688_i, Y
         => \REG_1_196\);
    
    PULSE_1_74 : MUX2H
      port map(A => \PULSE[2]\, B => N_2390, S => N_2454, Y => 
        \PULSE_1_74\);
    
    \VDBi_53_0_iv_0[2]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_138, C => 
        \REG_1_m[251]_net_1\, Y => \VDBi_53_0_iv_0_i[2]\);
    
    PIPEA_605 : MUX2H
      port map(A => \PIPEA_7[16]\, B => \PIPEA[16]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_605\);
    
    \REG_1[192]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_232\, CLR => 
        \un10_hwres_12\, Q => \REG[192]\);
    
    \PIPEA[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_591\, CLR => CLEAR_25, 
        Q => \PIPEA[2]_net_1\);
    
    \VDBi_53_0_iv_0[13]\ : AO21TTF
      port map(A => \REGMAP[12]_net_1\, B => REG_117, C => 
        \REG_1_m[262]_net_1\, Y => \VDBi_53_0_iv_0_i[13]\);
    
    BLTCYC_77 : OA21TTF
      port map(A => N_2434_i, B => \BLTCYC_0\, C => \TST_c_0[0]\, 
        Y => \BLTCYC_77\);
    
    WDOG_3_I_21 : XOR2
      port map(A => \WDOG[1]_net_1\, B => \DWACT_ADD_CI_0_TMP[0]\, 
        Y => \WDOG_3[1]\);
    
    un1_TCNT_1_I_5 : AND2
      port map(A => \TCNT[1]_net_1\, B => N_83, Y => 
        \DWACT_ADD_CI_0_g_array_0_1_0[0]\);
    
    \STATE2_ns_a3_0_a3[5]\ : AND2FT
      port map(A => N_1756, B => \STATE2[5]_net_1\, Y => 
        \STATE2_ns_i[5]\);
    
    \REG_1[194]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_234\, CLR => 
        \un10_hwres_12\, Q => \REG[194]\);
    
    VDBi_630 : MUX2H
      port map(A => \VDBi_92[9]\, B => \VDBi[9]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_630\);
    
    \OR_RDATA_5_i[3]\ : AND2
      port map(A => N_2572, B => LB_in(3), Y => N_21);
    
    \PULSE_1[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_72\, CLR => 
        \un10_hwres_4\, Q => \PULSE[0]\);
    
    \VDBm_0[3]\ : MUX2H
      port map(A => \PIPEB[3]_net_1\, B => \PIPEA[3]_net_1\, S
         => \BLTCYC\, Y => N_2299);
    
    un1_TCNT_1_I_32 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum_0[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, Y => I_32_1);
    
    PIPEA_604 : MUX2H
      port map(A => \PIPEA_7[15]\, B => \PIPEA[15]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_604\);
    
    REG_1_421_e_0 : OR2FT
      port map(A => \REGMAP_i_i_0[33]\, B => PULSE_0_sqmuxa_1_0, 
        Y => N_3104_i_0);
    
    RAMAD_VME_8 : MUX2H
      port map(A => \VAS[5]_net_1\, B => \RAMAD_VME[4]_net_1\, S
         => N_2523_0, Y => \RAMAD_VME_8\);
    
    un114_reg_ads_0_a3_0_a2_1 : NOR2FT
      port map(A => \VAS[5]_net_1\, B => \VAS[2]_net_1\, Y => 
        N_690);
    
    \VDBi_23[24]\ : MUX2H
      port map(A => \VDBi_18[24]_net_1\, B => \REG_i[506]_net_1\, 
        S => \REGMAP_1[13]_net_1\, Y => \VDBi_23[24]_net_1\);
    
    \REG_1[258]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_271\, CLR => 
        \un10_hwres_15\, Q => \REG[258]\);
    
    \REG_1[196]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_236\, CLR => 
        \un10_hwres_12\, Q => \REG[196]\);
    
    \VDBi_18[2]\ : MUX2H
      port map(A => \VDBi_16[2]\, B => \REG[50]\, S => \TST_c[5]\, 
        Y => \VDBi_18[2]_net_1\);
    
    \VADm[20]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[20]_net_1\, Y => 
        VADm(20));
    
    \LBUSTMO[3]\ : DFFS
      port map(CLK => ALICLK_c, D => \LBUSTMO_3[3]\, SET => 
        HWRES_c_13_0, Q => \LBUSTMO_i_0_i[3]\);
    
    \TCNT_10_s[2]\ : AO21TTF
      port map(A => \N_1897\, B => I_32_1, C => 
        \TCNT_0_sqmuxa_i_s\, Y => \TCNT_10[2]\);
    
    un1_TCNT_1_I_19 : XOR2
      port map(A => \TCNT_i_i[0]\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \REG_1[484]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_425\, SET => 
        \un10_hwres_25\, Q => \REG[484]\);
    
    \LB_i_6_1[1]\ : MUX2H
      port map(A => VDB_in_0(1), B => \LB_DOUT[1]_net_1\, S => 
        \STATE5[0]_net_1\, Y => N_2183);
    
    un10_hwres_8 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_8\);
    
    \VDBi_92_0_iv[9]\ : OAI21FTT
      port map(A => \VDBi_77[9]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[9]_net_1\, Y => \VDBi_92[9]\);
    
    WDOGTOi_1 : DFFC
      port map(CLK => CLK_c_c, D => \un12_wdog_0_a3\, CLR => 
        un15_hwres_i, Q => WDOGTO_1);
    
    REG_1_354 : MUX2H
      port map(A => VDB_in_0(12), B => \REG[389]\, S => 
        N_2976_i_0, Y => \REG_1_354\);
    
    LB_s_101 : MUX2H
      port map(A => LB_in(22), B => \LB_s[22]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_101\);
    
    \VDBi_66_0[10]\ : MUX2H
      port map(A => \REG[403]\, B => \REG[387]\, S => 
        \REGMAP_0[29]_net_1\, Y => N_2027);
    
    \REG_1[181]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_221\, CLR => 
        \un10_hwres_11\, Q => \REG[181]\);
    
    un120_reg_ads_0_a3_0_a2 : AND3
      port map(A => un120_reg_ads_1, B => \VAS[2]_net_1\, C => 
        \VAS[5]_net_1\, Y => \un120_reg_ads_0_a3_0_a2\);
    
    REG_1_374 : MUX2H
      port map(A => VDB_in_0(0), B => \REG[409]\, S => N_3072_i, 
        Y => \REG_1_374\);
    
    \REG3[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG3_115\, CLR => 
        \un10_hwres_6\, Q => \REG[2]\);
    
    REG_1_332 : MUX2H
      port map(A => VDB_in(22), B => \REG[367]\, S => N_2944_i_0, 
        Y => \REG_1_332\);
    
    LB_i_541 : MUX2H
      port map(A => \LB_i[29]_net_1\, B => \LB_i_6[29]\, S => 
        N_2570_0, Y => \LB_i_541\);
    
    REG_1_206 : MUX2H
      port map(A => VDB_in(13), B => \REG[166]\, S => N_2688_i_0, 
        Y => \REG_1_206\);
    
    \REG_1_m[159]\ : NAND2
      port map(A => \REGMAP[18]_net_1\, B => \REG[159]\, Y => 
        \REG_1_m[159]_net_1\);
    
    PIPEB_44 : MUX2H
      port map(A => \PIPEB[24]_net_1\, B => N_2635, S => N_1996_3, 
        Y => \PIPEB_44\);
    
    \VDBi_92_0_iv_0[16]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[16]_net_1\, C
         => \PIPEA_m[16]_net_1\, Y => \VDBi_92_0_iv_0[16]_net_1\);
    
    un5_noe16ri_0_0_a2_0_0_0 : NOR2FT
      port map(A => \MBLTCYC\, B => \ADACKCYC\, Y => 
        \NOEAD_c_0_0\);
    
    REG_1_438 : MUX2H
      port map(A => VDB_in_0(15), B => \REG[497]\, S => 
        N_3170_i_1, Y => \REG_1_438\);
    
    \VDBi_53_0_iv_1[6]\ : AO21TTF
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[239]\, C => 
        \REG_1_m[191]_net_1\, Y => \VDBi_53_0_iv_1_i[6]\);
    
    \PIPEA1_9_i[25]\ : AND2
      port map(A => DPR(25), B => N_85_3, Y => N_290);
    
    \OR_RDATA_5_i[0]\ : AND2
      port map(A => N_2572, B => LB_in(0), Y => N_13);
    
    \LB_ADDR[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_544\, CLR => 
        \un10_hwres_0\, Q => \LB_ADDR[1]_net_1\);
    
    REG_1_457 : MUX2H
      port map(A => VDB_in_0(2), B => \REG[50]\, S => N_3234_i, Y
         => \REG_1_457\);
    
    \STATE1_ns_0_iv_0_a2[7]\ : NAND2
      port map(A => N_2531, B => \STATE1[3]_net_1\, Y => N_2547);
    
    DS_i_a2 : OR2
      port map(A => DS0B_c, B => DS1B_c, Y => \DS_i_a2\);
    
    un7_ronly_0_a3_0_a2 : AND3FFT
      port map(A => un7_ronly_0_a3_0_a2_1_i, B => N_658, C => 
        \WRITES\, Y => \un7_ronly_0_a3_0_a2\);
    
    STATE5_0_sqmuxa_0_a3_0_a2_1 : NAND2FT
      port map(A => N_2608, B => N_2606_i_i, Y => 
        STATE5_0_sqmuxa_1);
    
    REG_1_477 : MUX2H
      port map(A => VDB_in(22), B => \REG[70]\, S => N_3234_i_0, 
        Y => \REG_1_477\);
    
    \REG_1[89]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_496\, CLR => 
        \un10_hwres_31\, Q => \REG[89]\);
    
    \PIPEB_4_0[30]\ : OR2FT
      port map(A => N_616_0, B => DPR(30), Y => \PIPEB_4[30]\);
    
    REG_1_224 : MUX2H
      port map(A => VDB_in(15), B => \REG[184]\, S => N_2720_i_0, 
        Y => \REG_1_224\);
    
    LB_s_108 : MUX2H
      port map(A => LB_in(29), B => \LB_s[29]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_108\);
    
    un1_STATE1_6_i_a2_0_o2 : OR2FT
      port map(A => N_2524, B => \STATE1_0[1]_net_1\, Y => N_83);
    
    REG_1_222 : MUX2H
      port map(A => VDB_in(13), B => \REG[182]\, S => N_2720_i_0, 
        Y => \REG_1_222\);
    
    \VDBi_58[12]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[12]\, B => N_412_i, C => 
        \VDBi_58_0[9]\, Y => \VDBi_58[12]_net_1\);
    
    \PULSE_42_r[10]\ : OA21
      port map(A => FWIMG2LOAD_0_sqmuxa, B => \PULSE[10]\, C => 
        N_2410, Y => \PULSE_42[10]\);
    
    \REGMAP_0[33]\ : DFF
      port map(CLK => CLK_c_c, D => \un114_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_i_i_0[33]\);
    
    \TCNT_10_0_a2[4]\ : AND2
      port map(A => N_2397, B => I_28, Y => \TCNT_10[4]\);
    
    REG_1_336 : MUX2H
      port map(A => VDB_in(26), B => \REG[371]\, S => N_2944_i_0, 
        Y => \REG_1_336\);
    
    WDOG_3_I_30 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \WDOG_i_0_i[4]\, Y => \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    \VDBi_77[5]\ : MUX2H
      port map(A => \VDBi_66[5]_net_1\, B => \VDBi_77_d[5]_net_1\, 
        S => \VDBi_77_s[8]_net_1\, Y => \VDBi_77[5]_net_1\);
    
    un1_NRDMEBi_2_sqmuxa_2_i_a2_0 : NAND2
      port map(A => DTEST_FIFO, B => \STATE2[5]_net_1\, Y => 
        N_2500);
    
    \LB_i[9]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_521\, CLR => 
        HWRES_c_16, Q => \LB_i[9]_net_1\);
    
    LB_i_515 : MUX2H
      port map(A => \LB_i[3]_net_1\, B => \LB_i_6[3]_net_1\, S
         => N_2570, Y => \LB_i_515\);
    
    \VDBi_16_r[13]\ : OA21TTF
      port map(A => N_2493_i, B => N_2492_i, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[13]\);
    
    REG_1_230 : MUX2H
      port map(A => VDB_in(5), B => \REG[190]\, S => N_2752_i, Y
         => \REG_1_230\);
    
    PIPEA_606 : MUX2H
      port map(A => \PIPEA_7[17]\, B => \PIPEA[17]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_606\);
    
    \RAMAD_VME[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \RAMAD_VME_12\, CLR => 
        \un10_hwres_5\, Q => \RAMAD_VME[8]_net_1\);
    
    \VDBi_16_1_a2_0[3]\ : AND2
      port map(A => N_2511, B => REG_34, Y => N_2467_i);
    
    REG_0_sqmuxa_0_a3_0 : NOR2FT
      port map(A => \REGMAP_0[16]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => REG_0_sqmuxa_0);
    
    un10_hwres_26 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_26\);
    
    REG_1_452 : MUX2H
      port map(A => VDB_in(29), B => \REG[511]\, S => N_3170_i_0, 
        Y => \REG_1_452\);
    
    \WDOG[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \WDOG_3[5]\, CLR => 
        un15_hwres_i, Q => \WDOG[5]_net_1\);
    
    \LB_i_6_0[4]\ : MUX2H
      port map(A => OR_RADDR(2), B => \LB_ADDR[4]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2174);
    
    \REG_1_m[233]\ : AND2
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[233]\, Y => 
        \REG_1_m_i[233]\);
    
    REG_1_472 : MUX2H
      port map(A => VDB_in(17), B => \REG[65]\, S => N_3234_i_1, 
        Y => \REG_1_472\);
    
    \REG_1[501]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_442\, CLR => 
        \un10_hwres_27\, Q => \REG[501]\);
    
    \REG_1[418]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_383\, SET => 
        \un10_hwres_22\, Q => \REG[418]\);
    
    \VDBi_92_0_iv_0_0_4[21]\ : AO21TTF
      port map(A => N_790, B => \REG[69]\, C => N_589, Y => 
        \VDBi_92_0_iv_0_0_4_i[21]\);
    
    \VDBm_0[29]\ : MUX2H
      port map(A => \PIPEB[29]_net_1\, B => \PIPEA[29]_net_1\, S
         => \BLTCYC_1\, Y => N_2325);
    
    un114_reg_ads_0_a3_0_a2 : AND2
      port map(A => N_690, B => un120_reg_ads_1, Y => 
        \un114_reg_ads_0_a3_0_a2\);
    
    SINGCYC_2 : DFFC
      port map(CLK => CLK_c_c, D => \SINGCYC_147\, CLR => 
        HWRES_c_21_0, Q => \SINGCYC_2\);
    
    \LB_i_6[2]\ : MUX2H
      port map(A => N_2172, B => N_2184, S => LB_i_6_sn_N_2, Y
         => N_2218);
    
    SELGEO : LD
      port map(EN => ASB_c, D => \un4_asb_NE\, Q => \TST_c[4]\);
    
    \REGMAP_0[28]\ : DFF
      port map(CLK => CLK_c_c, D => \un102_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[28]_net_1\);
    
    \VDBi_16_1_a2[12]\ : AND2
      port map(A => N_2511_0, B => REG_43, Y => N_2490_i);
    
    \REG_1[79]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_486\, CLR => 
        \un10_hwres_30\, Q => \REG[79]\);
    
    \VDBi_55[17]\ : NOR2
      port map(A => \REGMAP[26]_net_1\, B => \VDBi_23[17]_net_1\, 
        Y => \VDBi_55[17]_net_1\);
    
    MBLTCYC_78 : MUX2H
      port map(A => \MBLTCYC\, B => \TST_c_i_0[0]\, S => N_2385, 
        Y => \MBLTCYC_78\);
    
    REG_1_340 : MUX2H
      port map(A => VDB_in(30), B => \REG[375]\, S => N_2944_i_0, 
        Y => \REG_1_340\);
    
    \REGMAP[13]\ : DFF
      port map(CLK => CLK_c_c, D => \un84_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[13]_net_1\);
    
    \VDBi_23_d[5]\ : MUX2H
      port map(A => \REG[53]\, B => \REG[487]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23_d[5]_net_1\);
    
    PIPEA1_568 : MUX2H
      port map(A => N_264, B => \PIPEA1[12]_net_1\, S => 
        un1_STATE2_13_4_1, Y => \PIPEA1_568\);
    
    PIPEB_48 : MUX2H
      port map(A => \PIPEB_i_i[28]\, B => \PIPEB_4[28]\, S => 
        N_1996_3, Y => \PIPEB_48\);
    
    \VDBi_16_r[10]\ : OA21TTF
      port map(A => N_2487_i, B => N_2486_i, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[10]\);
    
    \VDBi_71[2]\ : MUX2H
      port map(A => \VDBi_60[2]_net_1\, B => \VDBi_71_d[2]_net_1\, 
        S => \VDBi_71_s[4]_net_1\, Y => \VDBi_71[2]_net_1\);
    
    \REG_1[364]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_329\, CLR => 
        \un10_hwres_17\, Q => \REG[364]\);
    
    \VDBi_71[28]\ : MUX2H
      port map(A => \VDBi_60[28]_net_1\, B => \REG[437]\, S => 
        \REGMAP_0[31]_net_1\, Y => \VDBi_71[28]_net_1\);
    
    \REG_1_m[168]\ : NAND2
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[168]\, Y => 
        \REG_1_m[168]_net_1\);
    
    REG_1_454_e_1 : OR2FT
      port map(A => \REGMAP_0[13]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => N_3170_i_1);
    
    \PIPEA1_9_i[9]\ : AND2
      port map(A => DPR(9), B => N_85_4, Y => N_258);
    
    REG_1_398 : MUX2H
      port map(A => VDB_in(24), B => \REG[433]\, S => N_3072_i_0, 
        Y => \REG_1_398\);
    
    \VDBi_92_0_iv_0[26]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[26]_net_1\, C
         => \PIPEA_m[26]_net_1\, Y => \VDBi_92_0_iv_0[26]_net_1\);
    
    \VDBm_0[17]\ : MUX2H
      port map(A => \PIPEB[17]_net_1\, B => \PIPEA[17]_net_1\, S
         => \BLTCYC_2\, Y => N_2313);
    
    \VDBi_92_0_iv_0_0[12]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[12]_net_1\, C
         => N_599, Y => \VDBi_92_0_iv_0_0[12]_net_1\);
    
    LB_i_528 : MUX2H
      port map(A => \LB_i[16]_net_1\, B => \LB_i_6[16]\, S => 
        N_2570_1, Y => \LB_i_528\);
    
    \PIPEA_m[13]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[13]_net_1\, Y => 
        \PIPEA_m[13]_net_1\);
    
    \LB_i_6_1[15]\ : MUX2H
      port map(A => VDB_in_0(15), B => \LB_DOUT[15]_net_1\, S => 
        \STATE5_2[0]_net_1\, Y => N_2197);
    
    \VDBi_53_0_iv_1[14]\ : AO21TTF
      port map(A => \REGMAP_i_i[23]\, B => \REG[247]\, C => 
        \REG_1_m[199]_net_1\, Y => \VDBi_53_0_iv_1_i[14]\);
    
    un776_regmap_21 : OR3FTT
      port map(A => \un776_regmap_17\, B => \REGMAP_0[16]_net_1\, 
        C => \REGMAP_0[26]_net_1\, Y => un776_regmap_21_i);
    
    PIPEB_29 : MUX2H
      port map(A => \PIPEB[9]_net_1\, B => N_2623, S => N_1996_4, 
        Y => \PIPEB_29\);
    
    \VDBi_66_d[11]\ : MUX2H
      port map(A => SPULSE0_c_c, B => N_2028, S => N_2033_0, Y
         => \VDBi_66_d[11]_net_1\);
    
    LB_s_83 : MUX2H
      port map(A => LB_in(4), B => \LB_s[4]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_83\);
    
    un2_nlbrdy_0_a2_2 : OR3
      port map(A => \LBUSTMO_i_0_i[0]\, B => \LBUSTMO_i_0_i[1]\, 
        C => \LBUSTMO[2]_net_1\, Y => un2_nlbrdy_0_a2_2_i);
    
    LB_i_524 : MUX2H
      port map(A => \LB_i[12]_net_1\, B => \LB_i_6[12]\, S => 
        N_2570_1, Y => \LB_i_524\);
    
    \STATE1_ns_0_0[0]\ : OA21FTT
      port map(A => \TST_c[2]\, B => N_2410, C => N_2429, Y => 
        \STATE1_ns_0_0[0]_net_1\);
    
    \REG_1_m[263]\ : NAND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[263]\, Y => 
        \REG_1_m[263]_net_1\);
    
    REG_1_404 : MUX2H
      port map(A => VDB_in(30), B => \REG[439]\, S => N_3072_i_0, 
        Y => \REG_1_404\);
    
    \PIPEA1[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_568\, CLR => CLEAR_21, 
        Q => \PIPEA1[12]_net_1\);
    
    REG_1_480 : MUX2H
      port map(A => VDB_in(25), B => \REG[73]\, S => N_3234_i_0, 
        Y => \REG_1_480\);
    
    \VDBi_53_0_iv_2[1]\ : AO21TTF
      port map(A => \REGMAP[20]_net_1\, B => \REG[186]\, C => 
        \REG_1_m[170]_net_1\, Y => \VDBi_53_0_iv_2_i[1]\);
    
    \LB_DOUT[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_166\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[18]_net_1\);
    
    \REGMAP[8]\ : DFF
      port map(CLK => CLK_c_c, D => \un37_reg_ads_0_a2_4_a2\, Q
         => \TST_c[5]\);
    
    REG_1_215 : MUX2H
      port map(A => VDB_in(6), B => \REG[175]\, S => N_2720_i, Y
         => \REG_1_215\);
    
    \VDBi_23_m[5]\ : AND2
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[5]_net_1\, Y
         => \VDBi_23_m_i[5]\);
    
    \REG_1[398]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_363\, CLR => 
        \un10_hwres_20\, Q => \REG[398]\);
    
    PIPEA_595 : MUX2H
      port map(A => \PIPEA_7[6]\, B => \PIPEA[6]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_595\);
    
    \LBUSTMO[2]\ : DFFS
      port map(CLK => ALICLK_c, D => \LBUSTMO_3[2]\, SET => 
        HWRES_c_13_0, Q => \LBUSTMO[2]_net_1\);
    
    un1_TCNT_1_I_31 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum_0[1]\, B => 
        \DWACT_ADD_CI_0_TMP_1[0]\, Y => I_31_1);
    
    REG_1_385 : MUX2H
      port map(A => VDB_in_0(11), B => \REG[420]\, S => 
        N_3072_i_1, Y => \REG_1_385\);
    
    \REG_1[233]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_246\, SET => 
        \un10_hwres_12\, Q => \REG[233]\);
    
    \PIPEA_7_i_m2[11]\ : MUX2H
      port map(A => DPR(11), B => \PIPEA1[11]_net_1\, S => 
        N_1996_1, Y => N_520);
    
    \REGMAP_0[18]\ : DFF
      port map(CLK => CLK_c_c, D => \un61_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_0[18]_net_1\);
    
    \VDBi_92_iv_0[7]\ : OAI21FTT
      port map(A => N_508, B => \N_2613_0\, C => 
        \VDBi_92_iv_0_2[7]_net_1\, Y => \VDBi_92[7]\);
    
    \PIPEB_4_i[16]\ : AND2
      port map(A => DPR(16), B => N_616_1, Y => N_186);
    
    \STATE2[5]\ : DFFS
      port map(CLK => CLK_c_c, D => \STATE2_ns[0]\, SET => CLEAR, 
        Q => \STATE2[5]_net_1\);
    
    \STATE1[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[1]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1[9]_net_1\);
    
    \VDBi[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_646\, CLR => 
        \un10_hwres_35\, Q => \VDBi[25]_net_1\);
    
    \REGMAP[10]\ : DFF
      port map(CLK => CLK_c_c, D => \un43_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[10]_net_1\);
    
    \REG_1[87]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_494\, CLR => 
        \un10_hwres_31\, Q => \REG[87]\);
    
    LB_i_519 : MUX2H
      port map(A => \LB_i[7]_net_1\, B => \LB_i_6[7]_net_1\, S
         => N_2570, Y => \LB_i_519\);
    
    \VDBi_53_0_iv_0[14]\ : AO21TTF
      port map(A => \REGMAP[12]_net_1\, B => REG_118, C => 
        \REG_1_m[263]_net_1\, Y => \VDBi_53_0_iv_0_i[14]\);
    
    PIPEB_40 : MUX2H
      port map(A => \PIPEB[20]_net_1\, B => N_2632, S => N_1996_3, 
        Y => \PIPEB_40\);
    
    \LB_s[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_79\, CLR => HWRES_c_17, 
        Q => \LB_s[0]_net_1\);
    
    \VDBi_58[11]\ : OA21
      port map(A => \VDBi_53_0_iv_5_i[11]\, B => 
        \VDBi_23_m_i[11]\, C => \VDBi_58_0[9]\, Y => 
        \VDBi_58[11]_net_1\);
    
    \OR_RDATA[5]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_187\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[5]_net_1\);
    
    \REG_1[237]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_250\, SET => 
        \un10_hwres_13\, Q => \REG[237]\);
    
    \VDBi_60[22]\ : MUX2H
      port map(A => \VDBi_55[22]_net_1\, B => LBSP_in_22, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[22]_net_1\);
    
    \VDBi_18[11]\ : MUX2H
      port map(A => \VDBi_16[11]\, B => \REG[59]\, S => 
        \TST_c[5]\, Y => \VDBi_18[11]_net_1\);
    
    REG_1_211 : MUX2H
      port map(A => VDB_in(2), B => \REG[171]\, S => N_2720_i, Y
         => \REG_1_211\);
    
    \STATE5_ns_0_0_0[1]\ : AO21TTF
      port map(A => N_2607, B => \OR_RREQ_sync\, C => N_2597, Y
         => \STATE5_ns_0_0_0_i[1]\);
    
    \REG_1[370]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_335\, CLR => 
        \un10_hwres_18\, Q => \REG[370]\);
    
    \VDBi_66[14]\ : MUX2H
      port map(A => \VDBi_60[14]_net_1\, B => N_2031, S => 
        N_2033_0, Y => \VDBi_66[14]_net_1\);
    
    MYBERRi : DFFS
      port map(CLK => CLK_c_c, D => \MYBERRi_19\, SET => 
        \un10_hwres_4\, Q => \MYBERR_c\);
    
    \VDBi_53_0_iv_5[11]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[11]\, B => 
        \VDBi_53_0_iv_0_i[11]\, C => \VDBi_53_0_iv_1_i[11]\, Y
         => \VDBi_53_0_iv_5_i[11]\);
    
    \REGMAP[1]\ : DFF
      port map(CLK => CLK_c_c, D => \un10_reg_ads_0_a2_1_a2\, Q
         => \REGMAP[1]_net_1\);
    
    PIPEA_592 : MUX2H
      port map(A => \PIPEA_7[3]\, B => \PIPEA[3]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_592\);
    
    un10_hwres_20 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_1, Y => 
        \un10_hwres_20\);
    
    un10_hwres_32 : OR2
      port map(A => HWRES_c_0_3, B => WDOGTO_0, Y => 
        \un10_hwres_32\);
    
    \VDBi_53_0_iv_3[11]\ : AO21TTF
      port map(A => \REGMAP_0[16]_net_1\, B => \REG[132]\, C => 
        \VDBi_53_0_iv_2[11]_net_1\, Y => \VDBi_53_0_iv_3_i[11]\);
    
    \REG_1[127]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_135\, CLR => 
        \un10_hwres_8\, Q => REG_126);
    
    \REGMAP[5]\ : DFF
      port map(CLK => CLK_c_c, D => \un25_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[5]_net_1\);
    
    un6_cycs_i_a2 : NOR2
      port map(A => \CYCS\, B => \TST_c[0]\, Y => N_2421);
    
    \REG_1[456]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_421\, CLR => 
        \un10_hwres_25\, Q => \REG[456]\);
    
    \LB_s[6]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_85\, CLR => HWRES_c_19, 
        Q => \LB_s[6]_net_1\);
    
    \VDBi_53_0_iv_1[10]\ : AO21TTF
      port map(A => \REGMAP_i_i[23]\, B => \REG[243]\, C => 
        \REG_1_m[195]_net_1\, Y => \VDBi_53_0_iv_1_i[10]\);
    
    \PIPEA[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_600\, CLR => CLEAR_23, 
        Q => \PIPEA[11]_net_1\);
    
    \VDBi_92_iv[3]\ : OAI21FTT
      port map(A => \VDBi_80[3]_net_1\, B => \N_2613_0\, C => 
        \VDBi_92_iv_2[3]_net_1\, Y => \VDBi_92[3]\);
    
    \VDBi_71[11]\ : MUX2H
      port map(A => \VDBi_66[11]_net_1\, B => \REG[420]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71[11]_net_1\);
    
    \PIPEA1_9_i[21]\ : AND2
      port map(A => DPR(21), B => N_85_3, Y => N_282);
    
    OR_RREQ_sync : DFFC
      port map(CLK => ALICLK_c, D => OR_RREQ, CLR => HWRES_c_20, 
        Q => \OR_RREQ_sync\);
    
    \VDBm_0_i_m2[11]\ : MUX2H
      port map(A => \PIPEB[11]_net_1\, B => \PIPEA[11]_net_1\, S
         => \BLTCYC_0\, Y => N_2540);
    
    \LB_DOUT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_150\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[2]_net_1\);
    
    \VDBm[7]\ : MUX2H
      port map(A => N_2303, B => \VDBi[7]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_7);
    
    \REG_88[88]\ : NOR2FT
      port map(A => N_2159, B => N_2566, Y => \REG_88[88]_net_1\);
    
    \VDBi_92_0_iv_1[17]\ : AOI21TTF
      port map(A => \LB_s[17]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[17]_net_1\, Y => 
        \VDBi_92_0_iv_1[17]_net_1\);
    
    \REG_1[408]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_373\, CLR => 
        \un10_hwres_21\, Q => \REG[408]\);
    
    \VADm[24]\ : AND2FT
      port map(A => N_2507_1, B => \PIPEA[24]_net_1\, Y => 
        VADm(24));
    
    EFS : DFFS
      port map(CLK => CLK_c_c, D => EF, SET => CLEAR_20, Q => 
        \EFS\);
    
    un1_NRDMEBi_2_sqmuxa_1_i_a3_i_o2_i_a2 : OR2FT
      port map(A => \STATE2[5]_net_1\, B => \REG[5]\, Y => N_584);
    
    \REG_i[400]\ : INV
      port map(A => \REG[400]\, Y => REG_i_0_395);
    
    \RAMDTS[6]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(6), CLR => HWRES_c_21, 
        Q => \RAMDTS[6]_net_1\);
    
    \VDBi_16_1_a3_2[0]\ : NAND3
      port map(A => N_2380_1, B => \VDBi_16_1_a3_2_0[0]_net_1\, C
         => \REGMAP[1]_net_1\, Y => N_2380);
    
    REG_1_334 : MUX2H
      port map(A => VDB_in(24), B => \REG[369]\, S => N_2944_i_0, 
        Y => \REG_1_334\);
    
    \REG_1[441]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_406\, CLR => 
        \un10_hwres_24\, Q => \REG[441]\);
    
    un1_TCNT_1_I_20 : XOR2
      port map(A => \TCNT[1]_net_1\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[1]\);
    
    un1_vas7_i_o2 : NOR2FT
      port map(A => \CYCS\, B => \CYCS1\, Y => N_2403);
    
    \PIPEA1[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_559\, CLR => CLEAR_22, 
        Q => \PIPEA1[3]_net_1\);
    
    \VDBi_77_0[0]\ : MUX2H
      port map(A => REG_456, B => \REG[441]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_2052);
    
    REG_1_198 : MUX2H
      port map(A => VDB_in(5), B => \REG[158]\, S => N_2688_i, Y
         => \REG_1_198\);
    
    \PIPEA_7_i_m2[29]\ : MUX2H
      port map(A => DPR(29), B => \PIPEA1[29]_net_1\, S => 
        N_1996_0, Y => N_538);
    
    \REG_1[77]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_484\, CLR => 
        \un10_hwres_30\, Q => \REG[77]\);
    
    PIPEB_45 : MUX2H
      port map(A => \PIPEB[25]_net_1\, B => N_229, S => N_1996_3, 
        Y => \PIPEB_45\);
    
    N_77_i_i_o2 : NOR3
      port map(A => N_449, B => N_440, C => N_77_i_i_o2_1_i, Y
         => N_472_i_0);
    
    \LB_i_6_0[8]\ : OR2FT
      port map(A => \STATE5_0[0]_net_1\, B => \LB_ADDR[8]_net_1\, 
        Y => N_2178);
    
    \REG_1[165]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_205\, CLR => 
        \un10_hwres_9\, Q => \REG[165]\);
    
    \PIPEB_4_i[19]\ : AND2
      port map(A => DPR(19), B => N_616_1, Y => N_2631);
    
    \REG_1_0[127]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_135\, CLR => 
        \un10_hwres_8_0\, Q => \REG_0[127]\);
    
    REG_1_265 : MUX2H
      port map(A => VDB_in(3), B => \REG[252]\, S => N_2816_i_0, 
        Y => \REG_1_265\);
    
    LB_WRITE_sync : DFFC
      port map(CLK => ALICLK_c, D => \LB_WRITE\, CLR => 
        HWRES_c_14, Q => \LB_WRITE_sync\);
    
    REG_1_341 : MUX2H
      port map(A => VDB_in(31), B => \REG[376]\, S => N_2944_i_0, 
        Y => \REG_1_341\);
    
    REG_1_437 : MUX2H
      port map(A => VDB_in_0(14), B => \REG[496]\, S => 
        N_3170_i_1, Y => \REG_1_437\);
    
    \LB_i_6_0[11]\ : AND2
      port map(A => \LB_ADDR[11]_net_1\, B => \STATE5_2[0]_net_1\, 
        Y => N_2181);
    
    \VDBi_80[3]\ : MUX2H
      port map(A => \VDBi_80_d[3]_net_1\, B => \VDBi_60[3]_net_1\, 
        S => \VDBi_80_s[3]_net_1\, Y => \VDBi_80[3]_net_1\);
    
    \PIPEB[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_29\, CLR => CLEAR_28, 
        Q => \PIPEB[9]_net_1\);
    
    \REG_1[200]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_240\, CLR => 
        \un10_hwres_12\, Q => \REG[200]\);
    
    \PIPEA_7_r[7]\ : AND2
      port map(A => N_85_2, B => N_516, Y => \PIPEA_7[7]\);
    
    \VADm[31]\ : NOR2FT
      port map(A => \PIPEA[31]_net_1\, B => N_2507_1, Y => 
        VADm(31));
    
    \VDBi_92_iv_0_m2[7]\ : MUX2H
      port map(A => N_476, B => REG_479, S => \REGMAP[35]_net_1\, 
        Y => N_508);
    
    \VDBi_53_0_iv_0[10]\ : AO21TTF
      port map(A => \REGMAP[12]_net_1\, B => REG_114, C => 
        \REG_1_m[259]_net_1\, Y => \VDBi_53_0_iv_0_i[10]\);
    
    \VDBi_71_i_m2_d[7]\ : MUX2H
      port map(A => N_2024, B => \REG[416]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71_i_m2_d[7]_net_1\);
    
    \VDBi_92_0_iv_1[28]\ : AOI21TTF
      port map(A => \LB_s[28]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[28]_net_1\, Y => 
        \VDBi_92_0_iv_1[28]_net_1\);
    
    \REG_1[507]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_448\, CLR => 
        \un10_hwres_27\, Q => \REG[507]\);
    
    un1_EVREAD_DS_1_sqmuxa_1_0_a2_0_0_o2 : NAND2
      port map(A => \STATE2[1]_net_1\, B => \TST_c[2]\, Y => 
        N_426);
    
    \VDBi[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_638\, CLR => 
        \un10_hwres_34\, Q => \VDBi[17]_net_1\);
    
    \REG_88[84]\ : NOR2FT
      port map(A => N_2155, B => N_2566, Y => \REG_88[84]_net_1\);
    
    \REG_1[198]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_238\, CLR => 
        \un10_hwres_12\, Q => \REG[198]\);
    
    \LB_i_6_r[22]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_0, C => N_2204, 
        Y => \LB_i_6[22]\);
    
    \VDBi_92_0_iv_0_0[25]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[25]_net_1\, C
         => N_603, Y => \VDBi_92_0_iv_0_0[25]_net_1\);
    
    \VDBi_92_iv[2]\ : OAI21FTT
      port map(A => \VDBi_80[2]_net_1\, B => \N_2613_0\, C => 
        \VDBi_92_iv_2[2]_net_1\, Y => \VDBi_92[2]\);
    
    \PIPEA_7_i_m2[24]\ : MUX2H
      port map(A => DPR(24), B => \PIPEA1[24]_net_1\, S => 
        N_1996_0, Y => N_533);
    
    \LB_i_6_r[19]\ : AND3
      port map(A => N_2572_1, B => LB_i_6_sn_N_2_1, C => N_2201, 
        Y => \LB_i_6[19]\);
    
    REG_1_423 : MUX2H
      port map(A => VDB_in_0(0), B => \REG[482]\, S => N_3170_i, 
        Y => \REG_1_423\);
    
    LB_s_107 : MUX2H
      port map(A => LB_in(28), B => \LB_s[28]_net_1\, S => 
        STATE5_0_sqmuxa_0, Y => \LB_s_107\);
    
    REG_1_261 : MUX2H
      port map(A => VDB_in(15), B => \REG[248]\, S => N_2784_i_0, 
        Y => \REG_1_261\);
    
    \LB_i_6_1[30]\ : MUX2H
      port map(A => VDB_in(30), B => \LB_DOUT[30]_net_1\, S => 
        \STATE5_0[0]_net_1\, Y => N_2212);
    
    STATE1_tr27_i_o4_0 : OAI21
      port map(A => \REGMAP[36]_net_1\, B => \REGMAP[10]_net_1\, 
        C => N_425, Y => N_2533);
    
    \LB_DOUT[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_175\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[27]_net_1\);
    
    un1_vas7_i : OAI21FTF
      port map(A => \STATE1[5]_net_1\, B => N_2403, C => N_2385, 
        Y => N_59);
    
    REG_1_299 : MUX2H
      port map(A => VDB_in(21), B => \REG[286]\, S => N_2880_i, Y
         => \REG_1_299\);
    
    \VDBi_16_1_a2[9]\ : AND2
      port map(A => N_2511_0, B => REG_40, Y => N_2484_i);
    
    REG_1_432 : MUX2H
      port map(A => VDB_in_0(9), B => \REG[491]\, S => N_3170_i, 
        Y => \REG_1_432\);
    
    \REG_1[425]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_390\, CLR => 
        \un10_hwres_22\, Q => \REG[425]\);
    
    \STATE1_ns_0_iv_0_a2_0[8]\ : OR3
      port map(A => N_2552_1, B => N_1898, C => N_2550_1, Y => 
        N_2550);
    
    \REG_1[417]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_382\, SET => 
        \un10_hwres_22\, Q => \REG[417]\);
    
    \OR_RDATA_5_i[4]\ : AND2
      port map(A => N_2572, B => LB_in(4), Y => N_2567);
    
    \PIPEB[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_41\, CLR => CLEAR_27, 
        Q => \PIPEB[21]_net_1\);
    
    REG1_0_sqmuxa_0_a3 : NOR2FT
      port map(A => \REGMAP[1]_net_1\, B => PULSE_0_sqmuxa_1_2, Y
         => REG1_0_sqmuxa);
    
    \PIPEA_7_r[12]\ : AND2
      port map(A => N_85_2, B => N_521, Y => \PIPEA_7[12]\);
    
    \PIPEA1[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_562\, CLR => CLEAR_23, 
        Q => \PIPEA1[6]_net_1\);
    
    PIPEB_37 : MUX2H
      port map(A => \PIPEB[17]_net_1\, B => N_2630, S => N_1996_4, 
        Y => \PIPEB_37\);
    
    VAS_56 : MUX2H
      port map(A => \VAS[5]_net_1\, B => VAD_in_4, S => 
        \TST_c[1]\, Y => \VAS_56\);
    
    \REG_1[187]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_227\, CLR => 
        \un10_hwres_11\, Q => \REG[187]\);
    
    \PIPEA[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_608\, CLR => CLEAR_24, 
        Q => \PIPEA[19]_net_1\);
    
    un1_REG_0_sqmuxa_i_a2_0 : NOR3
      port map(A => \STATE5[2]_net_1\, B => \OR_RREQ_sync\, C => 
        \LB_REQ_sync\, Y => N_2577_i);
    
    VDBi_636 : MUX2H
      port map(A => \VDBi_92[15]\, B => \VDBi[15]_net_1\, S => 
        un1_STATE1_34_1, Y => \VDBi_636\);
    
    \VDBi_92_0_iv_1[14]\ : AOI21TTF
      port map(A => \LB_s[14]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[14]_net_1\, Y => 
        \VDBi_92_0_iv_1[14]_net_1\);
    
    \PIPEA[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_589\, CLR => CLEAR_23, 
        Q => \PIPEA[0]_net_1\);
    
    LB_DOUT_167 : MUX2H
      port map(A => VDB_in(19), B => \LB_DOUT[19]_net_1\, S => 
        LB_DOUT_0_sqmuxa_1, Y => \LB_DOUT_167\);
    
    LB_s_94 : MUX2H
      port map(A => LB_in(15), B => \LB_s[15]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_94\);
    
    \REG_1[429]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_394\, CLR => 
        \un10_hwres_23\, Q => \REG[429]\);
    
    PIPEA1_578 : MUX2H
      port map(A => N_284, B => \PIPEA1[22]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_578\);
    
    \VDBi_53_0_iv_3[9]\ : AO21TTF
      port map(A => \REGMAP[16]_net_1\, B => \REG[130]\, C => 
        \VDBi_53_0_iv_2[9]_net_1\, Y => \VDBi_53_0_iv_3_i[9]\);
    
    REG_1_450 : MUX2H
      port map(A => VDB_in(27), B => \REG[509]\, S => N_3170_i_0, 
        Y => \REG_1_450\);
    
    \VDBi_16_1_a2_0[13]\ : AND2
      port map(A => N_2512_0, B => \REG[13]\, Y => N_2493_i);
    
    un10_hwres_3 : OR2
      port map(A => HWRES_c_0_6, B => \WDOGTO\, Y => 
        \un10_hwres_3\);
    
    REG_1_329 : MUX2H
      port map(A => VDB_in(19), B => \REG[364]\, S => N_2944_i, Y
         => \REG_1_329\);
    
    \REG_1[154]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_194\, CLR => 
        \un10_hwres_9\, Q => \REG[154]\);
    
    LB_DOUT_0_sqmuxa_0_a2_0_a2 : OR2FT
      port map(A => \REGMAP[36]_net_1\, B => PULSE_0_sqmuxa_1_2, 
        Y => LB_DOUT_0_sqmuxa);
    
    un81_reg_ads_0_a3_0_a2_0 : OR2FT
      port map(A => N_463, B => \VAS[1]_net_1\, Y => N_716);
    
    \VDBi_77_0[5]\ : MUX2H
      port map(A => REG_461, B => \REG[446]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_2057);
    
    REG_1_470 : MUX2H
      port map(A => VDB_in_0(15), B => \REG[63]\, S => N_3234_i_1, 
        Y => \REG_1_470\);
    
    \VDBi_77_0[6]\ : MUX2H
      port map(A => REG_462, B => \REG[447]\, S => 
        \REGMAP_i_i_0[33]\, Y => N_2058);
    
    un10_hwres_33 : OR2
      port map(A => HWRES_c_0_3, B => WDOGTO_0, Y => 
        \un10_hwres_33\);
    
    REG_1_355 : MUX2H
      port map(A => VDB_in_0(13), B => \REG[390]\, S => 
        N_2976_i_0, Y => \REG_1_355\);
    
    \REG_1[438]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_403\, CLR => 
        \un10_hwres_23\, Q => \REG[438]\);
    
    \REG_1_m[169]\ : NAND2
      port map(A => \REGMAP[19]_net_1\, B => \REG[169]\, Y => 
        \REG_1_m[169]_net_1\);
    
    \VDBi_23_d[14]\ : MUX2H
      port map(A => \REG[62]\, B => \REG[496]\, S => 
        \REGMAP_1[13]_net_1\, Y => \VDBi_23_d[14]_net_1\);
    
    \PIPEA1_9_i[13]\ : AND2
      port map(A => DPR(13), B => N_85_4, Y => N_266);
    
    \VDBi[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_643\, CLR => 
        \un10_hwres_34\, Q => \VDBi[22]_net_1\);
    
    \REG_1[412]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_377\, CLR => 
        \un10_hwres_21\, Q => \REG[412]\);
    
    REG_1_375 : MUX2H
      port map(A => VDB_in_0(1), B => \REG[410]\, S => N_3072_i, 
        Y => \REG_1_375\);
    
    un7_noe32ri_0_0_0 : OAI21FTF
      port map(A => \un7_noe32ri_0_0_a2_0\, B => \LWORDS\, C => 
        \NOEAD_c_0_0\, Y => un7_noe32ri_0);
    
    \REG_1[156]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_196\, CLR => 
        \un10_hwres_9\, Q => \REG[156]\);
    
    \VDBi_60_d[8]\ : MUX2H
      port map(A => LBSP_c(2), B => L2R_c_c, S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60_d[8]_net_1\);
    
    \VDBi_92_0_iv_1[9]\ : AOI21TTF
      port map(A => \LB_s[9]_net_1\, B => N_7_i, C => 
        \VDBi_92_0_iv_0[9]_net_1\, Y => \VDBi_92_0_iv_1[9]_net_1\);
    
    OR_RACK_1_sqmuxa_i_i_a2 : AND2
      port map(A => N_2597_1, B => \STATE5[2]_net_1\, Y => 
        \OR_RACK_1_sqmuxa_i_i_a2\);
    
    \REG_1[371]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_336\, CLR => 
        \un10_hwres_18\, Q => \REG[371]\);
    
    \PIPEA_7_r[2]\ : AND2
      port map(A => N_85_3, B => N_511, Y => \PIPEA_7[2]\);
    
    \VDBi_60_d[2]\ : MUX2H
      port map(A => L1R_c_c, B => LBSP_c(2), S => 
        \REGMAP[28]_net_1\, Y => \VDBi_60_d[2]_net_1\);
    
    \LBUSTMO_3_0[2]\ : OR2FT
      port map(A => N_2572_0, B => I_20_3, Y => \LBUSTMO_3[2]\);
    
    REG_1_310 : MUX2H
      port map(A => VDB_in_0(0), B => \REG[345]\, S => N_2944_i, 
        Y => \REG_1_310\);
    
    \PIPEB[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_23\, CLR => CLEAR_28, 
        Q => \PIPEB[3]_net_1\);
    
    \VDBi_60[23]\ : MUX2H
      port map(A => \VDBi_55[23]_net_1\, B => LBSP_in_23, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[23]_net_1\);
    
    \TCNT_10_r[7]\ : OA21FTT
      port map(A => \N_1897\, B => I_34_1, C => N_2523_0, Y => 
        \TCNT_10[7]\);
    
    \LB_i_6_0[6]\ : MUX2H
      port map(A => OR_RADDR(4), B => \LB_ADDR[6]_net_1\, S => 
        \STATE5_3[0]_net_1\, Y => N_2176);
    
    \VDBi_53_0_iv_5[4]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[4]\, B => 
        \VDBi_53_0_iv_0_i[4]\, C => \VDBi_53_0_iv_1_i[4]\, Y => 
        \VDBi_53_0_iv_5_i[4]\);
    
    REG_1_135 : MUX2H
      port map(A => \REG_0[127]\, B => VDB_in(6), S => 
        REG_0_sqmuxa, Y => \REG_1_135\);
    
    LB_i_518 : MUX2H
      port map(A => \LB_i[6]_net_1\, B => \LB_i_6[6]_net_1\, S
         => N_2570, Y => \LB_i_518\);
    
    \PIPEB[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_25\, CLR => CLEAR_28, 
        Q => \PIPEB[5]_net_1\);
    
    \VDBi_55[8]\ : OA21TTF
      port map(A => \VDBi_23_m_i[8]\, B => \VDBi_53_0_iv_6_i[8]\, 
        C => \REGMAP[26]_net_1\, Y => \VDBi_55[8]_net_1\);
    
    N_2522_i_i_o2_1 : AND3
      port map(A => N_425, B => \STATE1_0[9]_net_1\, C => 
        \REGMAP[0]_net_1\, Y => N_457_i_0_1);
    
    un78_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_689_i, B => un43_reg_ads_1, Y => 
        \un78_reg_ads_0_a3_0_a2\);
    
    \VDBi_92_0_iv_1[22]\ : AOI21TTF
      port map(A => \LB_s[22]_net_1\, B => N_7_i_0, C => 
        \VDBi_92_0_iv_0[22]_net_1\, Y => 
        \VDBi_92_0_iv_1[22]_net_1\);
    
    \PIPEA_m[15]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[15]_net_1\, Y => 
        \PIPEA_m[15]_net_1\);
    
    \REG_1_m[250]\ : AND2
      port map(A => \REGMAP[24]_net_1\, B => \REG[250]\, Y => 
        \REG_1_m_i[250]\);
    
    \PULSE_42_f0_i[3]\ : OA21TTF
      port map(A => \PULSE[3]\, B => N_2409, C => 
        \STATE1_0[7]_net_1\, Y => N_2391);
    
    LB_i_514 : MUX2H
      port map(A => \LB_i[2]_net_1\, B => \LB_i_6[2]_net_1\, S
         => N_2570, Y => \LB_i_514\);
    
    \VDBi_18[17]\ : NAND2
      port map(A => \REG[65]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[17]_net_1\);
    
    \VDBi_18[29]\ : NAND2
      port map(A => \REG[77]\, B => \TST_c_0[5]\, Y => 
        \VDBi_18[29]_net_1\);
    
    \FBOUT_m[1]\ : NAND2
      port map(A => FBOUT(1), B => \STATE1[2]_net_1\, Y => 
        \FBOUT_m[1]_net_1\);
    
    un1_TCNT_1_I_15 : XOR2
      port map(A => \TCNT[3]_net_1\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_2_0[0]\);
    
    un13_reg_ads_0_a2_0_a2 : NOR3FTT
      port map(A => \WRITES_0\, B => un13_reg_ads_1, C => N_681_i, 
        Y => \un13_reg_ads_0_a2_0_a2\);
    
    un1_LBUSTMO_1_I_28 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\);
    
    \REG_1[485]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_426\, CLR => 
        \un10_hwres_25\, Q => \REG[485]\);
    
    REG_1_405_e : OR2FT
      port map(A => \REGMAP_0[31]_net_1\, B => PULSE_0_sqmuxa_1, 
        Y => N_3072_i);
    
    \VDBi_92_0_iv[29]\ : OAI21FTT
      port map(A => \VDBi_71[29]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[29]_net_1\, Y => \VDBi_92[29]\);
    
    REG3_113 : MUX2H
      port map(A => \REG_c[0]\, B => VDB_in(0), S => 
        REG1_0_sqmuxa, Y => \REG3_113\);
    
    REG3_128 : MUX2H
      port map(A => \REG[15]\, B => VDB_in(15), S => 
        REG1_0_sqmuxa_0, Y => \REG3_128\);
    
    \PIPEB[29]\ : DFFS
      port map(CLK => CLK_c_c, D => \PIPEB_49\, SET => CLEAR_27, 
        Q => \PIPEB[29]_net_1\);
    
    un1_LBUSTMO_1_I_7 : NOR2FT
      port map(A => \LBUSTMO_i_0_i[3]\, B => N_66_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_3[0]\);
    
    un81_reg_ads_0_a3_0_a2 : NOR2FT
      port map(A => N_675, B => N_716, Y => 
        \un81_reg_ads_0_a3_0_a2\);
    
    REG_1_422_e : NOR2FT
      port map(A => \REGMAP[32]_net_1\, B => PULSE_0_sqmuxa_1_2, 
        Y => FWIMG2LOAD_0_sqmuxa);
    
    \LB_i_6_r[10]\ : AND2
      port map(A => N_2226, B => N_2572_2, Y => 
        \LB_i_6[10]_net_1\);
    
    \VDBi_53_0_iv_1[5]\ : AO21TTF
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[238]\, C => 
        \REG_1_m[190]_net_1\, Y => \VDBi_53_0_iv_1_i[5]\);
    
    VAS_55 : MUX2H
      port map(A => \VAS[4]_net_1\, B => VAD_in_3, S => 
        \TST_c[1]\, Y => \VAS_55\);
    
    REG_1_228 : MUX2H
      port map(A => VDB_in(3), B => \REG[188]\, S => N_2752_i, Y
         => \REG_1_228\);
    
    un2_reg_ads_0_a3_0_a2 : AND3FTT
      port map(A => N_724, B => N_685, C => N_674, Y => 
        \un2_reg_ads_0_a3_0_a2\);
    
    LB_DOUT_149 : MUX2H
      port map(A => VDB_in(1), B => \LB_DOUT[1]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_149\);
    
    \RAMRD\ : DFFS
      port map(CLK => CLK_c_c, D => \TCNT_0_sqmuxa_i_s\, SET => 
        \un10_hwres_5\, Q => RAMRD);
    
    un776_regmap_14_i_0_o2 : OR2
      port map(A => \REGMAP_i_i[33]\, B => \REGMAP[34]_net_1\, Y
         => \N_441\);
    
    REG_1_199 : MUX2H
      port map(A => VDB_in(6), B => \REG[159]\, S => N_2688_i, Y
         => \REG_1_199\);
    
    \VDBm[10]\ : MUX2H
      port map(A => N_2306, B => \VDBi[10]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_10);
    
    un1_TCNT_1_I_27 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[6]\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => I_27);
    
    \VDBi_92_0_iv_0[18]\ : AOI21TTF
      port map(A => \STATE1_1[2]_net_1\, B => \VDBi[18]_net_1\, C
         => \PIPEA_m[18]_net_1\, Y => \VDBi_92_0_iv_0[18]_net_1\);
    
    \PIPEB_4_i[17]\ : AND2
      port map(A => DPR(17), B => N_616_1, Y => N_2630);
    
    \LB_s[17]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_96\, CLR => HWRES_c_17, 
        Q => \LB_s[17]_net_1\);
    
    \REG_1[489]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_430\, CLR => 
        \un10_hwres_26\, Q => \REG[489]\);
    
    un1_STATE5_15_i_a2_0 : AND2FT
      port map(A => \LB_WRITE_sync\, B => N_2607, Y => N_2602_i);
    
    \VDBi_71_d[3]\ : MUX2H
      port map(A => N_2020, B => \REG[412]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71_d[3]_net_1\);
    
    \REG_1[365]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_330\, CLR => 
        \un10_hwres_17\, Q => \REG[365]\);
    
    \VDBi_18[16]\ : NAND2
      port map(A => \REG[64]\, B => \TST_c_1[5]\, Y => 
        \VDBi_18[16]_net_1\);
    
    \LBUSTMO_3_0[0]\ : OR2FT
      port map(A => N_2572_0, B => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, Y => \LBUSTMO_3[0]\);
    
    \VDBi_92_0_iv[23]\ : OAI21FTT
      port map(A => \VDBi_71[23]_net_1\, B => N_2613, C => 
        \VDBi_92_0_iv_1[23]_net_1\, Y => \VDBi_92[23]\);
    
    \STATE5_ns_0_0_a2_0[1]\ : OR2
      port map(A => \STATE5_0[2]_net_1\, B => LB_i_6_sn_N_2_0, Y
         => N_2596);
    
    \LB_i_6_r[4]\ : AND2
      port map(A => N_2220, B => N_2572_3, Y => \LB_i_6[4]_net_1\);
    
    PIPEB_31 : MUX2H
      port map(A => \PIPEB[11]_net_1\, B => N_2625, S => N_1996_4, 
        Y => \PIPEB_31\);
    
    REG_1_360 : MUX2H
      port map(A => VDB_in_0(2), B => \REG[395]\, S => N_3008_i, 
        Y => \REG_1_360\);
    
    \PIPEA_m[17]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[17]_net_1\, Y => 
        \PIPEA_m[17]_net_1\);
    
    \STATE1_ns_0_iv_0_a2[9]\ : AND2
      port map(A => N_2531, B => \STATE1_0[1]_net_1\, Y => 
        N_2551_i);
    
    \REG_1[199]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_239\, CLR => 
        \un10_hwres_12\, Q => \REG[199]\);
    
    \VDBm[20]\ : MUX2H
      port map(A => N_2316, B => \VDBi[20]_net_1\, S => 
        \SINGCYC_1\, Y => VDBm_20);
    
    \REG_1[407]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_372\, CLR => 
        \un10_hwres_21\, Q => \REG[407]\);
    
    \REG_i[397]\ : INV
      port map(A => \REG[397]\, Y => REG_i_0_392);
    
    LB_i_532 : MUX2H
      port map(A => \LB_i[20]_net_1\, B => \LB_i_6[20]\, S => 
        N_2570_1, Y => \LB_i_532\);
    
    \VDBi_18_i_m2[12]\ : MUX2H
      port map(A => \VDBi_16[12]\, B => \REG[60]\, S => 
        \TST_c[5]\, Y => N_497);
    
    un2_vsel_1_i_a2_1_0 : NAND2
      port map(A => IACKB_c, B => \TST_c[4]\, Y => 
        un2_vsel_1_i_a2_1_0_i);
    
    PIPEB_51 : MUX2H
      port map(A => \PIPEB[31]_net_1\, B => N_236, S => N_1996_2, 
        Y => \PIPEB_51\);
    
    \PIPEB[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_21\, CLR => CLEAR_27, 
        Q => \PIPEB[1]_net_1\);
    
    un108_reg_ads_0_a3_0_a2 : NOR2
      port map(A => N_684_i, B => un105_reg_ads_1_0, Y => 
        \un108_reg_ads_0_a3_0_a2\);
    
    \REG_1_m[164]\ : NAND2
      port map(A => \REGMAP_0[18]_net_1\, B => \REG[164]\, Y => 
        \REG_1_m[164]_net_1\);
    
    REG_1_296 : MUX2H
      port map(A => VDB_in(18), B => \REG[283]\, S => N_2880_i, Y
         => \REG_1_296\);
    
    \OR_RDATA_5_i_o2_0[0]\ : OR2
      port map(A => N_66_0, B => \STATE5_0[2]_net_1\, Y => 
        N_2572_0);
    
    \VDBi_58[6]\ : MUX2H
      port map(A => \VDBi_55[6]_net_1\, B => REG_334, S => 
        \REGMAP[27]_net_1\, Y => \VDBi_58[6]_net_1\);
    
    \VDBi_71_d_0[1]\ : MUX2H
      port map(A => L1A_c_c, B => \VDBi_71_d[1]_net_1\, S => 
        \VDBi_71_s[1]_net_1\, Y => \VDBi_71_d_0[1]_net_1\);
    
    \STATE1_ns_0_iv_0_0[1]\ : NAND3FTT
      port map(A => \STATE1_ns_0_iv_0_0_0_i[1]\, B => N_627, C
         => N_2431, Y => \STATE1_ns[1]\);
    
    REG_1_343 : MUX2H
      port map(A => VDB_in_0(1), B => \REG[378]\, S => N_2976_i, 
        Y => \REG_1_343\);
    
    \VDBi_16_1_a2_1[3]\ : NAND2
      port map(A => N_2512, B => \REG[3]\, Y => N_2468);
    
    \VDBi_92_0_iv_0_a2_8[21]\ : NOR2FT
      port map(A => \REGMAP_0[31]_net_1\, B => \N_2613_0\, Y => 
        N_723);
    
    \STATE2_ns_o2_0_0[0]\ : OR2FT
      port map(A => N_1756_1, B => \REG[5]\, Y => N_1756);
    
    \VDBi_16_r[12]\ : OA21TTF
      port map(A => N_2491_i, B => N_2490_i, C => 
        \REGMAP[7]_net_1\, Y => \VDBi_16[12]\);
    
    un120_reg_ads_0_a3_0_a2_1 : NOR2FT
      port map(A => N_674, B => N_672, Y => un120_reg_ads_1);
    
    \PIPEA_m[8]\ : NAND2
      port map(A => N_457_i_0, B => \PIPEA[8]_net_1\, Y => 
        \PIPEA_m[8]_net_1\);
    
    LB_DOUT_155 : MUX2H
      port map(A => VDB_in(7), B => \LB_DOUT[7]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_155\);
    
    \VDBm_0[22]\ : MUX2H
      port map(A => \PIPEB[22]_net_1\, B => \PIPEA[22]_net_1\, S
         => \BLTCYC_1\, Y => N_2318);
    
    \VDBi_53_0_iv_5[15]\ : OR3
      port map(A => \VDBi_53_0_iv_3_i[15]\, B => 
        \VDBi_53_0_iv_0_i[15]\, C => \VDBi_53_0_iv_1_i[15]\, Y
         => \VDBi_53_0_iv_5_i[15]\);
    
    \REG_1[402]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_367\, CLR => 
        \un10_hwres_20\, Q => \REG[402]\);
    
    \STATE1_i[8]\ : INV
      port map(A => \STATE1[8]_net_1\, Y => \STATE1_i_0[8]\);
    
    \STATE5_ns_0_0[0]\ : NAND3FTT
      port map(A => \STATE5_ns_0_0_0_i[0]\, B => 
        STATE5_0_sqmuxa_0, C => N_2596, Y => \STATE5_ns[0]\);
    
    \LBUSTMO[4]\ : DFFS
      port map(CLK => ALICLK_c, D => \LBUSTMO_3[4]\, SET => 
        HWRES_c_14, Q => \LBUSTMO[4]_net_1\);
    
    \VDBi_16_1_0[7]\ : AO21TTF
      port map(A => \REGMAP[2]_net_1\, B => REG_c_23, C => N_2480, 
        Y => \VDBi_16_1_0_i[7]\);
    
    un1_LBUSTMO_1_I_26 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0[0]\, B => 
        \DWACT_ADD_CI_0_TMP_0[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\);
    
    \VDBi_53_0_iv_3[15]\ : AO21TTF
      port map(A => \REGMAP_0[16]_net_1\, B => \REG[136]\, C => 
        \VDBi_53_0_iv_2[15]_net_1\, Y => \VDBi_53_0_iv_3_i[15]\);
    
    \REG_1[296]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_309\, CLR => 
        \un10_hwres_17\, Q => \REG[296]\);
    
    \VDBi_92_0_iv[14]\ : OAI21FTT
      port map(A => \VDBi_77[14]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[14]_net_1\, Y => \VDBi_92[14]\);
    
    \LB_DOUT[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_161\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[13]_net_1\);
    
    un10_hwres_6 : OR2
      port map(A => HWRES_c_0_6, B => WDOGTO_2, Y => 
        \un10_hwres_6\);
    
    REG1_0_sqmuxa_1_0_a3 : OR2FT
      port map(A => \REGMAP[14]_net_1\, B => PULSE_0_sqmuxa_1_2, 
        Y => REG1_0_sqmuxa_1);
    
    N_7_i_0_a2_1 : NOR2FT
      port map(A => \STATE1_0[9]_net_1\, B => N_425, Y => N_7_i_1);
    
    \VDBi_53_0_iv_2[4]\ : AOI21TTF
      port map(A => \REGMAP[19]_net_1\, B => \REG[173]\, C => 
        \REG_1_m[157]_net_1\, Y => \VDBi_53_0_iv_2[4]_net_1\);
    
    \REGMAP[19]\ : DFF
      port map(CLK => CLK_c_c, D => \un64_reg_ads_0_a3_0_a2\, Q
         => \REGMAP[19]_net_1\);
    
    PIPEA1_582 : MUX2H
      port map(A => N_292, B => \PIPEA1[26]_net_1\, S => 
        un1_STATE2_13_4_0, Y => \PIPEA1_582\);
    
    REG_1_311 : MUX2H
      port map(A => VDB_in_0(1), B => \REG[346]\, S => N_2944_i, 
        Y => \REG_1_311\);
    
    \TCNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \TCNT_10[0]\, CLR => 
        \un10_hwres_33\, Q => \TCNT_i_i[0]\);
    
    \PIPEB_4_i[15]\ : AND2
      port map(A => DPR(15), B => N_616_1, Y => N_2629);
    
    \LB_DOUT[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_173\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[25]_net_1\);
    
    \VDBm_0[15]\ : MUX2H
      port map(A => \PIPEB[15]_net_1\, B => \PIPEA[15]_net_1\, S
         => \BLTCYC_2\, Y => N_2311);
    
    un2_vsel_5_i_a2 : AOI21FTT
      port map(A => N_222_i, B => N_232, C => N_2434_1, Y => 
        N_2436_i);
    
    \PIPEA_m[16]\ : NAND2
      port map(A => N_457_i_0_1, B => \PIPEA[16]_net_1\, Y => 
        \PIPEA_m[16]_net_1\);
    
    \PIPEA[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_620\, CLR => CLEAR_25, 
        Q => \PIPEA[31]_net_1\);
    
    \LB_i_6_1[24]\ : MUX2H
      port map(A => VDB_in(24), B => \LB_DOUT[24]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2206);
    
    \VDBi_16_1_0[8]\ : AO21TTF
      port map(A => \REGMAP_0[2]_net_1\, B => \REG[24]\, C => 
        N_2483, Y => \VDBi_16_1_0_i[8]\);
    
    un10_hwres_5 : OR2
      port map(A => HWRES_c_0_6, B => \WDOGTO\, Y => 
        \un10_hwres_5\);
    
    un1_STATE2_12_0_0_a2_0 : NOR3FFT
      port map(A => \END_PK\, B => \STATE2[1]_net_1\, C => 
        \EVREAD_DS\, Y => N_620_i_i);
    
    \VDBi_92_0_iv_0[28]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[28]_net_1\, C
         => \PIPEA_m[28]_net_1\, Y => \VDBi_92_0_iv_0[28]_net_1\);
    
    \VDBi_23_m[8]\ : AND2
      port map(A => \VDBi_9_sqmuxa_0\, B => \VDBi_23[8]_net_1\, Y
         => \VDBi_23_m_i[8]\);
    
    un57_reg_ads_0_a3_0_a2_0 : NAND2
      port map(A => N_675, B => \WRITES\, Y => N_791);
    
    LB_DOUT_154 : MUX2H
      port map(A => VDB_in(6), B => \LB_DOUT[6]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_154\);
    
    \PIPEA_7_i_m2[4]\ : MUX2H
      port map(A => DPR(4), B => \PIPEA1[4]_net_1\, S => N_1996_2, 
        Y => N_513);
    
    VDBi_9_sqmuxa_i_1 : NOR2
      port map(A => \REGMAP_i_i[17]\, B => \REGMAP[18]_net_1\, Y
         => \VDBi_9_sqmuxa_i_1\);
    
    \REG_1_m[191]\ : NAND2
      port map(A => \REGMAP[20]_net_1\, B => \REG[191]\, Y => 
        \REG_1_m[191]_net_1\);
    
    \VDBi_58_d[0]\ : MUX2H
      port map(A => SPULSE0_c_c, B => L0_c_c, S => 
        \REGMAP[27]_net_1\, Y => \VDBi_58_d[0]_net_1\);
    
    \REG_1_m[241]\ : AND2
      port map(A => \REGMAP_i_i[23]\, B => \REG[241]\, Y => 
        \REG_1_m_i[241]\);
    
    LB_DOUT_0_sqmuxa_0_a2_0_a2_0 : OR2FT
      port map(A => \REGMAP[36]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => LB_DOUT_0_sqmuxa_0);
    
    \VDBi_92_0_iv_0[12]\ : OAI21FTT
      port map(A => N_502, B => N_2613_1, C => 
        \VDBi_92_0_iv_0_1[12]_net_1\, Y => \VDBi_92[12]\);
    
    SINGCYC_1 : DFFC
      port map(CLK => CLK_c_c, D => \SINGCYC_147\, CLR => 
        HWRES_c_21_0, Q => \SINGCYC_1\);
    
    \VDBm_0[8]\ : MUX2H
      port map(A => \PIPEB[8]_net_1\, B => \PIPEA[8]_net_1\, S
         => \BLTCYC_2\, Y => N_2304);
    
    REG_1_405 : MUX2H
      port map(A => VDB_in(31), B => \REG[440]\, S => N_3072_i_0, 
        Y => \REG_1_405\);
    
    REG_1_430 : MUX2H
      port map(A => VDB_in_0(7), B => \REG[489]\, S => N_3170_i, 
        Y => \REG_1_430\);
    
    RAMAD_VME_10 : MUX2H
      port map(A => \VAS[7]_net_1\, B => \RAMAD_VME[6]_net_1\, S
         => N_2523_0, Y => \RAMAD_VME_10\);
    
    \VDBi_16_1_a2[11]\ : AND2
      port map(A => N_2511_0, B => REG_42, Y => N_2488_i);
    
    \VADm[8]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[8]_net_1\, Y => VADm(8));
    
    un7_ronly_0_a3_0_a2_1 : NAND3FTT
      port map(A => N_2369, B => \LWORDS\, C => \VAS[15]_net_1\, 
        Y => un7_ronly_0_a3_0_a2_1_i);
    
    OR_RDATA_184 : MUX2H
      port map(A => N_19, B => \OR_RDATA[2]_net_1\, S => N_1832, 
        Y => \OR_RDATA_184\);
    
    \PIPEA1[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_563\, CLR => CLEAR_23, 
        Q => \PIPEA1[7]_net_1\);
    
    un1_STATE1_28_i : OAI21
      port map(A => \STATE1_0[9]_net_1\, B => LB_DOUT_0_sqmuxa_0, 
        C => \un1_STATE1_28_i_0\, Y => N_2384);
    
    \VADm[3]\ : NOR2FT
      port map(A => \PIPEA[3]_net_1\, B => N_2507_0, Y => VADm(3));
    
    LB_DOUT_153 : MUX2H
      port map(A => VDB_in(5), B => \LB_DOUT[5]_net_1\, S => 
        LB_DOUT_0_sqmuxa, Y => \LB_DOUT_153\);
    
    REG_1_335 : MUX2H
      port map(A => VDB_in(25), B => \REG[370]\, S => N_2944_i_0, 
        Y => \REG_1_335\);
    
    BLTCYC : DFFC
      port map(CLK => CLK_c_c, D => \BLTCYC_77\, CLR => 
        HWRES_c_13, Q => \BLTCYC\);
    
    un776_regmap_19 : NOR2
      port map(A => \REGMAP_0[31]_net_1\, B => 
        \REGMAP_0[28]_net_1\, Y => \un776_regmap_19\);
    
    \REG_1[437]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_402\, CLR => 
        \un10_hwres_23\, Q => \REG[437]\);
    
    un7_cycs_0_a2 : NOR2FT
      port map(A => \CYCS\, B => \TST_c_0[0]\, Y => 
        \un7_cycs_0_a2\);
    
    \REGMAP_1[28]\ : DFF
      port map(CLK => CLK_c_c, D => \un102_reg_ads_0_a3_0_a2\, Q
         => \REGMAP_1[28]_net_1\);
    
    LB_i_521 : MUX2H
      port map(A => \LB_i[9]_net_1\, B => \LB_i_6[9]_net_1\, S
         => N_2570, Y => \LB_i_521\);
    
    WRITES_0 : DFFC
      port map(CLK => CLK_c_c, D => \WRITES_2\, CLR => 
        HWRES_c_23_0, Q => \WRITES_0\);
    
    \REG_i[291]\ : INV
      port map(A => \REG[291]\, Y => REG_i_0_286);
    
    un1_STATE1_15_0_a2 : OR2
      port map(A => \STATE1_0[8]_net_1\, B => \STATE1[9]_net_1\, 
        Y => N_231);
    
    REG_1_409 : MUX2H
      port map(A => VDB_in_0(3), B => \REG[444]\, S => N_3104_i, 
        Y => \REG_1_409\);
    
    \REG_1[373]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_338\, CLR => 
        \un10_hwres_18\, Q => \REG[373]\);
    
    un10_hwres_16 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_16\);
    
    \PIPEA1_9_i[0]\ : AND2
      port map(A => DPR(0), B => N_85, Y => N_238);
    
    \VDBi_16_r[0]\ : OA21TTF
      port map(A => \VDBi_16_1_1_i[0]\, B => N_2377_i, C => 
        \REGMAP_0[7]_net_1\, Y => \VDBi_16[0]\);
    
    \VADm[5]\ : NOR2FT
      port map(A => \PIPEA[5]_net_1\, B => N_2507_0, Y => VADm(5));
    
    VDBi_621 : MUX2H
      port map(A => \VDBi_92[0]\, B => \VDBi[0]_net_1\, S => 
        un1_STATE1_34, Y => \VDBi_621\);
    
    \STATE5_2[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns[0]\, CLR => 
        HWRES_c_21_0, Q => \STATE5_2[0]_net_1\);
    
    REG_1_254 : MUX2H
      port map(A => VDB_in(8), B => \REG[241]\, S => N_2784_i_0, 
        Y => \REG_1_254\);
    
    REG_1_252 : MUX2H
      port map(A => VDB_in(6), B => \REG[239]\, S => N_2784_i, Y
         => \REG_1_252\);
    
    REG_1_494 : MUX2H
      port map(A => \REG_88[87]_net_1\, B => \REG[87]\, S => 
        un1_STATE1_15, Y => \REG_1_494\);
    
    REG_1_361 : MUX2H
      port map(A => VDB_in_0(3), B => \REG[396]\, S => N_3008_i, 
        Y => \REG_1_361\);
    
    \REG_1[410]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_375\, CLR => 
        \un10_hwres_21\, Q => \REG[410]\);
    
    \OR_RDATA[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \OR_RDATA_182\, CLR => 
        HWRES_c_20, Q => \OR_RDATA[0]_net_1\);
    
    REG_1_274 : MUX2H
      port map(A => VDB_in(12), B => \REG[261]\, S => 
        N_2816_i_0_0, Y => \REG_1_274\);
    
    un1_TCNT_1_I_18 : XOR2
      port map(A => \TCNT_i_i[2]\, B => N_83_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_1_0[0]\);
    
    REG_1_272 : MUX2H
      port map(A => VDB_in(10), B => \REG[259]\, S => 
        N_2816_i_0_0, Y => \REG_1_272\);
    
    \REG_1[432]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_397\, CLR => 
        \un10_hwres_23\, Q => \REG[432]\);
    
    \VDBi_23_d[7]\ : MUX2H
      port map(A => \REG[55]\, B => \REG[489]\, S => 
        \REGMAP[13]_net_1\, Y => \VDBi_23_d[7]_net_1\);
    
    PIPEB_49 : MUX2H
      port map(A => \PIPEB[29]_net_1\, B => \PIPEB_4[29]\, S => 
        N_1996_3, Y => \PIPEB_49\);
    
    \REG_1[243]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_256\, SET => 
        \un10_hwres_13\, Q => \REG[243]\);
    
    \VADm[10]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[10]_net_1\, Y => VADm(10));
    
    \STATE5_ns_i_o4_0_o2[2]\ : NAND2
      port map(A => \STATE5[0]_net_1\, B => \STATE5[1]_net_1\, Y
         => N_1861);
    
    \VDBi_92_iv_0[5]\ : AOI21TTF
      port map(A => \RAMDTS[5]_net_1\, B => \STATE1[1]_net_1\, C
         => \FBOUT_m[5]_net_1\, Y => \VDBi_92_iv_0[5]_net_1\);
    
    OR_RDATA_191 : MUX2H
      port map(A => N_33, B => \OR_RDATA[9]_net_1\, S => N_1832, 
        Y => \OR_RDATA_191\);
    
    REG_1_347 : MUX2H
      port map(A => VDB_in_0(5), B => \REG[382]\, S => N_2976_i, 
        Y => \REG_1_347\);
    
    \VDBi[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_635\, CLR => 
        \un10_hwres_34\, Q => \VDBi[14]_net_1\);
    
    \STATE1[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[3]\, CLR => 
        \un10_hwres_32_0\, Q => \STATE1[7]_net_1\);
    
    \PIPEA[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_594\, CLR => CLEAR_25, 
        Q => \PIPEA[5]_net_1\);
    
    \REG_1[158]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_198\, CLR => 
        \un10_hwres_9\, Q => \REG[158]\);
    
    \PIPEA[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_595\, CLR => CLEAR_25, 
        Q => \PIPEA[6]_net_1\);
    
    \STATE1_ns_0[0]\ : OAI21FTT
      port map(A => \STATE1[10]_net_1\, B => N_436, C => 
        \STATE1_ns_0_0[0]_net_1\, Y => \STATE1_ns[0]\);
    
    \REG_1_m[259]\ : NAND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[259]\, Y => 
        \REG_1_m[259]_net_1\);
    
    REG_1_441 : MUX2H
      port map(A => VDB_in(18), B => \REG[500]\, S => N_3170_i_1, 
        Y => \REG_1_441\);
    
    NOEDTKi_192 : MUX2H
      port map(A => NOEDTKi_10, B => \TST_c_c[3]\, S => 
        un1_STATE1_32, Y => \NOEDTKi_192\);
    
    PIPEA_603 : MUX2H
      port map(A => \PIPEA_7[14]\, B => \PIPEA[14]_net_1\, S => 
        un1_STATE2_16_1, Y => \PIPEA_603\);
    
    un1_STATE1_32_0 : AO21TTF
      port map(A => N_2413, B => \STATE1[9]_net_1\, C => 
        \un1_STATE1_32_0_3\, Y => un1_STATE1_32);
    
    REG_1_426 : MUX2H
      port map(A => VDB_in_0(3), B => \REG[485]\, S => N_3170_i, 
        Y => \REG_1_426\);
    
    \REG_1[247]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_260\, SET => 
        \un10_hwres_14\, Q => \REG[247]\);
    
    \REG_1[494]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_435\, SET => 
        \un10_hwres_26\, Q => \REG[494]\);
    
    \VDBi_71[9]\ : MUX2H
      port map(A => \VDBi_66[9]_net_1\, B => \REG[418]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71[9]_net_1\);
    
    \REG_1[180]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_220\, CLR => 
        \un10_hwres_11\, Q => \REG[180]\);
    
    \REG_1[191]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_231\, CLR => 
        \un10_hwres_12\, Q => \REG[191]\);
    
    \VDBi_92_0_iv_0[22]\ : AOI21TTF
      port map(A => \STATE1_0[2]_net_1\, B => \VDBi[22]_net_1\, C
         => \PIPEA_m[22]_net_1\, Y => \VDBi_92_0_iv_0[22]_net_1\);
    
    \LBUSTMO_3_0[3]\ : OR2FT
      port map(A => N_2572_0, B => I_21_1, Y => \LBUSTMO_3[3]\);
    
    un10_hwres_31 : OR2
      port map(A => HWRES_c_0_4, B => WDOGTO_0, Y => 
        \un10_hwres_31\);
    
    \REG_1[63]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_470\, CLR => 
        \un10_hwres_29\, Q => \REG[63]\);
    
    DSSF1 : DFFS
      port map(CLK => CLK_c_c, D => \DSSF1_13\, SET => 
        HWRES_c_13_0, Q => \DSSF1\);
    
    LB_ACK_sync : DFFC
      port map(CLK => CLK_c_c, D => \LB_ACK\, CLR => 
        \un10_hwres_0\, Q => \LB_ACK_sync\);
    
    \PIPEA[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_592\, CLR => CLEAR_25, 
        Q => \PIPEA[3]_net_1\);
    
    \VDBi_18[0]\ : MUX2H
      port map(A => \VDBi_16[0]\, B => \REG[48]\, S => \TST_c[5]\, 
        Y => \VDBi_18[0]_net_1\);
    
    PIPEA_596 : MUX2H
      port map(A => \PIPEA_7[7]\, B => \PIPEA[7]_net_1\, S => 
        un1_STATE2_16, Y => \PIPEA_596\);
    
    un114_reg_ads_0_a3_0_a2_2 : OR2
      port map(A => \VAS[4]_net_1\, B => \VAS[1]_net_1\, Y => 
        N_664);
    
    \PIPEA1[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_580\, CLR => CLEAR_22, 
        Q => \PIPEA1[24]_net_1\);
    
    REG_1_483 : MUX2H
      port map(A => VDB_in(28), B => \REG[76]\, S => N_3234_i_0, 
        Y => \REG_1_483\);
    
    un1_STATE2_8_0_0_0_o2 : NAND2
      port map(A => N_426, B => \STATE2_i_0[3]\, Y => N_1996);
    
    \VDBm_0[4]\ : MUX2H
      port map(A => \PIPEB[4]_net_1\, B => \PIPEA[4]_net_1\, S
         => \BLTCYC\, Y => N_2300);
    
    \REG_1[259]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_272\, CLR => 
        \un10_hwres_15\, Q => \REG[259]\);
    
    \LB_DOUT[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_164\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[16]_net_1\);
    
    \REG_1[135]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_143\, CLR => 
        \un10_hwres_8_0\, Q => \REG[135]\);
    
    \RAMDTS[3]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(3), CLR => HWRES_c_21, 
        Q => \RAMDTS[3]_net_1\);
    
    un1_WDOGRES_0_sqmuxa_0_a2_0_2 : NAND3FTT
      port map(A => \WDOG[0]_net_1\, B => \STATE1[10]_net_1\, C
         => \WDOG[3]_net_1\, Y => un1_WDOGRES_0_sqmuxa_0_a2_0_2_i);
    
    \REG_1[504]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_445\, SET => 
        \un10_hwres_27\, Q => \REG[504]\);
    
    \VDBi_60[14]\ : MUX2H
      port map(A => \VDBi_58[14]_net_1\, B => \REG_c[0]\, S => 
        \REGMAP_1[28]_net_1\, Y => \VDBi_60[14]_net_1\);
    
    \REG_i[287]\ : INV
      port map(A => \REG[287]\, Y => REG_i_0_282);
    
    \VDBi_92_iv_1[0]\ : AO21TTF
      port map(A => N_457_i_0, B => \PIPEA[0]_net_1\, C => 
        \VDBi_92_iv_0[0]_net_1\, Y => \VDBi_92_iv_1_i[0]\);
    
    \VDBi_16_1_0[2]\ : AO21TTF
      port map(A => LOS_c_c, B => \REGMAP_0[2]_net_1\, C => 
        N_2465, Y => \VDBi_16_1_0_i[2]\);
    
    \VDBi_16_1_a2_1[6]\ : NAND2
      port map(A => N_2512, B => \REG[6]\, Y => N_2477);
    
    un1_TCNT_1_I_26 : XOR2
      port map(A => \TCNT_i_i[6]\, B => N_83, Y => 
        \DWACT_ADD_CI_0_partial_sum[6]\);
    
    N_77_i_i_o2_1_2 : NAND3FFT
      port map(A => N_652, B => \END_PK\, C => \MBLTCYC\, Y => 
        N_77_i_i_o2_1_i);
    
    LB_s_84 : MUX2H
      port map(A => LB_in(5), B => \LB_s[5]_net_1\, S => 
        STATE5_0_sqmuxa, Y => \LB_s_84\);
    
    \REG_i[283]\ : INV
      port map(A => \REG[283]\, Y => REG_i_0_278);
    
    \REGMAP_0[2]\ : DFF
      port map(CLK => CLK_c_c, D => \un13_reg_ads_0_a2_0_a2\, Q
         => \REGMAP_0[2]_net_1\);
    
    \REG_1[264]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_277\, CLR => 
        \un10_hwres_15\, Q => \REG[264]\);
    
    \REG_1[262]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_275\, CLR => 
        \un10_hwres_15\, Q => \REG[262]\);
    
    un7_ronly_0_a3_0_a2_0_0 : OR2
      port map(A => \VAS[11]_net_1\, B => \VAS[12]_net_1\, Y => 
        \un7_ronly_0_a3_0_a2_0_0\);
    
    LB_s_98 : MUX2H
      port map(A => LB_in(19), B => \LB_s[19]_net_1\, S => 
        STATE5_0_sqmuxa_1, Y => \LB_s_98\);
    
    \VDBi_23[5]\ : MUX2H
      port map(A => \VDBi_16[5]\, B => \VDBi_23_d[5]_net_1\, S
         => \VDBi_23_s[7]_net_1\, Y => \VDBi_23[5]_net_1\);
    
    \REG_1_m[260]\ : NAND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[260]\, Y => 
        \REG_1_m[260]_net_1\);
    
    un2_vsel_5_i_a2_0 : AND3
      port map(A => AMB_c(1), B => AMB_c(2), C => AMB_c(5), Y => 
        N_222_i);
    
    \REG_1[64]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_471\, CLR => 
        \un10_hwres_29\, Q => \REG[64]\);
    
    \VDBi_53_0_iv_3[6]\ : AO21TTF
      port map(A => \REGMAP[16]_net_1\, B => \REG_0[127]\, C => 
        \VDBi_53_0_iv_2[6]_net_1\, Y => \VDBi_53_0_iv_3_i[6]\);
    
    \STATE1_ns_0_iv_0_a2_0_1[8]\ : NAND2
      port map(A => \REGMAP[10]_net_1\, B => \WRITES\, Y => 
        N_2550_1);
    
    \STATE5_1[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns[0]\, CLR => 
        HWRES_c_21_0, Q => \STATE5_1[0]_net_1\);
    
    \LB_i_6[4]\ : MUX2H
      port map(A => N_2174, B => N_2186, S => LB_i_6_sn_N_2, Y
         => N_2220);
    
    \VDBi_16_1_a2_0[10]\ : AND2
      port map(A => N_2512_0, B => \REG[10]\, Y => N_2487_i);
    
    \VDBi_23_m[6]\ : AND2
      port map(A => \VDBi_9_sqmuxa\, B => \VDBi_23[6]_net_1\, Y
         => \VDBi_23_m_i[6]\);
    
    \LB_i[8]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_520\, CLR => 
        HWRES_c_16, Q => \LB_i[8]_net_1\);
    
    WDOGRES1 : DFFS
      port map(CLK => CLK_c_c, D => \WDOGRES_i\, SET => 
        HWRES_c_23, Q => WDOGRES1_i);
    
    \VDBi_53_0_iv_2[9]\ : AOI21TTF
      port map(A => \REGMAP_0[19]_net_1\, B => \REG[178]\, C => 
        \REG_1_m[162]_net_1\, Y => \VDBi_53_0_iv_2[9]_net_1\);
    
    REG_1_508 : MUX2H
      port map(A => \REG[101]\, B => VDB_in_0(12), S => N_2416_i, 
        Y => \REG_1_508\);
    
    un2_vsel_1_i_a2_1_1 : NAND2FT
      port map(A => AMB_c(4), B => AMB_c(3), Y => 
        un2_vsel_1_i_a2_1_1_i);
    
    \VDBm[6]\ : MUX2H
      port map(A => N_2302, B => \VDBi[6]_net_1\, S => 
        \SINGCYC_2\, Y => VDBm_6);
    
    REG_1_389 : MUX2H
      port map(A => VDB_in_0(15), B => \REG[424]\, S => 
        N_3072_i_1, Y => \REG_1_389\);
    
    \LB_i_6_1[26]\ : MUX2H
      port map(A => VDB_in(26), B => \LB_DOUT[26]_net_1\, S => 
        \STATE5_1[0]_net_1\, Y => N_2208);
    
    un10_hwres_10 : OR2
      port map(A => HWRES_c_0_5, B => WDOGTO_2, Y => 
        \un10_hwres_10\);
    
    \LB_ADDR[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_ADDR_551\, CLR => 
        \un10_hwres_1\, Q => \LB_ADDR[8]_net_1\);
    
    \REG_1[377]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_342\, CLR => 
        \un10_hwres_18\, Q => \REG[377]\);
    
    \STATE5[2]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns_i_0[2]_net_1\, 
        CLR => HWRES_c_22, Q => \STATE5[2]_net_1\);
    
    \STATE2_ns_0_0[4]\ : NAND2
      port map(A => N_580, B => N_725, Y => \STATE2_ns[4]\);
    
    \PIPEA_7_i_m2[12]\ : MUX2H
      port map(A => DPR(12), B => \PIPEA1[12]_net_1\, S => 
        N_1996_1, Y => N_521);
    
    \VDBi_23[18]\ : MUX2H
      port map(A => \VDBi_18[18]_net_1\, B => \REG[500]\, S => 
        \REGMAP_1[13]_net_1\, Y => \VDBi_23[18]_net_1\);
    
    REG_1_143 : MUX2H
      port map(A => \REG[135]\, B => VDB_in(14), S => 
        REG_0_sqmuxa_0, Y => \REG_1_143\);
    
    \PIPEB_4_i[18]\ : AND2
      port map(A => DPR(18), B => N_616_1, Y => N_199);
    
    \VDBi_16_1_a2_0[8]\ : AND2
      port map(A => N_2511_0, B => REG_39, Y => N_2482_i);
    
    \VDBi_53_0_iv_6[0]\ : NOR3
      port map(A => \VDBi_53_0_iv_5_i[0]\, B => 
        \VDBi_53_0_iv_2_i[0]\, C => \VDBi_53_0_iv_0_i[0]\, Y => 
        \VDBi_53_0_iv_6[0]_net_1\);
    
    \PIPEB_4_i[22]\ : AND2
      port map(A => DPR(22), B => N_616_0, Y => N_2634);
    
    REG3_119 : MUX2H
      port map(A => \REG[6]\, B => VDB_in(6), S => REG1_0_sqmuxa, 
        Y => \REG3_119\);
    
    REG1_0_sqmuxa_0_a3_0 : NOR2FT
      port map(A => \REGMAP[1]_net_1\, B => PULSE_0_sqmuxa_1_0, Y
         => REG1_0_sqmuxa_0);
    
    \REG_i[398]\ : INV
      port map(A => \REG[398]\, Y => REG_i_0_393);
    
    un1_REG_0_sqmuxa_i_o2 : OR2
      port map(A => \STATE5_0[0]_net_1\, B => \STATE5[1]_net_1\, 
        Y => N_66);
    
    un1_STATE2_8_0_0_0_o2_4 : NAND2
      port map(A => N_426, B => \STATE2_i_0[3]\, Y => N_1996_4);
    
    \RAMDTS[1]\ : DFFC
      port map(CLK => CLK_c_c, D => RAMDT(1), CLR => HWRES_c_21, 
        Q => \RAMDTS[1]_net_1\);
    
    un12_wdog_0_a3_0 : NAND2
      port map(A => \WDOG_i_0_i[4]\, B => \WDOG[5]_net_1\, Y => 
        un12_wdog_0_a3_0_i);
    
    \REG_1[400]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_365\, CLR => 
        \un10_hwres_20\, Q => \REG[400]\);
    
    \PIPEA[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA_604\, CLR => CLEAR_23, 
        Q => \PIPEA[15]_net_1\);
    
    REG_1_341_e_0 : OR2FT
      port map(A => \REGMAP_0[28]_net_1\, B => PULSE_0_sqmuxa_1_1, 
        Y => N_2944_i_0);
    
    \VDBi_66_0[11]\ : MUX2H
      port map(A => \REG[404]\, B => \REG[388]\, S => 
        \REGMAP_0[29]_net_1\, Y => N_2028);
    
    \PULSE_1[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_245\, CLR => 
        \un10_hwres_4\, Q => \PULSE[10]\);
    
    \REG_1[85]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_492\, CLR => 
        \un10_hwres_31\, Q => \REG[85]\);
    
    \LB_s[30]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_109\, CLR => 
        HWRES_c_19, Q => \LB_s[30]_net_1\);
    
    \VDBi_77_0_i_m2[12]\ : MUX2H
      port map(A => REG_468, B => \REG[453]\, S => 
        \REGMAP_i_i[33]\, Y => N_496);
    
    un1_MYBERRi_1_sqmuxa_0_a2 : NAND2
      port map(A => \STATE1[4]_net_1\, B => \TST_c[2]\, Y => 
        N_2424);
    
    \VDBi_92_0_iv[17]\ : OAI21FTT
      port map(A => \VDBi_71[17]_net_1\, B => N_2613_1, C => 
        \VDBi_92_0_iv_1[17]_net_1\, Y => \VDBi_92[17]\);
    
    \FWIMG2LOAD\ : DFFS
      port map(CLK => CLK_c_c, D => \FWIMG2LOAD_111\, SET => 
        \un10_hwres_0\, Q => FWIMG2LOAD_net_1);
    
    \VDBi_77[15]\ : MUX2H
      port map(A => \VDBi_66[15]_net_1\, B => 
        \VDBi_77_d[15]_net_1\, S => \VDBi_77_s[8]_net_1\, Y => 
        \VDBi_77[15]_net_1\);
    
    LB_DOUT_0_sqmuxa_0_a2_0_a2_1 : OR2FT
      port map(A => \REGMAP[36]_net_1\, B => PULSE_0_sqmuxa_1_0, 
        Y => LB_DOUT_0_sqmuxa_1);
    
    \VDBi_55[19]\ : NOR2FT
      port map(A => \VDBi_23[19]_net_1\, B => 
        \REGMAP_0[26]_net_1\, Y => \VDBi_55[19]_net_1\);
    
    un1_STATE2_12_0_0_2 : OAI21FTF
      port map(A => \STATE2[2]_net_1\, B => N_472_i_0, C => 
        un1_STATE2_12_0_0_1_i, Y => un1_STATE2_13_4_1);
    
    \VDBi_92_0_iv_1[16]\ : AOI21TTF
      port map(A => \LB_s[16]_net_1\, B => N_7_i_1, C => 
        \VDBi_92_0_iv_0[16]_net_1\, Y => 
        \VDBi_92_0_iv_1[16]_net_1\);
    
    \REG_1_m[258]\ : NAND2
      port map(A => \REGMAP_0[24]_net_1\, B => \REG[258]\, Y => 
        \REG_1_m[258]_net_1\);
    
    \PIPEA1_9_i[27]\ : AND2
      port map(A => DPR(27), B => N_85_3, Y => N_294);
    
    \PIPEB_4_i[14]\ : AND2
      port map(A => DPR(14), B => N_616_1, Y => N_2628);
    
    \REG_1[448]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_413\, CLR => 
        \un10_hwres_24\, Q => \REG[448]\);
    
    \STATE1[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[7]\, CLR => 
        \un10_hwres_32\, Q => \STATE1[3]_net_1\);
    
    NRDMEBi : DFFS
      port map(CLK => CLK_c_c, D => \NRDMEBi_588\, SET => 
        CLEAR_20, Q => \NRDMEB\);
    
    \VDBi_23[10]\ : MUX2H
      port map(A => \VDBi_16[10]\, B => \VDBi_23_d[10]_net_1\, S
         => \VDBi_23_s[7]_net_1\, Y => \VDBi_23[10]_net_1\);
    
    \STATE5[1]\ : DFFC
      port map(CLK => ALICLK_c, D => \STATE5_ns[1]\, CLR => 
        HWRES_c_21_0, Q => \STATE5[1]_net_1\);
    
    \PIPEA_7_r[26]\ : AND2
      port map(A => N_85_0, B => N_535, Y => \PIPEA_7[26]\);
    
    N_1897_1 : AOI21TTF
      port map(A => N_1898, B => \WRITES\, C => \N_1897_0\, Y => 
        \N_1897_1\);
    
    \VDBi[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \VDBi_648\, CLR => 
        \un10_hwres_35\, Q => \VDBi[27]_net_1\);
    
    \LB_DOUT[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_157\, CLR => 
        \un10_hwres_3\, Q => \LB_DOUT[9]_net_1\);
    
    \PIPEA1_9_i[6]\ : AND2
      port map(A => DPR(6), B => N_85, Y => N_252);
    
    \PIPEA_7_i_m2[21]\ : MUX2H
      port map(A => DPR(21), B => \PIPEA1[21]_net_1\, S => 
        N_1996_0, Y => N_530);
    
    \VDBi_16_1_0[1]\ : AO21TTF
      port map(A => \REGMAP[2]_net_1\, B => REG_16, C => N_2462, 
        Y => \VDBi_16_1_0_i[1]\);
    
    \STATE1_ns_0_iv_0[7]\ : OAI21FTT
      port map(A => N_2430, B => \REGMAP[36]_net_1\, C => N_2547, 
        Y => \STATE1_ns[7]\);
    
    \REG_1[346]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_311\, SET => 
        \un10_hwres_17\, Q => \REG[346]\);
    
    \REG_1[159]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_199\, CLR => 
        \un10_hwres_9\, Q => \REG[159]\);
    
    \LB_DOUT[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_167\, CLR => 
        \un10_hwres_2\, Q => \LB_DOUT[19]_net_1\);
    
    \VAS[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \VAS_53\, CLR => HWRES_c_22_0, 
        Q => \VAS[2]_net_1\);
    
    \PULSE_1[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_1_243\, CLR => 
        \un10_hwres_4\, Q => \PULSE[8]\);
    
    \PIPEA1_9_0[30]\ : OR2FT
      port map(A => N_85_0, B => DPR(30), Y => \PIPEA1_9[30]\);
    
    REG_1_19_70 : MUX2H
      port map(A => \STATE5[2]_net_1\, B => \REG[19]\, S => N_11, 
        Y => \REG_1_19_70\);
    
    \VDBi_92_0_iv_1[8]\ : AOI21TTF
      port map(A => \LB_s[8]_net_1\, B => N_7_i, C => 
        \VDBi_92_0_iv_0[8]_net_1\, Y => \VDBi_92_0_iv_1[8]_net_1\);
    
    \VDBi_92_iv_1[5]\ : AOI21TTF
      port map(A => N_457_i_0, B => \PIPEA[5]_net_1\, C => 
        \VDBi_92_iv_0[5]_net_1\, Y => \VDBi_92_iv_1[5]_net_1\);
    
    NOEDTKi_10_r : OA21
      port map(A => N_425, B => PULSE_0_sqmuxa_1, C => 
        un1_LB_DOUT_0_sqmuxa, Y => NOEDTKi_10);
    
    \FBOUT_m[4]\ : NAND2
      port map(A => FBOUT(4), B => \STATE1[2]_net_1\, Y => 
        \FBOUT_m[4]_net_1\);
    
    \VDBi_53_0_iv_0[1]\ : AO21TTF
      port map(A => \REGMAP_i_i[17]\, B => REG_137, C => 
        \REG_m[106]_net_1\, Y => \VDBi_53_0_iv_0_i[1]\);
    
    \REG_1[240]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_253\, SET => 
        \un10_hwres_13\, Q => \REG[240]\);
    
    \PIPEA_7_r[13]\ : AND2
      port map(A => N_85_2, B => N_522, Y => \PIPEA_7[13]\);
    
    \REG_1[75]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_482\, CLR => 
        \un10_hwres_30\, Q => \REG[75]\);
    
    REG_1_234 : MUX2H
      port map(A => VDB_in(9), B => \REG[194]\, S => N_2752_i_0, 
        Y => \REG_1_234\);
    
    \VDBi_60[8]\ : MUX2H
      port map(A => \VDBi_60_d[8]_net_1\, B => \VDBi_55[8]_net_1\, 
        S => \VDBi_60_s[5]_net_1\, Y => \VDBi_60[8]_net_1\);
    
    un1_LBUSTMO_1_I_5 : NOR2FT
      port map(A => \LBUSTMO_i_0_i[1]\, B => N_66_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_1[0]\);
    
    REG_1_232 : MUX2H
      port map(A => VDB_in(7), B => \REG[192]\, S => N_2752_i, Y
         => \REG_1_232\);
    
    \LB_i[4]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_i_516\, CLR => 
        HWRES_c_16, Q => \LB_i[4]_net_1\);
    
    ADACKCYC : DFFC
      port map(CLK => CLK_c_c, D => \ADACKCYC_76\, CLR => 
        HWRES_c_12, Q => \ADACKCYC\);
    
    \VDBi_92_iv_0[3]\ : AOI21TTF
      port map(A => \RAMDTS[3]_net_1\, B => \STATE1[1]_net_1\, C
         => \FBOUT_m[3]_net_1\, Y => \VDBi_92_iv_0[3]_net_1\);
    
    \VDBm_0[16]\ : MUX2H
      port map(A => \PIPEB[16]_net_1\, B => \PIPEA[16]_net_1\, S
         => \BLTCYC_2\, Y => N_2312);
    
    \VDBi_77_s[8]\ : OR2
      port map(A => \REGMAP_0[31]_net_1\, B => N_441_0, Y => 
        \VDBi_77_s[8]_net_1\);
    
    \VDBi_23[30]\ : MUX2H
      port map(A => \VDBi_18[30]_net_1\, B => \REG_i[512]_net_1\, 
        S => \REGMAP_0[13]_net_1\, Y => \VDBi_23[30]_net_1\);
    
    un90_reg_ads_0_a3_0_a2 : AND3FTT
      port map(A => un90_reg_ads_0_a3_0_a2_0_i, B => N_688, C => 
        N_674, Y => \un90_reg_ads_0_a3_0_a2\);
    
    \PIPEA1_9_i[5]\ : AND2
      port map(A => DPR(5), B => N_85, Y => N_250);
    
    \REG_1[80]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_487\, CLR => 
        \un10_hwres_30\, Q => \REG[80]\);
    
    PIPEA1_586 : MUX2H
      port map(A => \PIPEA1_9[30]\, B => \PIPEA1[30]_net_1\, S
         => un1_STATE2_13_4_0, Y => \PIPEA1_586\);
    
    PULSE_0_sqmuxa_1_0_a2_0_i2_0_a2_0_a2 : OR2FT
      port map(A => \STATE1_0[8]_net_1\, B => \WRITES_0\, Y => 
        PULSE_0_sqmuxa_1);
    
    \VDBi_77_d[8]\ : MUX2H
      port map(A => \REG[417]\, B => N_2060, S => \N_441\, Y => 
        \VDBi_77_d[8]_net_1\);
    
    REG_1_363 : MUX2H
      port map(A => VDB_in_0(5), B => \REG[398]\, S => N_3008_i, 
        Y => \REG_1_363\);
    
    \REG_1[173]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_213\, CLR => 
        \un10_hwres_10\, Q => \REG[173]\);
    
    \PIPEB[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEB_45\, CLR => CLEAR_27, 
        Q => \PIPEB[25]_net_1\);
    
    \LB_s[19]\ : DFFC
      port map(CLK => ALICLK_c, D => \LB_s_98\, CLR => HWRES_c_17, 
        Q => \LB_s[19]_net_1\);
    
    PIPEB_23 : MUX2H
      port map(A => \PIPEB[3]_net_1\, B => N_2617, S => N_1996, Y
         => \PIPEB_23\);
    
    REG_1_453 : MUX2H
      port map(A => VDB_in(30), B => \REG[512]\, S => N_3170_i_0, 
        Y => \REG_1_453\);
    
    \VADm[14]\ : AND2FT
      port map(A => N_2507, B => \PIPEA[14]_net_1\, Y => VADm(14));
    
    \LB_i_6[8]\ : MUX2H
      port map(A => N_2178, B => N_2190, S => LB_i_6_sn_N_2, Y
         => N_2224);
    
    LB_DOUT_175 : MUX2H
      port map(A => VDB_in(27), B => \LB_DOUT[27]_net_1\, S => 
        LB_DOUT_0_sqmuxa_0, Y => \LB_DOUT_175\);
    
    PULSE_1_243 : MUX2H
      port map(A => N_2386, B => \PULSE[8]\, S => un1_STATE1_17, 
        Y => \PULSE_1_243\);
    
    REG_1_473 : MUX2H
      port map(A => VDB_in(18), B => \REG[66]\, S => N_3234_i_1, 
        Y => \REG_1_473\);
    
    \REG_1[285]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_298\, CLR => 
        \un10_hwres_16\, Q => \REG[285]\);
    
    \PIPEA1[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PIPEA1_557\, CLR => CLEAR_21, 
        Q => \PIPEA1[1]_net_1\);
    
    \VDBi_53_0_iv_1[4]\ : AO21TTF
      port map(A => \REGMAP_i_i_0[23]\, B => \REG[237]\, C => 
        \REG_1_m[189]_net_1\, Y => \VDBi_53_0_iv_1_i[4]\);
    
    \VDBi_71_d[4]\ : MUX2H
      port map(A => N_2021, B => \REG[413]\, S => 
        \REGMAP[31]_net_1\, Y => \VDBi_71_d[4]_net_1\);
    
    \REG_1[256]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_269\, CLR => 
        \un10_hwres_14\, Q => \REG[256]\);
    
    \VDBi_92_0_iv_0_1[31]\ : AO21TTF
      port map(A => N_457_i_0_0, B => \PIPEA[31]_net_1\, C => 
        N_615, Y => \VDBi_92_0_iv_0_1_i[31]\);
    
    \REG_88[81]\ : NOR2FT
      port map(A => N_2152, B => N_2566, Y => \REG_88[81]_net_1\);
    
    \REG_1[430]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_395\, CLR => 
        \un10_hwres_23\, Q => \REG[430]\);
    
    \LB_DOUT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \LB_DOUT_148\, CLR => 
        \un10_hwres_1\, Q => \LB_DOUT[0]_net_1\);
    
    REG3_124 : MUX2H
      port map(A => \REG[11]\, B => VDB_in(11), S => 
        REG1_0_sqmuxa_0, Y => \REG3_124\);
    
    \VADm[0]\ : NOR2FT
      port map(A => \PIPEA[0]_net_1\, B => N_2507_0, Y => VADm(0));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity CROM is

    port( CROMWDT   : in    std_logic_vector(7 downto 0);
          RAMAD_VME : in    std_logic_vector(8 downto 0);
          CROMWAD   : in    std_logic_vector(8 downto 0);
          RAMDT     : out   std_logic_vector(7 downto 0);
          WRCROM    : in    std_logic;
          RAMRD     : in    std_logic;
          CLK_c_c   : in    std_logic
        );

end CROM;

architecture DEF_ARCH of CROM is 

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DMUX
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFF
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM256x9SSTP
    generic (MEMORYFILE:string := "");

    port( DO8    : out   std_logic;
          DO7    : out   std_logic;
          DO6    : out   std_logic;
          DO5    : out   std_logic;
          DO4    : out   std_logic;
          DO3    : out   std_logic;
          DO2    : out   std_logic;
          DO1    : out   std_logic;
          DO0    : out   std_logic;
          DOS    : out   std_logic;
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          DI8    : in    std_logic := 'U';
          DI7    : in    std_logic := 'U';
          DI6    : in    std_logic := 'U';
          DI5    : in    std_logic := 'U';
          DI4    : in    std_logic := 'U';
          DI3    : in    std_logic := 'U';
          DI2    : in    std_logic := 'U';
          DI1    : in    std_logic := 'U';
          DI0    : in    std_logic := 'U';
          WRB    : in    std_logic := 'U';
          RDB    : in    std_logic := 'U';
          WBLKB  : in    std_logic := 'U';
          RBLKB  : in    std_logic := 'U';
          PARODD : in    std_logic := 'U';
          WCLKS  : in    std_logic := 'U';
          RCLKS  : in    std_logic := 'U';
          DIS    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal net00048, net00047, net00013, net00046, net00011, 
        net00043, net00042, net00041, \GND\, net00038, net00037, 
        net00036, net00033, net00032, net00031, net00028, 
        net00027, net00026, net00023, net00022, net00021, 
        net00018, net00017, net00016, net00012, net00010, 
        net00009, net00004, net00002, net00003, net00052, 
        net00050, \VCC\ : std_logic;

begin 


    U2 : MUX2H
      port map(A => RAMAD_VME(8), B => net00002, S => RAMRD, Y
         => net00003);
    
    U6 : DMUX
      port map(A => net00009, B => \GND\, S => net00011, Y => 
        net00010);
    
    U20 : DMUX
      port map(A => net00046, B => \GND\, S => net00011, Y => 
        net00047);
    
    U19 : DMUX
      port map(A => net00043, B => net00042, S => net00013, Y => 
        RAMDT(6));
    
    U9 : DMUX
      port map(A => net00018, B => net00017, S => net00013, Y => 
        RAMDT(1));
    
    U3 : DFF
      port map(CLK => CLK_c_c, D => net00003, Q => net00002);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    U4 : INV
      port map(A => CROMWAD(8), Y => net00004);
    
    U17 : DMUX
      port map(A => net00038, B => net00037, S => net00013, Y => 
        RAMDT(5));
    
    U15 : DMUX
      port map(A => net00033, B => net00032, S => net00013, Y => 
        RAMDT(4));
    
    M1 : RAM256x9SSTP
      generic map(MEMORYFILE => "CROM_M1.mem")

      port map(DO8 => net00052, DO7 => net00048, DO6 => net00043, 
        DO5 => net00038, DO4 => net00033, DO3 => net00028, DO2
         => net00023, DO1 => net00018, DO0 => net00012, DOS => 
        net00013, WADDR7 => CROMWAD(7), WADDR6 => CROMWAD(6), 
        WADDR5 => CROMWAD(5), WADDR4 => CROMWAD(4), WADDR3 => 
        CROMWAD(3), WADDR2 => CROMWAD(2), WADDR1 => CROMWAD(1), 
        WADDR0 => CROMWAD(0), RADDR7 => RAMAD_VME(7), RADDR6 => 
        RAMAD_VME(6), RADDR5 => RAMAD_VME(5), RADDR4 => 
        RAMAD_VME(4), RADDR3 => RAMAD_VME(3), RADDR2 => 
        RAMAD_VME(2), RADDR1 => RAMAD_VME(1), RADDR0 => 
        RAMAD_VME(0), DI8 => \GND\, DI7 => CROMWDT(7), DI6 => 
        CROMWDT(6), DI5 => CROMWDT(5), DI4 => CROMWDT(4), DI3 => 
        CROMWDT(3), DI2 => CROMWDT(2), DI1 => CROMWDT(1), DI0 => 
        CROMWDT(0), WRB => WRCROM, RDB => RAMRD, WBLKB => 
        CROMWAD(8), RBLKB => \GND\, PARODD => \GND\, WCLKS => 
        CLK_c_c, RCLKS => CLK_c_c, DIS => net00002);
    
    U14 : DMUX
      port map(A => net00031, B => \GND\, S => net00011, Y => 
        net00032);
    
    U10 : DMUX
      port map(A => net00021, B => \GND\, S => net00011, Y => 
        net00022);
    
    U8 : DMUX
      port map(A => net00016, B => \GND\, S => net00011, Y => 
        net00017);
    
    U13 : DMUX
      port map(A => net00028, B => net00027, S => net00013, Y => 
        RAMDT(3));
    
    GND_i : GND
      port map(Y => \GND\);
    
    U21 : DMUX
      port map(A => net00048, B => net00047, S => net00013, Y => 
        RAMDT(7));
    
    U12 : DMUX
      port map(A => net00026, B => \GND\, S => net00011, Y => 
        net00027);
    
    U18 : DMUX
      port map(A => net00041, B => \GND\, S => net00011, Y => 
        net00042);
    
    M0 : RAM256x9SSTP
      generic map(MEMORYFILE => "CROM_M0.mem")

      port map(DO8 => net00050, DO7 => net00046, DO6 => net00041, 
        DO5 => net00036, DO4 => net00031, DO3 => net00026, DO2
         => net00021, DO1 => net00016, DO0 => net00009, DOS => 
        net00011, WADDR7 => CROMWAD(7), WADDR6 => CROMWAD(6), 
        WADDR5 => CROMWAD(5), WADDR4 => CROMWAD(4), WADDR3 => 
        CROMWAD(3), WADDR2 => CROMWAD(2), WADDR1 => CROMWAD(1), 
        WADDR0 => CROMWAD(0), RADDR7 => RAMAD_VME(7), RADDR6 => 
        RAMAD_VME(6), RADDR5 => RAMAD_VME(5), RADDR4 => 
        RAMAD_VME(4), RADDR3 => RAMAD_VME(3), RADDR2 => 
        RAMAD_VME(2), RADDR1 => RAMAD_VME(1), RADDR0 => 
        RAMAD_VME(0), DI8 => \GND\, DI7 => CROMWDT(7), DI6 => 
        CROMWDT(6), DI5 => CROMWDT(5), DI4 => CROMWDT(4), DI3 => 
        CROMWDT(3), DI2 => CROMWDT(2), DI1 => CROMWDT(1), DI0 => 
        CROMWDT(0), WRB => WRCROM, RDB => RAMRD, WBLKB => 
        net00004, RBLKB => \GND\, PARODD => \GND\, WCLKS => 
        CLK_c_c, RCLKS => CLK_c_c, DIS => \GND\);
    
    U16 : DMUX
      port map(A => net00036, B => \GND\, S => net00011, Y => 
        net00037);
    
    U11 : DMUX
      port map(A => net00023, B => net00022, S => net00013, Y => 
        RAMDT(2));
    
    U7 : DMUX
      port map(A => net00012, B => net00010, S => net00013, Y => 
        RAMDT(0));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity RESET_MOD is

    port( TICK_2_d0     : out   std_logic;
          TICK_1_d0     : out   std_logic;
          TICK_0_d0     : out   std_logic;
          LBSP_c        : out   std_logic_vector(2 to 2);
          PULSE         : in    std_logic_vector(1 to 1);
          LBSP_c_0      : out   std_logic_vector(2 to 2);
          LBSP_c_1      : out   std_logic_vector(2 to 2);
          TST_c         : out   std_logic_vector(15 downto 13);
          TICK_0_2      : out   std_logic;
          TICK_0_0      : out   std_logic;
          TICK_1        : out   std_logic_vector(0 to 0);
          TICK_2        : out   std_logic_vector(0 to 0);
          REG_464       : out   std_logic;
          REG_463       : out   std_logic;
          REG_462       : out   std_logic;
          REG_461       : out   std_logic;
          REG_460       : out   std_logic;
          REG_459       : out   std_logic;
          REG_458       : out   std_logic;
          REG_456       : out   std_logic;
          REG_455       : out   std_logic;
          REG_454       : out   std_logic;
          REG_453       : out   std_logic;
          REG_451       : out   std_logic;
          REG_457       : out   std_logic;
          REG_452       : out   std_logic;
          REG_449       : out   std_logic;
          REG_450       : out   std_logic;
          REG_0         : in    std_logic;
          PON_LOAD_i    : out   std_logic;
          EV_RES_c      : out   std_logic;
          RUN_c         : in    std_logic;
          LOAD_RES      : in    std_logic;
          CLEAR         : out   std_logic;
          BNCRES_c      : in    std_logic;
          EVRES_c       : in    std_logic;
          WDOGTO        : in    std_logic;
          HWRES_c       : out   std_logic;
          HWRES_c_i_0   : out   std_logic;
          CLEAR_i_0     : out   std_logic;
          RUN_c_0       : in    std_logic;
          ALICLK_c      : in    std_logic;
          HWRES_c_0     : out   std_logic;
          HWRES_c_1     : out   std_logic;
          HWRES_c_2     : out   std_logic;
          HWRES_c_3     : out   std_logic;
          HWRES_c_4     : out   std_logic;
          HWRES_c_5     : out   std_logic;
          NPWON_c       : in    std_logic;
          HWRES_c_6     : out   std_logic;
          HWRES_c_7     : out   std_logic;
          HWRES_c_8     : out   std_logic;
          HWRES_c_9     : out   std_logic;
          HWRES_c_10    : out   std_logic;
          HWRES_c_11    : out   std_logic;
          HWRES_c_12    : out   std_logic;
          HWRES_c_13    : out   std_logic;
          HWRES_c_14    : out   std_logic;
          HWRES_c_15    : out   std_logic;
          HWRES_c_16    : out   std_logic;
          HWRES_c_17    : out   std_logic;
          HWRES_c_18    : out   std_logic;
          HWRES_c_19    : out   std_logic;
          HWRES_c_20    : out   std_logic;
          HWRES_c_21    : out   std_logic;
          HWRES_c_22    : out   std_logic;
          HWRES_c_23    : out   std_logic;
          HWRES_c_24    : out   std_logic;
          HWRES_c_25    : out   std_logic;
          HWRES_c_26    : out   std_logic;
          HWRES_c_27    : out   std_logic;
          HWRES_c_28    : out   std_logic;
          HWRES_c_29    : out   std_logic;
          HWRES_c_30    : out   std_logic;
          HWRES_c_31    : out   std_logic;
          HWRES_c_32    : out   std_logic;
          HWRES_c_33    : out   std_logic;
          HWRES_c_34    : out   std_logic;
          HWRES_c_35    : out   std_logic;
          HWRES_c_36    : out   std_logic;
          CLEAR_0       : out   std_logic;
          CLEAR_2       : out   std_logic;
          CLEAR_3       : out   std_logic;
          CLEAR_4       : out   std_logic;
          CLEAR_5       : out   std_logic;
          CLEAR_6       : out   std_logic;
          CLEAR_7       : out   std_logic;
          CLEAR_8       : out   std_logic;
          LOAD_RES_2    : in    std_logic;
          CLEAR_9       : out   std_logic;
          CLEAR_10      : out   std_logic;
          CLEAR_11      : out   std_logic;
          CLEAR_12      : out   std_logic;
          CLEAR_13      : out   std_logic;
          CLEAR_14      : out   std_logic;
          CLEAR_15      : out   std_logic;
          CLEAR_16      : out   std_logic;
          CLEAR_17      : out   std_logic;
          CLEAR_18      : out   std_logic;
          LOAD_RES_1    : in    std_logic;
          CLEAR_19      : out   std_logic;
          CLEAR_20      : out   std_logic;
          CLEAR_21      : out   std_logic;
          CLEAR_22      : out   std_logic;
          CLEAR_23      : out   std_logic;
          CLEAR_24      : out   std_logic;
          CLEAR_25      : out   std_logic;
          CLEAR_26      : out   std_logic;
          CLEAR_27      : out   std_logic;
          LOAD_RES_0    : in    std_logic;
          CLEAR_28      : out   std_logic;
          HWRES_c_36_0  : out   std_logic;
          HWRES_c_32_0  : out   std_logic;
          NPWON_c_1     : in    std_logic;
          HWRES_c_23_0  : out   std_logic;
          HWRES_c_22_0  : out   std_logic;
          HWRES_c_21_0  : out   std_logic;
          HWRES_c_13_0  : out   std_logic;
          HWRES_c_10_0  : out   std_logic;
          HWRES_c_0_0   : out   std_logic;
          HWRES_c_0_2   : out   std_logic;
          HWRES_c_0_3   : out   std_logic;
          HWRES_c_0_4   : out   std_logic;
          HWRES_c_0_5   : out   std_logic;
          HWRES_c_0_6   : out   std_logic;
          RUN_c_0_0     : in    std_logic;
          NLBCLR_c      : out   std_logic;
          SYSRESB_c     : in    std_logic;
          CLK_c_c       : in    std_logic;
          NPWON_c_2     : in    std_logic;
          HWRES_c_27_0  : out   std_logic;
          NPWON_c_3     : in    std_logic;
          HWRES_c_7_0   : out   std_logic;
          NPWON_c_0     : in    std_logic;
          HWRES_c_0_6_0 : out   std_logic
        );

end RESET_MOD;

architecture DEF_ARCH of RESET_MOD is 

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFF
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NAND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_259_0, \TST_c_0[15]\, N_259_3, \TST_c_3[15]\, 
        N_259_2, \TST_c_2[15]\, LongSoftPON_1_i, \TST_c_1[15]\, 
        N_259_1, CLEAR_0_i_1, CLEAR_0_i_0, \NLBCLR_c\, 
        HWRES_c_0_1, N_269_i_0, \un12_tcnt3_i\, \HWRES_c_0_0\, 
        CLEAR_0_i, \HWRES_c_0_2\, \CLEAR_1\, stop2_1, 
        stop2_40_i_a3, stop2_0, N_259, \TST_c[15]\, un8_hwresi_i, 
        \BNC_RESi_1\, \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_TMP[0]\, \TCNT2[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, 
        \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, \TCNT2_i_i[4]\, 
        \DWACT_ADD_CI_0_g_array_12[0]\, \TCNT2_i_i[2]\, 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, \TCNT2_i_i[6]\, 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, 
        \DWACT_ADD_CI_0_TMP_0[0]\, \TCNT3[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_2_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_11_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_12_1_0[0]\, \TCNT3_i_i[4]\, 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, \TCNT3_i_i[2]\, 
        \DWACT_ADD_CI_0_g_array_12_2_0[0]\, \TCNT3_i_i[6]\, 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, 
        \DWACT_ADD_CI_0_TMP_1[0]\, \TCNT4[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, \TCNT4_i_0_i[2]\, N_63, 
        N_55, \DWACT_FINC_E[0]\, N_32, \DWACT_FINC_E[4]\, N_17, 
        \DWACT_FINC_E[7]\, \DWACT_FINC_E[6]\, N_157, 
        \cnt2[1]_net_1\, \cnt2[0]_net_1\, N_149, \cnt2[3]\, 
        \DWACT_FINC_E_0[0]\, N_126, \cnt2[8]\, 
        \DWACT_FINC_E_0[4]\, N_111, \DWACT_FINC_E_0[7]\, 
        \DWACT_FINC_E_0[6]\, N_7, \cnt1[1]\, \cnt1[0]\, N_15, 
        \TCNT1_i_i[1]\, \TCNT1[0]_net_1\, N_7_0, \TCNT1[3]_net_1\, 
        \DWACT_FINC_E_1[0]\, \stop_0_sqmuxa_i\, \stop_0_sqmuxa\, 
        N_270_i_0, \un10_tcnt2_i_o3\, un6_tcnt1_i_0_2_i, 
        un6_tcnt1_i_0_1_i, \TCNT1_i_i[2]\, \TCNT1_i_i[4]\, 
        \TCNT1[5]_net_1\, \HWRES_c_0\, CLEAR_0_net_1, \HWRES_c_3\, 
        \HWCLEARi_2\, un7_stop2_i, \un11_tcnt3_i_0\, 
        un10_tcnt2_i_o3_4_i, un10_tcnt2_i_o3_5_i, 
        un10_tcnt2_i_o3_0_i, \TCNT2[5]_net_1\, \TCNT2[7]_net_1\, 
        un10_tcnt2_i_o3_2_i, \TCNT2_i_i[0]\, \TCNT2[3]_net_1\, 
        cnt2_39, \cnt2_2_i_i[31]\, \cnt2[31]\, cnt2_38, 
        \cnt2_2[30]\, \cnt2[30]\, cnt2_37, \cnt2_2_i_i[29]\, 
        \cnt2[29]\, cnt2_36, \cnt2_2[28]\, \cnt2[28]\, cnt2_35, 
        \cnt2_2[27]\, \cnt2[27]\, cnt2_34, \cnt2_2[26]\, 
        \cnt2[26]\, cnt2_33, \cnt2_2_i_i[25]\, \cnt2[25]\, 
        cnt2_32, \cnt2_2[24]\, \cnt2[24]\, cnt2_31, 
        \cnt2_2_i_i[23]\, \cnt2[23]\, cnt2_30, \cnt2_2[22]\, 
        \cnt2[22]\, cnt2_29, \cnt2_2_i_i[21]\, \cnt2[21]\, 
        cnt2_28, \cnt2_2[20]\, \cnt2[20]\, cnt2_27, 
        \cnt2_2_i_i[19]\, \cnt2[19]\, cnt2_26, \cnt2_2[18]\, 
        \cnt2[18]\, cnt2_25, \cnt2_2[17]\, \cnt2[17]\, cnt2_24, 
        \cnt2_2[16]\, \cnt2[16]\, cnt2_23, \cnt2_2_i_i[15]\, 
        \cnt2[15]\, cnt2_22, \cnt2_2[14]\, \cnt2[14]\, cnt2_21, 
        \cnt2_2_i_i[13]\, \cnt2[13]\, cnt2_20, \cnt2_2[12]\, 
        \cnt2[12]\, cnt2_19, \cnt2_2[11]\, \cnt2[11]\, stop2, 
        cnt2_18, \cnt2_2[10]\, \cnt2[10]\, cnt2_17, \cnt2_2[9]\, 
        \cnt2[9]\, cnt2_16, \cnt2_2[8]\, cnt2_15, \cnt2_2[7]\, 
        \cnt2[7]\, cnt2_14, \cnt2_2[6]\, \cnt2[6]\, cnt2_13, 
        \cnt2_2[5]\, \cnt2[5]\, cnt2_12, \cnt2_2[4]\, \cnt2[4]\, 
        cnt2_11, \cnt2_2[3]\, cnt2_10, \cnt2_2[2]\, \cnt2[2]\, 
        cnt2_9, \cnt2_2[1]\, cnt2_8, \cnt2_2[0]\, \stop_7\, 
        \stop\, \cnt2_0[1]\, \un4_ticki\, \cnt2_0[0]\, cnt1_6, 
        I_13_2, \cnt1[3]\, \un1_stop2_1_0\, cnt1_5, I_9_1, 
        \cnt1[2]\, cnt1_4, I_5_1, cnt1_3, I_4_1, stop1, \cnt2_2\, 
        N_254, \cnt2_1\, \TICK[3]\, \SoftPON_2_0\, 
        \SoftPON_2_0_a3_0\, \SoftPON_2_0_a3\, \TST_c[14]\, 
        un3_stop2_i, un7_stop2_i_29_i, un7_stop2_i_25_i, 
        un7_stop2_i_24_i, un7_stop2_i_17_i, un7_stop2_i_19, 
        un7_stop2_i_7_i, un7_stop2_i_6_i, un7_stop2_i_4, 
        un7_stop2_i_2_i, un7_stop2_i_1, un7_stop2_i_26_i, 
        un7_stop2_i_23_i, un7_stop2_i_21_i, un7_stop2_i_8_i, 
        un7_stop2_i_9_i, un7_stop2_i_10_i, un7_stop2_i_20_i, 
        un7_stop2_i_12_i, stop1_1_0, un3_stop2_i_0, 
        \un15_tcnt4_0_a3\, un15_tcnt4_0_a3_2_i, 
        un11_tcnt3_i_0_4_i, un11_tcnt3_i_0_0_i, 
        un11_tcnt3_i_0_1_i, \TCNT3[5]_net_1\, \TCNT3[7]_net_1\, 
        un11_tcnt3_i_0_2_i, \TCNT3_i_i[0]\, \TCNT3[3]_net_1\, 
        un15_tcnt4_0_a3_0_i, \TCNT4_i_0_i[0]\, \TCNT4[3]_net_1\, 
        \EV_RESi_1\, \EV_RES1\, \BNC_RES1\, \TST_c[13]\, I_4_0, 
        I_5_0, I_9_0, I_13_1, I_20_0, I_24_0, 
        \DWACT_ADD_CI_0_partial_sum[0]\, \TCNT2_2[1]\, 
        \TCNT2_2[2]\, \TCNT2_2[3]\, \TCNT2_2[4]\, \TCNT2_2[5]\, 
        \TCNT2_2[6]\, \TCNT2_2[7]\, 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, \TCNT3_2[1]\, 
        \TCNT3_2[2]\, \TCNT3_2[3]\, \TCNT3_2[4]\, \TCNT3_2[5]\, 
        \TCNT3_2[6]\, \TCNT3_2[7]\, \REG[457]\, I_4, \REG[458]\, 
        I_5, I_9, \REG[460]\, I_13_0, I_20, I_24, CLEAR_2_net_1, 
        I_31, I_38, \REG[465]\, I_45, I_52, I_56, I_66, I_73, 
        I_77, I_84, I_91, \DWACT_ADD_CI_0_partial_sum_1[0]\, 
        \TCNT4_2[1]\, \TCNT4_2[2]\, \TCNT4_2[3]\, \TICK[2]\, N_4, 
        N_12, N_4_0, N_4_1, \DWACT_FINC_E[24]\, 
        \DWACT_FINC_E[23]\, \DWACT_FINC_E[27]\, 
        \DWACT_FINC_E[26]\, N_9, N_14, \DWACT_FINC_E[25]\, N_19, 
        \DWACT_FINC_E[29]\, \DWACT_FINC_E[30]\, N_24, 
        \DWACT_FINC_E[15]\, \DWACT_FINC_E[17]\, 
        \DWACT_FINC_E[22]\, N_31, \DWACT_FINC_E[21]\, 
        \DWACT_FINC_E[9]\, \DWACT_FINC_E[12]\, \DWACT_FINC_E[20]\, 
        N_40, \DWACT_FINC_E[13]\, \DWACT_FINC_E[19]\, N_45, 
        \DWACT_FINC_E[18]\, N_52, \DWACT_FINC_E[33]\, 
        \DWACT_FINC_E[34]\, \DWACT_FINC_E[2]\, \DWACT_FINC_E[5]\, 
        N_61, \DWACT_FINC_E[28]\, \DWACT_FINC_E[16]\, N_66, N_71, 
        \DWACT_FINC_E[14]\, N_76, N_81, \DWACT_FINC_E[10]\, N_88, 
        \DWACT_FINC_E[11]\, N_93, N_98, N_103, \DWACT_FINC_E[8]\, 
        N_108, N_116, N_123, \DWACT_FINC_E[3]\, N_131, N_136, 
        N_141, \DWACT_FINC_E[1]\, N_146, N_154, N_4_2, \REG[472]\, 
        \DWACT_FINC_E_0[9]\, \REG[469]\, \REG[470]\, \REG[471]\, 
        N_9_0, \DWACT_FINC_E_0[8]\, N_14_0, \REG[466]\, 
        \REG[467]\, \REG[468]\, N_22, \DWACT_FINC_E_0[2]\, 
        \DWACT_FINC_E_0[5]\, \REG[463]\, \REG[464]\, N_29, 
        \DWACT_FINC_E_0[3]\, N_37, N_42, \REG[461]\, \REG[462]\, 
        N_47, \DWACT_FINC_E_0[1]\, N_52_0, \REG[459]\, N_60, 
        \TICK[1]\, \TICK[0]\, \GND\, \VCC\ : std_logic;

begin 

    TICK_2_d0 <= \TICK[2]\;
    TICK_1_d0 <= \TICK[1]\;
    TICK_0_d0 <= \TICK[0]\;
    TST_c(15) <= \TST_c[15]\;
    TST_c(14) <= \TST_c[14]\;
    TST_c(13) <= \TST_c[13]\;
    REG_464 <= \REG[472]\;
    REG_463 <= \REG[471]\;
    REG_462 <= \REG[470]\;
    REG_461 <= \REG[469]\;
    REG_460 <= \REG[468]\;
    REG_459 <= \REG[467]\;
    REG_458 <= \REG[466]\;
    REG_456 <= \REG[464]\;
    REG_455 <= \REG[463]\;
    REG_454 <= \REG[462]\;
    REG_453 <= \REG[461]\;
    REG_451 <= \REG[459]\;
    REG_457 <= \REG[465]\;
    REG_452 <= \REG[460]\;
    REG_449 <= \REG[457]\;
    REG_450 <= \REG[458]\;
    HWRES_c_0 <= \HWRES_c_0\;
    HWRES_c_3 <= \HWRES_c_3\;
    CLEAR_0 <= CLEAR_0_net_1;
    CLEAR_2 <= CLEAR_2_net_1;
    HWRES_c_0_0 <= \HWRES_c_0_0\;
    HWRES_c_0_2 <= \HWRES_c_0_2\;
    NLBCLR_c <= \NLBCLR_c\;

    un2_hwresi_0 : OR2
      port map(A => REG_0, B => SYSRESB_c, Y => N_259_0);
    
    SOFT_PON_GENERATE_cnt2_11 : MUX2H
      port map(A => \cnt2_2[3]\, B => \cnt2[3]\, S => stop2, Y
         => cnt2_11);
    
    HWRES_27 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_27);
    
    HWRES_36_0 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_36_0);
    
    \CLEAR\ : OR3FTT
      port map(A => LOAD_RES, B => \HWRES_c_0\, C => CLEAR_0_i, Y
         => CLEAR);
    
    un1_tcnt1_I_19 : AND2
      port map(A => \TCNT1[3]_net_1\, B => \DWACT_FINC_E_1[0]\, Y
         => N_7_0);
    
    \TCNT2[3]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT2_2[3]\, Q => 
        \TCNT2[3]_net_1\);
    
    SOFT_PON_GENERATE_cnt2_17 : MUX2H
      port map(A => \cnt2_2[9]\, B => \cnt2[9]\, S => stop2, Y
         => cnt2_17);
    
    un10_tcnt2_i_o3 : NAND3FFT
      port map(A => un10_tcnt2_i_o3_4_i, B => un10_tcnt2_i_o3_5_i, 
        C => N_269_i_0, Y => \un10_tcnt2_i_o3\);
    
    \TICKi[2]\ : DFF
      port map(CLK => CLK_c_c, D => \un12_tcnt3_i\, Q => 
        \TICK[2]\);
    
    un2_cnt2_1_SUM1 : XOR2
      port map(A => \cnt2_0[0]\, B => \cnt2_0[1]\, Y => N_254);
    
    SOFT_PON_GENERATE_cnt2_39 : MUX2H
      port map(A => \cnt2_2_i_i[31]\, B => \cnt2[31]\, S => 
        stop2_0, Y => cnt2_39);
    
    \CLEAR_7\ : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => CLEAR_7);
    
    BNC_RESi_1_0 : DFFC
      port map(CLK => ALICLK_c, D => \BNC_RESi_1\, CLR => 
        un8_hwresi_i, Q => LBSP_c_1(2));
    
    HWRES_35 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_35);
    
    un6_tcnt1_i_0_1 : OR2
      port map(A => \TCNT1_i_i[2]\, B => \TCNT1[3]_net_1\, Y => 
        un6_tcnt1_i_0_1_i);
    
    TCNT4_2_I_19 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_1[0]\, B => 
        \TCNT4[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1_1[0]\);
    
    \TCNT1[0]\ : DFF
      port map(CLK => CLK_c_c, D => I_4_0, Q => \TCNT1[0]_net_1\);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_6 : NAND3
      port map(A => un7_stop2_i_4, B => \cnt2_2[4]\, C => 
        \cnt2_2[5]\, Y => un7_stop2_i_6_i);
    
    HWRES_23_0 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_23_0);
    
    cnt2_2_0_I_84 : XOR2
      port map(A => N_103, B => \cnt2[14]\, Y => \cnt2_2[14]\);
    
    un3_activity_I_37 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E_0[2]\, 
        C => \REG[463]\, Y => N_42);
    
    cnt2_2_0_I_41 : AND2
      port map(A => \cnt2[6]\, B => \cnt2[7]\, Y => 
        \DWACT_FINC_E[3]\);
    
    HWRES_13 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_13);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_23 : OR3
      port map(A => un7_stop2_i_9_i, B => un7_stop2_i_10_i, C => 
        \cnt2_2[28]\, Y => un7_stop2_i_23_i);
    
    un10_tcnt2_i_o3_5 : OR3
      port map(A => un10_tcnt2_i_o3_0_i, B => \TCNT2_i_i[4]\, C
         => \TCNT2[5]_net_1\, Y => un10_tcnt2_i_o3_5_i);
    
    cnt2_2_0_I_179 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        C => \DWACT_FINC_E[20]\, Y => \DWACT_FINC_E[21]\);
    
    un3_activity_I_66 : XOR2
      port map(A => N_22, B => \REG[468]\, Y => I_66);
    
    un3_activity_I_55 : AND3
      port map(A => \DWACT_FINC_E[4]\, B => \REG[465]\, C => 
        \REG[466]\, Y => N_29);
    
    cnt2_2_0_I_77 : XOR2
      port map(A => N_108, B => \cnt2[13]\, Y => \cnt2_2_i_i[13]\);
    
    SOFT_PON_GENERATE_cnt2_21 : MUX2H
      port map(A => \cnt2_2_i_i[13]\, B => \cnt2[13]\, S => 
        stop2_1, Y => cnt2_21);
    
    TCNT2_2_I_39 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    cnt2_2_0_I_5 : XOR2
      port map(A => \cnt2[0]_net_1\, B => \cnt2[1]_net_1\, Y => 
        \cnt2_2[1]\);
    
    \ACTIVITY[15]\ : DFFC
      port map(CLK => ALICLK_c, D => I_91, CLR => \CLEAR_1\, Q
         => \REG[472]\);
    
    SOFT_PON_GENERATE_P_SoftPON_cnt1_4 : MUX2H
      port map(A => I_5_1, B => \cnt1[1]\, S => \un1_stop2_1_0\, 
        Y => cnt1_4);
    
    \SOFT_PON_GENERATE_cnt2[10]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_18, Q => \cnt2[10]\);
    
    cnt2_2_0_I_45 : XOR2
      port map(A => N_131, B => \cnt2[8]\, Y => \cnt2_2[8]\);
    
    SOFT_PON_GENERATE_cnt2_35 : MUX2H
      port map(A => \cnt2_2[27]\, B => \cnt2[27]\, S => stop2_0, 
        Y => cnt2_35);
    
    cnt2_2_0_I_173 : XOR2
      port map(A => N_40, B => \cnt2[25]\, Y => \cnt2_2_i_i[25]\);
    
    SOFT_PON_GENERATE_cnt2_27 : MUX2H
      port map(A => \cnt2_2_i_i[19]\, B => \cnt2[19]\, S => 
        stop2_1, Y => cnt2_27);
    
    SOFT_PON_GENERATE_cnt2_30 : MUX2H
      port map(A => \cnt2_2[22]\, B => \cnt2[22]\, S => stop2_1, 
        Y => cnt2_30);
    
    TCNT2_2_I_36 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    cnt2_2_0_I_156 : XOR2
      port map(A => N_52, B => \cnt2[23]\, Y => \cnt2_2_i_i[23]\);
    
    TCNT3_2_I_31 : XOR2
      port map(A => \TCNT3[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP_0[0]\, Y => \TCNT3_2[1]\);
    
    HWRES_22 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_22);
    
    \SOFT_PON_GENERATE_P_SoftPON_cnt1[0]\ : DFF
      port map(CLK => CLK_c_c, D => cnt1_3, Q => \cnt1[0]\);
    
    \SOFT_PON_GENERATE_cnt2[26]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_34, Q => \cnt2[26]\);
    
    EV_RES1 : DFFC
      port map(CLK => ALICLK_c, D => EVRES_c, CLR => un8_hwresi_i, 
        Q => \EV_RES1\);
    
    HWRES_34 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_34);
    
    un3_activity_I_77 : XOR2
      port map(A => N_14_0, B => \REG[470]\, Y => I_77);
    
    HWRES_6 : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        HWRES_c_6);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i : OR3
      port map(A => un7_stop2_i_29_i, B => un7_stop2_i_25_i, C
         => un7_stop2_i_24_i, Y => un7_stop2_i);
    
    HWRES_c_i : INV
      port map(A => \HWRES_c_3\, Y => HWRES_c_i_0);
    
    cnt2_2_0_I_23 : AND3
      port map(A => \DWACT_FINC_E_0[0]\, B => \cnt2[3]\, C => 
        \cnt2[4]\, Y => N_146);
    
    HWRES_4 : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        HWRES_c_4);
    
    cnt2_2_0_I_166 : XOR2
      port map(A => N_45, B => \cnt2[24]\, Y => \cnt2_2[24]\);
    
    \CLEAR_3\ : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => CLEAR_3);
    
    un3_activity_I_59 : AND3
      port map(A => \REG[463]\, B => \REG[464]\, C => \REG[465]\, 
        Y => \DWACT_FINC_E_0[5]\);
    
    \CLEAR_13\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_13);
    
    \ACTIVITY[2]\ : DFFC
      port map(CLK => ALICLK_c, D => I_9, CLR => \CLEAR_1\, Q => 
        \REG[459]\);
    
    un1_tcnt1_I_4 : INV
      port map(A => \TCNT1[0]_net_1\, Y => I_4_0);
    
    \CLEAR_23\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_23);
    
    cnt2_2_0_I_20 : XOR2
      port map(A => N_149, B => \cnt2[4]\, Y => \cnt2_2[4]\);
    
    cnt2_2_0_I_104 : AND3
      port map(A => \DWACT_FINC_E_0[6]\, B => \DWACT_FINC_E[10]\, 
        C => \DWACT_FINC_E[11]\, Y => N_88);
    
    HWRES_21 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_21);
    
    un3_activity_I_30 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E_0[1]\, 
        C => \REG[462]\, Y => N_47);
    
    un1_tcnt1_I_9 : XOR2
      port map(A => N_15, B => \TCNT1_i_i[2]\, Y => I_9_0);
    
    SoftPON : DFF
      port map(CLK => CLK_c_c, D => \SoftPON_2_0\, Q => 
        \TST_c[14]\);
    
    un2_hwresi_2 : OR2
      port map(A => REG_0, B => SYSRESB_c, Y => N_259_2);
    
    \SOFT_PON_GENERATE_cnt2[22]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_30, Q => \cnt2[22]\);
    
    cnt2_2_0_I_135 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[15]\, Y => N_66);
    
    TCNT3_2_I_42 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \TCNT3_i_i[4]\, Y => \DWACT_ADD_CI_0_g_array_12_1_0[0]\);
    
    LongSoftPON_3 : DFF
      port map(CLK => CLK_c_c, D => LongSoftPON_1_i, Q => 
        \TST_c_3[15]\);
    
    SOFT_PON_GENERATE_cnt2_31 : MUX2H
      port map(A => \cnt2_2_i_i[23]\, B => \cnt2[23]\, S => 
        stop2_1, Y => cnt2_31);
    
    cnt2_2_0_I_59 : AND3
      port map(A => \cnt2[6]\, B => \cnt2[7]\, C => \cnt2[8]\, Y
         => \DWACT_FINC_E[5]\);
    
    cnt2_2_0_I_122 : XOR2
      port map(A => N_76, B => \cnt2[19]\, Y => \cnt2_2_i_i[19]\);
    
    un3_activity_I_19 : AND2
      port map(A => \REG[460]\, B => \DWACT_FINC_E[0]\, Y => N_55);
    
    un15_tcnt4_0_a3_0 : OR2
      port map(A => \TCNT4_i_0_i[2]\, B => \TCNT4[3]_net_1\, Y
         => un15_tcnt4_0_a3_0_i);
    
    cnt2_2_0_I_13 : XOR2
      port map(A => N_154, B => \cnt2[3]\, Y => \cnt2_2[3]\);
    
    cnt2_2_0_I_105 : XOR2
      port map(A => N_88, B => \cnt2[17]\, Y => \cnt2_2[17]\);
    
    cnt2_2_0_I_27 : AND2
      port map(A => \cnt2[3]\, B => \cnt2[4]\, Y => 
        \DWACT_FINC_E[1]\);
    
    cnt2_2_0_I_202 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \cnt2[27]\, Y => N_19);
    
    SOFT_PON_GENERATE_cnt2_37 : MUX2H
      port map(A => \cnt2_2_i_i[29]\, B => \cnt2[29]\, S => 
        stop2_0, Y => cnt2_37);
    
    HWRES_10 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_10);
    
    TCNT3_2_I_47 : AND2
      port map(A => \TCNT3_i_i[2]\, B => \TCNT3[3]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\);
    
    cnt2_2_0_I_31 : XOR2
      port map(A => N_141, B => \cnt2[6]\, Y => \cnt2_2[6]\);
    
    cnt2_2_0_I_203 : XOR2
      port map(A => N_19, B => \cnt2[28]\, Y => \cnt2_2[28]\);
    
    un11_tcnt3_i_0_0 : OR2
      port map(A => \TCNT3_i_i[6]\, B => \TCNT3[7]_net_1\, Y => 
        un11_tcnt3_i_0_0_i);
    
    SoftPON_2_0_a3_0 : NAND3
      port map(A => un7_stop2_i, B => \TST_c[14]\, C => stop1, Y
         => \SoftPON_2_0_a3_0\);
    
    HWRES_1 : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        HWRES_c_1);
    
    TCNT2_2_I_48 : AND2
      port map(A => \TCNT2_i_i[4]\, B => \TCNT2[5]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    HWRES_0 : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        \HWRES_c_0\);
    
    \SOFT_PON_GENERATE_cnt2[31]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_39, Q => \cnt2[31]\);
    
    TCNT3_2_I_44 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_0[0]\, B => 
        \TCNT3_i_i[2]\, Y => \DWACT_ADD_CI_0_g_array_12_0[0]\);
    
    HWRES_0_5 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_0_5);
    
    cnt2_2_0_I_48 : AND3
      port map(A => \DWACT_FINC_E_0[0]\, B => \DWACT_FINC_E[2]\, 
        C => \DWACT_FINC_E[3]\, Y => \DWACT_FINC_E_0[4]\);
    
    TCNT3_2_I_35 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_0[0]\, B => 
        \TCNT3[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1_0[0]\);
    
    HWRES_32 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_32);
    
    un11_tcnt3_i_0_4 : OR3
      port map(A => un11_tcnt3_i_0_2_i, B => \TCNT3_i_i[0]\, C
         => \TCNT3[1]_net_1\, Y => un11_tcnt3_i_0_4_i);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_25 : NAND3FTT
      port map(A => \cnt2_2[17]\, B => un7_stop2_i_19, C => 
        \cnt2_2[11]\, Y => un7_stop2_i_25_i);
    
    cnt2_2_0_I_90 : AND3
      port map(A => \DWACT_FINC_E_0[6]\, B => \DWACT_FINC_E_0[7]\, 
        C => \DWACT_FINC_E[9]\, Y => N_98);
    
    \SOFT_PON_GENERATE_cnt2[17]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_25, Q => \cnt2[17]\);
    
    BNC_RESi : DFFC
      port map(CLK => ALICLK_c, D => \BNC_RESi_1\, CLR => 
        un8_hwresi_i, Q => LBSP_c(2));
    
    TCNT3_2_I_1 : AND2
      port map(A => \TCNT3_i_i[0]\, B => \TICK[1]\, Y => 
        \DWACT_ADD_CI_0_TMP_0[0]\);
    
    stop_0_sqmuxa_i : INV
      port map(A => \stop_0_sqmuxa\, Y => \stop_0_sqmuxa_i\);
    
    LongSoftPON_2 : DFF
      port map(CLK => CLK_c_c, D => LongSoftPON_1_i, Q => 
        \TST_c_2[15]\);
    
    un2_hwresi_3 : OR2
      port map(A => REG_0, B => SYSRESB_c, Y => N_259_3);
    
    SoftPON_2_0_a3 : OR3FFT
      port map(A => un3_stop2_i, B => un7_stop2_i, C => stop1, Y
         => \SoftPON_2_0_a3\);
    
    un11_tcnt3_i_0 : OR3
      port map(A => un11_tcnt3_i_0_4_i, B => un11_tcnt3_i_0_0_i, 
        C => un11_tcnt3_i_0_1_i, Y => \un11_tcnt3_i_0\);
    
    un3_activity_I_62 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E_0[2]\, 
        C => \DWACT_FINC_E_0[5]\, Y => \DWACT_FINC_E[6]\);
    
    un1_tcnt1_I_8 : AND2
      port map(A => \TCNT1_i_i[1]\, B => \TCNT1[0]_net_1\, Y => 
        N_15);
    
    \ACTIVITY[3]\ : DFFC
      port map(CLK => ALICLK_c, D => I_13_0, CLR => \CLEAR_1\, Q
         => \REG[460]\);
    
    un1_cnt1_1_I_13 : XOR2
      port map(A => N_4_0, B => \cnt1[3]\, Y => I_13_2);
    
    GND_i : GND
      port map(Y => \GND\);
    
    cnt2_2_0_I_186 : XOR2
      port map(A => N_31, B => \cnt2[26]\, Y => \cnt2_2[26]\);
    
    HWRES_10_0 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_10_0);
    
    \ACTIVITY[0]\ : DFFC
      port map(CLK => ALICLK_c, D => I_4, CLR => \CLEAR_1\, Q => 
        \REG[457]\);
    
    un3_activity_I_45 : XOR2
      port map(A => N_37, B => \REG[465]\, Y => I_45);
    
    un3_activity_I_24 : XOR2
      port map(A => N_52_0, B => \REG[462]\, Y => I_24);
    
    \TCNT1[2]\ : DFF
      port map(CLK => CLK_c_c, D => I_9_0, Q => \TCNT1_i_i[2]\);
    
    HWRES_23 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_23);
    
    \CLEAR_9\ : OR3FTT
      port map(A => LOAD_RES_2, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_9);
    
    \CLEAR_16\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_16);
    
    un11_tcnt3_i_0_2 : OR2
      port map(A => \TCNT3_i_i[2]\, B => \TCNT3[3]_net_1\, Y => 
        un11_tcnt3_i_0_2_i);
    
    HWRES_31 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_31);
    
    cnt2_2_0_I_129 : XOR2
      port map(A => N_71, B => \cnt2[20]\, Y => \cnt2_2[20]\);
    
    cnt2_2_0_I_72 : AND2
      port map(A => \DWACT_FINC_E_0[7]\, B => \DWACT_FINC_E_0[6]\, 
        Y => N_111);
    
    \CLEAR_26\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_26);
    
    cnt2_2_0_I_152 : AND3
      port map(A => \DWACT_FINC_E[34]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[5]\, Y => \DWACT_FINC_E[29]\);
    
    un15_tcnt4_0_a3_i : INV
      port map(A => \un10_tcnt2_i_o3\, Y => N_270_i_0);
    
    cnt2_2_0_I_97 : AND3
      port map(A => \DWACT_FINC_E_0[6]\, B => \DWACT_FINC_E[10]\, 
        C => \cnt2[15]\, Y => N_93);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_20 : OR3
      port map(A => un7_stop2_i_12_i, B => \cnt2_2_i_i[19]\, C
         => \cnt2_2[20]\, Y => un7_stop2_i_20_i);
    
    TCNT3_2_I_27 : XOR2
      port map(A => \TCNT3_i_i[6]\, B => 
        \DWACT_ADD_CI_0_g_array_11_0[0]\, Y => \TCNT3_2[6]\);
    
    \TCNT3[4]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT3_2[4]\, Q => 
        \TCNT3_i_i[4]\);
    
    HWRES_13_0 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_13_0);
    
    cnt2_2_0_I_162 : AND2
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        Y => \DWACT_FINC_E[18]\);
    
    \ACTIVITY[1]\ : DFFC
      port map(CLK => ALICLK_c, D => I_5, CLR => \CLEAR_1\, Q => 
        \REG[458]\);
    
    SOFT_PON_GENERATE_P_SoftPON_LongSoftPON_1_i : AND2
      port map(A => \TST_c[13]\, B => \TST_c[14]\, Y => 
        LongSoftPON_1_i);
    
    BNC_RES1 : DFFC
      port map(CLK => ALICLK_c, D => BNCRES_c, CLR => 
        un8_hwresi_i, Q => \BNC_RES1\);
    
    \TICKi_2[0]\ : DFF
      port map(CLK => CLK_c_c, D => N_269_i_0, Q => TICK_2(0));
    
    SOFT_PON_GENERATE_cnt2_9 : MUX2H
      port map(A => \cnt2_2[1]\, B => \cnt2[1]_net_1\, S => stop2, 
        Y => cnt2_9);
    
    CLEAR_i : INV
      port map(A => CLEAR_0_net_1, Y => CLEAR_i_0);
    
    \ACTIVITY[14]\ : DFFC
      port map(CLK => ALICLK_c, D => I_84, CLR => \CLEAR_1\, Q
         => \REG[471]\);
    
    \ACTIVITY[13]\ : DFFC
      port map(CLK => ALICLK_c, D => I_77, CLR => \CLEAR_1\, Q
         => \REG[470]\);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_21 : OR3
      port map(A => \cnt2_2_i_i[31]\, B => un7_stop2_i_8_i, C => 
        \cnt2_2[18]\, Y => un7_stop2_i_21_i);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_2 : NAND3FTT
      port map(A => \cnt2[0]_net_1\, B => un7_stop2_i_1, C => 
        \cnt2_2[1]\, Y => un7_stop2_i_2_i);
    
    \TCNT4[1]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT4_2[1]\, Q => 
        \TCNT4[1]_net_1\);
    
    TCNT3_2_I_33 : XOR2
      port map(A => \TCNT3[5]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_1_0[0]\, Y => \TCNT3_2[5]\);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_4 : AND2
      port map(A => \cnt2_2[6]\, B => \cnt2_2[7]\, Y => 
        un7_stop2_i_4);
    
    \SOFT_PON_GENERATE_cnt2[28]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_36, Q => \cnt2[28]\);
    
    \cnt2[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \cnt2_1\, CLR => \HWRES_c_3\, 
        Q => \cnt2_0[0]\);
    
    CLEAR_0_1 : NAND2
      port map(A => \NLBCLR_c\, B => RUN_c_0_0, Y => CLEAR_0_i_1);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_29 : OR3
      port map(A => un7_stop2_i_26_i, B => un7_stop2_i_23_i, C
         => un7_stop2_i_21_i, Y => un7_stop2_i_29_i);
    
    un1_cnt1_1_I_9 : XOR2
      port map(A => N_7, B => \cnt1[2]\, Y => I_9_1);
    
    \ACTIVITY[11]\ : DFFC
      port map(CLK => ALICLK_c, D => I_66, CLR => \CLEAR_1\, Q
         => \REG[468]\);
    
    un10_tcnt2_i_o3_4 : OR3
      port map(A => un10_tcnt2_i_o3_2_i, B => \TCNT2_i_i[0]\, C
         => \TCNT2[1]_net_1\, Y => un10_tcnt2_i_o3_4_i);
    
    cnt2_2_0_I_4 : INV
      port map(A => \cnt2[0]_net_1\, Y => \cnt2_2[0]\);
    
    un10_tcnt2_i_o3_0 : OR2
      port map(A => \TCNT2_i_i[6]\, B => \TCNT2[7]_net_1\, Y => 
        un10_tcnt2_i_o3_0_i);
    
    un3_activity_I_56 : XOR2
      port map(A => N_29, B => \REG[467]\, Y => I_56);
    
    SOFT_PON_GENERATE_cnt2_18 : MUX2H
      port map(A => \cnt2_2[10]\, B => \cnt2[10]\, S => stop2, Y
         => cnt2_18);
    
    \SOFT_PON_GENERATE_cnt2[21]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_29, Q => \cnt2[21]\);
    
    \TCNT3[1]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT3_2[1]\, Q => 
        \TCNT3[1]_net_1\);
    
    SOFT_PON_GENERATE_P_SoftPON_cnt1_6 : MUX2H
      port map(A => I_13_2, B => \cnt1[3]\, S => \un1_stop2_1_0\, 
        Y => cnt1_6);
    
    SOFT_PON_GENERATE_P_SoftPON_stop1_1_0 : OAI21TTF
      port map(A => stop2_0, B => un3_stop2_i, C => stop1, Y => 
        stop1_1_0);
    
    SOFT_PON_GENERATE_cnt2_13 : MUX2H
      port map(A => \cnt2_2[5]\, B => \cnt2[5]\, S => stop2, Y
         => cnt2_13);
    
    TCNT2_2_I_19 : XOR2
      port map(A => \TCNT2_i_i[0]\, B => \TICK[0]\, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    HWRES : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        HWRES_c);
    
    cnt2_2_0_I_159 : AND3
      port map(A => \cnt2[21]\, B => \cnt2[22]\, C => \cnt2[23]\, 
        Y => \DWACT_FINC_E[17]\);
    
    un3_activity_I_23 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \REG[460]\, C => 
        \REG[461]\, Y => N_52_0);
    
    un1_tcnt1_I_5 : XOR2
      port map(A => \TCNT1[0]_net_1\, B => \TCNT1_i_i[1]\, Y => 
        I_5_0);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_8 : NAND2FT
      port map(A => \cnt2_2[27]\, B => \cnt2_2[9]\, Y => 
        un7_stop2_i_8_i);
    
    \SOFT_PON_GENERATE_cnt2[24]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_32, Q => \cnt2[24]\);
    
    \SOFT_PON_GENERATE_P_SoftPON_cnt1[1]\ : DFF
      port map(CLK => CLK_c_c, D => cnt1_4, Q => \cnt1[1]\);
    
    TCNT2_2_I_30 : XOR2
      port map(A => \TCNT2[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => \TCNT2_2[3]\);
    
    \SOFT_PON_GENERATE_cnt2[29]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_37, Q => \cnt2[29]\);
    
    cnt2_2_0_I_220 : AND2
      port map(A => \DWACT_FINC_E[26]\, B => \cnt2[30]\, Y => 
        \DWACT_FINC_E[27]\);
    
    un4_ticki : AND2FT
      port map(A => \stop\, B => \TICK[3]\, Y => \un4_ticki\);
    
    cnt2_2_0_I_38 : XOR2
      port map(A => N_136, B => \cnt2[7]\, Y => \cnt2_2[7]\);
    
    cnt2_2_0_I_169 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        C => \cnt2[24]\, Y => \DWACT_FINC_E[19]\);
    
    cnt2_2_0_I_83 : AND3
      port map(A => \DWACT_FINC_E_0[6]\, B => \DWACT_FINC_E_0[7]\, 
        C => \DWACT_FINC_E[8]\, Y => N_103);
    
    cnt2_2_0_I_76 : AND3
      port map(A => \DWACT_FINC_E_0[6]\, B => \DWACT_FINC_E_0[7]\, 
        C => \cnt2[12]\, Y => N_108);
    
    \CLEAR_4\ : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => CLEAR_4);
    
    \SOFT_PON_GENERATE_cnt2[5]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_13, Q => \cnt2[5]\);
    
    PON_LOAD : DFFS
      port map(CLK => CLK_c_c, D => \stop_0_sqmuxa_i\, SET => 
        \HWRES_c_3\, Q => PON_LOAD_i);
    
    un1_stop2_1_0 : OR2
      port map(A => stop2_0, B => stop1, Y => \un1_stop2_1_0\);
    
    HWRES_33 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_33);
    
    HWRES_7 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_7);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \TCNT2[2]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT2_2[2]\, Q => 
        \TCNT2_i_i[2]\);
    
    cnt2_2_0_I_80 : AND2
      port map(A => \cnt2[12]\, B => \cnt2[13]\, Y => 
        \DWACT_FINC_E[8]\);
    
    cnt2_2_0_I_44 : AND3
      port map(A => \DWACT_FINC_E_0[0]\, B => \DWACT_FINC_E[2]\, 
        C => \DWACT_FINC_E[3]\, Y => N_131);
    
    un3_activity_I_16 : AND3
      port map(A => \REG[457]\, B => \REG[458]\, C => \REG[459]\, 
        Y => \DWACT_FINC_E[0]\);
    
    HWRES_20 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_20);
    
    HWRES_2 : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        HWRES_c_2);
    
    SOFT_PON_GENERATE_cnt2_28 : MUX2H
      port map(A => \cnt2_2[20]\, B => \cnt2[20]\, S => stop2_1, 
        Y => cnt2_28);
    
    un15_tcnt4_0_a3 : NOR3
      port map(A => \un10_tcnt2_i_o3\, B => \un11_tcnt3_i_0\, C
         => un15_tcnt4_0_a3_2_i, Y => \un15_tcnt4_0_a3\);
    
    \TICKi_0[0]\ : DFF
      port map(CLK => CLK_c_c, D => N_269_i_0, Q => TICK_0_0);
    
    \TCNT4[0]\ : DFF
      port map(CLK => CLK_c_c, D => 
        \DWACT_ADD_CI_0_partial_sum_1[0]\, Q => \TCNT4_i_0_i[0]\);
    
    TCNT2_2_I_27 : XOR2
      port map(A => \TCNT2_i_i[6]\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => \TCNT2_2[6]\);
    
    \SOFT_PON_GENERATE_cnt2[4]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_12, Q => \cnt2[4]\);
    
    un1_tcnt1_I_20 : XOR2
      port map(A => N_7_0, B => \TCNT1_i_i[4]\, Y => I_20_0);
    
    cnt2_2_0_I_182 : AND3
      port map(A => \DWACT_FINC_E_0[7]\, B => \DWACT_FINC_E[9]\, 
        C => \DWACT_FINC_E[12]\, Y => \DWACT_FINC_E[30]\);
    
    SOFT_PON_GENERATE_cnt2_23 : MUX2H
      port map(A => \cnt2_2_i_i[15]\, B => \cnt2[15]\, S => 
        stop2_1, Y => cnt2_23);
    
    HWRES_5 : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        HWRES_c_5);
    
    \SOFT_PON_GENERATE_cnt2[15]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_23, Q => \cnt2[15]\);
    
    cnt2_2_0_I_146 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \cnt2[21]\, C => 
        \cnt2[22]\, Y => \DWACT_FINC_E[33]\);
    
    \SOFT_PON_GENERATE_P_SoftPON_cnt1[3]\ : DFF
      port map(CLK => CLK_c_c, D => cnt1_6, Q => \cnt1[3]\);
    
    LongSoftPON : DFF
      port map(CLK => CLK_c_c, D => LongSoftPON_1_i, Q => 
        \TST_c[15]\);
    
    cnt2_2_0_I_206 : AND2
      port map(A => \cnt2[27]\, B => \cnt2[28]\, Y => 
        \DWACT_FINC_E[25]\);
    
    un10_tcnt2_i_o3_i : NOR3
      port map(A => un6_tcnt1_i_0_2_i, B => un6_tcnt1_i_0_1_i, C
         => \TCNT1[0]_net_1\, Y => N_269_i_0);
    
    un1_tcnt1_I_13 : XOR2
      port map(A => N_12, B => \TCNT1[3]_net_1\, Y => I_13_1);
    
    un1_tcnt1_I_23 : AND3
      port map(A => \DWACT_FINC_E_1[0]\, B => \TCNT1[3]_net_1\, C
         => \TCNT1_i_i[4]\, Y => N_4);
    
    cnt2_2_0_I_210 : XOR2
      port map(A => N_14, B => \cnt2[29]\, Y => \cnt2_2_i_i[29]\);
    
    cnt2_2_0_I_125 : AND2
      port map(A => \cnt2[18]\, B => \cnt2[19]\, Y => 
        \DWACT_FINC_E[14]\);
    
    \SOFT_PON_GENERATE_cnt2[7]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_15, Q => \cnt2[7]\);
    
    TCNT2_2_I_32 : XOR2
      port map(A => \TCNT2_i_i[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => \TCNT2_2[2]\);
    
    \SOFT_PON_GENERATE_cnt2[30]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_38, Q => \cnt2[30]\);
    
    \ACTIVITY[6]\ : DFFC
      port map(CLK => ALICLK_c, D => I_31, CLR => CLEAR_2_net_1, 
        Q => \REG[463]\);
    
    TCNT4_2_I_17 : XOR2
      port map(A => \TCNT4[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, Y => \TCNT4_2[3]\);
    
    cnt2_2_0_I_87 : AND3
      port map(A => \cnt2[12]\, B => \cnt2[13]\, C => \cnt2[14]\, 
        Y => \DWACT_FINC_E[9]\);
    
    cnt2_2_0_I_223 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \DWACT_FINC_E[27]\, Y => N_4_1);
    
    BNC_RESi_1 : AND2FT
      port map(A => \BNC_RES1\, B => BNCRES_c, Y => \BNC_RESi_1\);
    
    \TCNT4[3]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT4_2[3]\, Q => 
        \TCNT4[3]_net_1\);
    
    cnt2_2_0_I_114 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[10]\, 
        C => \DWACT_FINC_E[12]\, Y => N_81);
    
    cnt2_2_0_I_12 : AND3
      port map(A => \cnt2[0]_net_1\, B => \cnt2[1]_net_1\, C => 
        \cnt2[2]\, Y => N_154);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_7 : NAND3FTT
      port map(A => un7_stop2_i_2_i, B => \cnt2_2[10]\, C => 
        \cnt2_2[8]\, Y => un7_stop2_i_7_i);
    
    cnt2_2_0_I_196 : XOR2
      port map(A => N_24, B => \cnt2[27]\, Y => \cnt2_2[27]\);
    
    TCNT3_2_I_45 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11_0[0]\, B => 
        \TCNT3_i_i[6]\, Y => \DWACT_ADD_CI_0_g_array_12_2_0[0]\);
    
    \SOFT_PON_GENERATE_cnt2[23]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_31, Q => \cnt2[23]\);
    
    cnt2_2_0_I_62 : AND3
      port map(A => \DWACT_FINC_E_0[0]\, B => \DWACT_FINC_E[2]\, 
        C => \DWACT_FINC_E[5]\, Y => \DWACT_FINC_E_0[6]\);
    
    HWRES_18 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_18);
    
    un1_cnt1_1_I_5 : XOR2
      port map(A => \cnt1[0]\, B => \cnt1[1]\, Y => I_5_1);
    
    TCNT2_2_I_34 : XOR2
      port map(A => \TCNT2[7]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => \TCNT2_2[7]\);
    
    SOFT_PON_GENERATE_cnt2_14 : MUX2H
      port map(A => \cnt2_2[6]\, B => \cnt2[6]\, S => stop2, Y
         => cnt2_14);
    
    un3_activity_I_27 : AND2
      port map(A => \REG[460]\, B => \REG[461]\, Y => 
        \DWACT_FINC_E_0[1]\);
    
    HWRES_0_3 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_0_3);
    
    cnt2_2_0_I_189 : AND3
      port map(A => \cnt2[24]\, B => \cnt2[25]\, C => \cnt2[26]\, 
        Y => \DWACT_FINC_E[22]\);
    
    un3_activity_I_9 : XOR2
      port map(A => N_63, B => \REG[459]\, Y => I_9);
    
    cnt2_2_0_I_115 : XOR2
      port map(A => N_81, B => \cnt2[18]\, Y => \cnt2_2[18]\);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_10 : OR2
      port map(A => \cnt2_2_i_i[23]\, B => \cnt2_2[24]\, Y => 
        un7_stop2_i_10_i);
    
    un3_activity_I_8 : AND2
      port map(A => \REG[458]\, B => \REG[457]\, Y => N_63);
    
    SOFT_PON_GENERATE_cnt2_38 : MUX2H
      port map(A => \cnt2_2[30]\, B => \cnt2[30]\, S => stop2_0, 
        Y => cnt2_38);
    
    un3_activity_I_52 : XOR2
      port map(A => N_32, B => \REG[466]\, Y => I_52);
    
    \TCNT2[0]\ : DFF
      port map(CLK => CLK_c_c, D => 
        \DWACT_ADD_CI_0_partial_sum[0]\, Q => \TCNT2_i_i[0]\);
    
    cnt2_2_0_I_213 : AND3
      port map(A => \cnt2[27]\, B => \cnt2[28]\, C => \cnt2[29]\, 
        Y => \DWACT_FINC_E[26]\);
    
    cnt2_2_0_I_209 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \DWACT_FINC_E[25]\, Y => N_14);
    
    HWRES_30 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_30);
    
    SOFT_PON_GENERATE_cnt2_33 : MUX2H
      port map(A => \cnt2_2_i_i[25]\, B => \cnt2[25]\, S => 
        stop2_0, Y => cnt2_33);
    
    SOFT_PON_GENERATE_P_SoftPON_stop2_0 : DFF
      port map(CLK => CLK_c_c, D => stop2_40_i_a3, Q => stop2_0);
    
    SOFT_PON_GENERATE_cnt2_12 : MUX2H
      port map(A => \cnt2_2[4]\, B => \cnt2[4]\, S => stop2, Y
         => cnt2_12);
    
    HWRES_3 : NAND3
      port map(A => N_259, B => NPWON_c, C => \TST_c[15]\, Y => 
        \HWRES_c_3\);
    
    HWCLEARi_2 : NOR2
      port map(A => PULSE(1), B => WDOGTO, Y => \HWCLEARi_2\);
    
    cnt2_2_0_I_155 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[33]\, Y => N_52);
    
    un3_activity_I_5 : XOR2
      port map(A => \REG[457]\, B => \REG[458]\, Y => I_5);
    
    EV_RESi_i : OR2FT
      port map(A => RUN_c_0, B => \HWRES_c_0\, Y => un8_hwresi_i);
    
    \CLEAR_0\ : NAND2
      port map(A => \NLBCLR_c\, B => RUN_c, Y => CLEAR_0_i);
    
    un2_hwresi_1 : OR2
      port map(A => REG_0, B => SYSRESB_c, Y => N_259_1);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_1 : AND2
      port map(A => \cnt2_2[2]\, B => \cnt2_2[3]\, Y => 
        un7_stop2_i_1);
    
    SOFT_PON_GENERATE_P_SoftPON_stop1 : DFF
      port map(CLK => CLK_c_c, D => stop1_1_0, Q => stop1);
    
    un1_tcnt1_I_24 : XOR2
      port map(A => N_4, B => \TCNT1[5]_net_1\, Y => I_24_0);
    
    un1_cnt1_1_I_12 : AND3
      port map(A => \cnt1[0]\, B => \cnt1[1]\, C => \cnt1[2]\, Y
         => N_4_0);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_17 : OR2
      port map(A => \cnt2_2_i_i[15]\, B => \cnt2_2[16]\, Y => 
        un7_stop2_i_17_i);
    
    HWRES_16 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_16);
    
    cnt2_2_0_I_91 : XOR2
      port map(A => N_98, B => \cnt2[15]\, Y => \cnt2_2_i_i[15]\);
    
    cnt2_2_0_I_34 : AND3
      port map(A => \cnt2[3]\, B => \cnt2[4]\, C => \cnt2[5]\, Y
         => \DWACT_FINC_E[2]\);
    
    un3_activity_I_91 : XOR2
      port map(A => N_4_2, B => \REG[472]\, Y => I_91);
    
    \SOFT_PON_GENERATE_cnt2[0]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_8, Q => \cnt2[0]_net_1\);
    
    cnt2_2_0_I_165 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[18]\, Y => N_45);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_19 : NOR3
      port map(A => un7_stop2_i_7_i, B => un7_stop2_i_6_i, C => 
        \cnt2_2[12]\, Y => un7_stop2_i_19);
    
    \TCNT1[5]\ : DFF
      port map(CLK => CLK_c_c, D => I_24_0, Q => \TCNT1[5]_net_1\);
    
    SOFT_PON_GENERATE_cnt2_24 : MUX2H
      port map(A => \cnt2_2[16]\, B => \cnt2[16]\, S => stop2_1, 
        Y => cnt2_24);
    
    cnt2_2_0_I_108 : AND3
      port map(A => \cnt2[15]\, B => \cnt2[16]\, C => \cnt2[17]\, 
        Y => \DWACT_FINC_E[12]\);
    
    \ACTIVITY[8]\ : DFFC
      port map(CLK => ALICLK_c, D => I_45, CLR => CLEAR_2_net_1, 
        Q => \REG[465]\);
    
    TCNT3_2_I_39 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_0[0]\);
    
    \TCNT1[3]\ : DFF
      port map(CLK => CLK_c_c, D => I_13_1, Q => \TCNT1[3]_net_1\);
    
    cnt2_2_0_I_16 : AND3
      port map(A => \cnt2[0]_net_1\, B => \cnt2[1]_net_1\, C => 
        \cnt2[2]\, Y => \DWACT_FINC_E_0[0]\);
    
    HWRES_9 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_9);
    
    cnt2_2_0_I_65 : AND3
      port map(A => \DWACT_FINC_E_0[6]\, B => \cnt2[9]\, C => 
        \cnt2[10]\, Y => N_116);
    
    \SOFT_PON_GENERATE_cnt2[20]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_28, Q => \cnt2[20]\);
    
    un3_activity_I_51 : AND2
      port map(A => \REG[465]\, B => \DWACT_FINC_E[4]\, Y => N_32);
    
    un3_activity_I_12 : AND3
      port map(A => \REG[457]\, B => \REG[458]\, C => \REG[459]\, 
        Y => N_60);
    
    un3_activity_I_76 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[7]\, C
         => \REG[469]\, Y => N_14_0);
    
    HWRES_0_6 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_0_6);
    
    un3_activity_I_20 : XOR2
      port map(A => N_55, B => \REG[461]\, Y => I_20);
    
    cnt2_2_0_I_66 : XOR2
      port map(A => N_116, B => \cnt2[11]\, Y => \cnt2_2[11]\);
    
    cnt2_2_0_I_142 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[16]\, Y => N_61);
    
    TCNT4_2_I_11 : XOR2
      port map(A => \TCNT4_i_0_i[0]\, B => \TICK[2]\, Y => 
        \DWACT_ADD_CI_0_partial_sum_1[0]\);
    
    TCNT3_2_I_36 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\);
    
    SOFT_PON_GENERATE_cnt2_22 : MUX2H
      port map(A => \cnt2_2[14]\, B => \cnt2[14]\, S => stop2_1, 
        Y => cnt2_22);
    
    \TICKi[3]\ : DFF
      port map(CLK => CLK_c_c, D => \un15_tcnt4_0_a3\, Q => 
        \TICK[3]\);
    
    \TICKi[1]\ : DFF
      port map(CLK => CLK_c_c, D => N_270_i_0, Q => \TICK[1]\);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_9 : OR2
      port map(A => \cnt2_2_i_i[25]\, B => \cnt2_2[26]\, Y => 
        un7_stop2_i_9_i);
    
    \SOFT_PON_GENERATE_cnt2[6]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_14, Q => \cnt2[6]\);
    
    \ACTIVITY[7]\ : DFFC
      port map(CLK => ALICLK_c, D => I_38, CLR => CLEAR_2_net_1, 
        Q => \REG[464]\);
    
    HWRES_22_0 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_22_0);
    
    \ACTIVITY[5]\ : DFFC
      port map(CLK => ALICLK_c, D => I_24, CLR => \CLEAR_1\, Q
         => \REG[462]\);
    
    TCNT2_2_I_31 : XOR2
      port map(A => \TCNT2[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => \TCNT2_2[1]\);
    
    \SOFT_PON_GENERATE_cnt2[16]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_24, Q => \cnt2[16]\);
    
    CLEAR_1 : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => \CLEAR_1\);
    
    \TCNT2[5]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT2_2[5]\, Q => 
        \TCNT2[5]_net_1\);
    
    un3_activity_I_84 : XOR2
      port map(A => N_9_0, B => \REG[471]\, Y => I_84);
    
    \CLEAR_2\ : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => CLEAR_2_net_1);
    
    SOFT_PON_GENERATE_cnt2_8 : MUX2H
      port map(A => \cnt2_2[0]\, B => \cnt2[0]_net_1\, S => stop2, 
        Y => cnt2_8);
    
    cnt2_2_0_I_192 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        C => \DWACT_FINC_E[22]\, Y => \DWACT_FINC_E[23]\);
    
    \CLEAR_14\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_14);
    
    TCNT3_2_I_19 : XOR2
      port map(A => \TCNT3_i_i[0]\, B => \TICK[1]\, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\);
    
    \SOFT_PON_GENERATE_cnt2[9]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_17, Q => \cnt2[9]\);
    
    \CLEAR_24\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_24);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_24 : OR3
      port map(A => un7_stop2_i_17_i, B => \cnt2_2_i_i[13]\, C
         => \cnt2_2[14]\, Y => un7_stop2_i_24_i);
    
    SOFT_PON_GENERATE_cnt2_16 : MUX2H
      port map(A => \cnt2_2[8]\, B => \cnt2[8]\, S => stop2, Y
         => cnt2_16);
    
    \TCNT1[1]\ : DFF
      port map(CLK => CLK_c_c, D => I_5_0, Q => \TCNT1_i_i[1]\);
    
    \TCNT2[6]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT2_2[6]\, Q => 
        \TCNT2_i_i[6]\);
    
    TCNT4_2_I_1 : AND2
      port map(A => \TCNT4_i_0_i[0]\, B => \TICK[2]\, Y => 
        \DWACT_ADD_CI_0_TMP_1[0]\);
    
    \TCNT4[2]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT4_2[2]\, Q => 
        \TCNT4_i_0_i[2]\);
    
    SOFT_PON_GENERATE_cnt2_34 : MUX2H
      port map(A => \cnt2_2[26]\, B => \cnt2[26]\, S => stop2_0, 
        Y => cnt2_34);
    
    \TCNT3[2]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT3_2[2]\, Q => 
        \TCNT3_i_i[2]\);
    
    \TCNT3[3]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT3_2[3]\, Q => 
        \TCNT3[3]_net_1\);
    
    \CLEAR_11\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_11);
    
    \TICKi_1[0]\ : DFF
      port map(CLK => CLK_c_c, D => N_269_i_0, Q => TICK_1(0));
    
    cnt2_2_0_I_185 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[30]\, 
        C => \DWACT_FINC_E[21]\, Y => N_31);
    
    cnt2_2_0_I_149 : AND3
      port map(A => \cnt2[0]_net_1\, B => \cnt2[1]_net_1\, C => 
        \cnt2[2]\, Y => \DWACT_FINC_E[34]\);
    
    \SOFT_PON_GENERATE_cnt2[12]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_20, Q => \cnt2[12]\);
    
    EV_RESi_1 : AND2FT
      port map(A => \EV_RES1\, B => EVRES_c, Y => \EV_RESi_1\);
    
    \CLEAR_21\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_21);
    
    HWRES_28 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_28);
    
    HWRES_19 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_19);
    
    cnt2_2_0_I_101 : AND2
      port map(A => \cnt2[15]\, B => \cnt2[16]\, Y => 
        \DWACT_FINC_E[11]\);
    
    \CLEAR_5\ : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => CLEAR_5);
    
    TCNT3_2_I_48 : AND2
      port map(A => \TCNT3_i_i[4]\, B => \TCNT3[5]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1_0[0]\);
    
    un1_tcnt1_I_16 : AND3
      port map(A => \TCNT1[0]_net_1\, B => \TCNT1_i_i[1]\, C => 
        \TCNT1_i_i[2]\, Y => \DWACT_FINC_E_1[0]\);
    
    cnt2_2_0_I_143 : XOR2
      port map(A => N_61, B => \cnt2[22]\, Y => \cnt2_2[22]\);
    
    \cnt2[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \cnt2_2\, CLR => \HWRES_c_3\, 
        Q => \cnt2_0[1]\);
    
    TCNT2_2_I_42 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \TCNT2_i_i[4]\, Y => \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    HWRES_0_0 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => \HWRES_c_0_0\);
    
    SOFT_PON_GENERATE_cnt2_32 : MUX2H
      port map(A => \cnt2_2[24]\, B => \cnt2[24]\, S => stop2_0, 
        Y => cnt2_32);
    
    \SOFT_PON_GENERATE_cnt2[1]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_9, Q => \cnt2[1]_net_1\);
    
    \TCNT3[7]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT3_2[7]\, Q => 
        \TCNT3[7]_net_1\);
    
    \TCNT1[4]\ : DFF
      port map(CLK => CLK_c_c, D => I_20_0, Q => \TCNT1_i_i[4]\);
    
    un1_cnt1_1_I_4 : INV
      port map(A => \cnt1[0]\, Y => I_4_1);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_26 : OR3
      port map(A => un7_stop2_i_20_i, B => \cnt2_2_i_i[29]\, C
         => \cnt2_2[30]\, Y => un7_stop2_i_26_i);
    
    cnt2_2_0_I_199 : AND2
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[30]\, 
        Y => \DWACT_FINC_E[24]\);
    
    TCNT4_2_I_15 : XOR2
      port map(A => \TCNT4[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP_1[0]\, Y => \TCNT4_2[1]\);
    
    SOFT_PON_GENERATE_cnt2_26 : MUX2H
      port map(A => \cnt2_2[18]\, B => \cnt2[18]\, S => stop2_1, 
        Y => cnt2_26);
    
    cnt2_2_0_I_98 : XOR2
      port map(A => N_93, B => \cnt2[16]\, Y => \cnt2_2[16]\);
    
    \CLEAR_19\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_0, Y => CLEAR_19);
    
    HWRES_27_0 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_27_0);
    
    un3_activity_I_83 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[7]\, C
         => \DWACT_FINC_E_0[8]\, Y => N_9_0);
    
    un3_activity_I_4 : INV
      port map(A => \REG[457]\, Y => I_4);
    
    \ACTIVITY[12]\ : DFFC
      port map(CLK => ALICLK_c, D => I_73, CLR => \CLEAR_1\, Q
         => \REG[469]\);
    
    TCNT2_2_I_47 : AND2
      port map(A => \TCNT2_i_i[2]\, B => \TCNT2[3]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    stop_7 : OR2
      port map(A => \stop\, B => \stop_0_sqmuxa\, Y => \stop_7\);
    
    \SOFT_PON_GENERATE_cnt2[27]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_35, Q => \cnt2[27]\);
    
    HWRES_15 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_15);
    
    HWRES_0_1 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_0_1);
    
    \ACTIVITY[10]\ : DFFC
      port map(CLK => ALICLK_c, D => I_56, CLR => \CLEAR_1\, Q
         => \REG[467]\);
    
    cnt2_2_0_I_52 : XOR2
      port map(A => N_126, B => \cnt2[9]\, Y => \cnt2_2[9]\);
    
    \TCNT3[0]\ : DFF
      port map(CLK => CLK_c_c, D => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, Q => \TCNT3_i_i[0]\);
    
    SOFT_PON_GENERATE_P_SoftPON_stop2_40_i_a3 : OR2FT
      port map(A => un7_stop2_i, B => stop2_0, Y => stop2_40_i_a3);
    
    TCNT2_2_I_35 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \TCNT2[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \TCNT2[1]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT2_2[1]\, Q => 
        \TCNT2[1]_net_1\);
    
    \CLEAR_10\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_10);
    
    un3_activity_I_38 : XOR2
      port map(A => N_42, B => \REG[464]\, Y => I_38);
    
    TCNT2_2_I_44 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \TCNT2_i_i[2]\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    cnt2_2_0_I_216 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \DWACT_FINC_E[26]\, Y => N_9);
    
    HWRES_26 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_26);
    
    \CLEAR_20\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_20);
    
    \CLEAR_12\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_12);
    
    cnt2_2_0_I_136 : XOR2
      port map(A => N_66, B => \cnt2[21]\, Y => \cnt2_2_i_i[21]\);
    
    un3_activity_I_48 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E_0[2]\, 
        C => \DWACT_FINC_E_0[3]\, Y => \DWACT_FINC_E[4]\);
    
    un1_tcnt1_I_12 : AND3
      port map(A => \TCNT1[0]_net_1\, B => \TCNT1_i_i[1]\, C => 
        \TCNT1_i_i[2]\, Y => N_12);
    
    \CLEAR_22\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_22);
    
    un3_activity_I_31 : XOR2
      port map(A => N_47, B => \REG[463]\, Y => I_31);
    
    un3_activity_I_72 : AND2
      port map(A => \DWACT_FINC_E[7]\, B => \DWACT_FINC_E[6]\, Y
         => N_17);
    
    SOFT_PON_GENERATE_P_SoftPON_cnt1_3 : MUX2H
      port map(A => I_4_1, B => \cnt1[0]\, S => \un1_stop2_1_0\, 
        Y => cnt1_3);
    
    HWRES_7_0 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_7_0);
    
    un15_tcnt4_0_a3_2 : OR3
      port map(A => un15_tcnt4_0_a3_0_i, B => \TCNT4_i_0_i[0]\, C
         => \TCNT4[1]_net_1\, Y => un15_tcnt4_0_a3_2_i);
    
    un3_activity_I_41 : AND2
      port map(A => \REG[463]\, B => \REG[464]\, Y => 
        \DWACT_FINC_E_0[3]\);
    
    \TICKi_0[2]\ : DFF
      port map(CLK => CLK_c_c, D => \un12_tcnt3_i\, Q => TICK_0_2);
    
    SOFT_PON_GENERATE_P_SoftPON_stop2_1 : DFF
      port map(CLK => CLK_c_c, D => stop2_40_i_a3, Q => stop2_1);
    
    \SOFT_PON_GENERATE_cnt2[2]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_10, Q => \cnt2[2]\);
    
    TCNT3_2_I_28 : XOR2
      port map(A => \TCNT3_i_i[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\, Y => \TCNT3_2[4]\);
    
    \ACTIVITY[9]\ : DFFC
      port map(CLK => ALICLK_c, D => I_52, CLR => CLEAR_2_net_1, 
        Q => \REG[466]\);
    
    stop_0_sqmuxa : AND3FTT
      port map(A => \cnt2_0[1]\, B => \un4_ticki\, C => 
        \cnt2_0[0]\, Y => \stop_0_sqmuxa\);
    
    SoftPON_2_0 : OR3FFT
      port map(A => \SoftPON_2_0_a3_0\, B => \SoftPON_2_0_a3\, C
         => stop2_0, Y => \SoftPON_2_0\);
    
    HWRES_14 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_14);
    
    cnt2_2_0_I_51 : AND2
      port map(A => \cnt2[8]\, B => \DWACT_FINC_E_0[4]\, Y => 
        N_126);
    
    cnt2_2_0_I_24 : XOR2
      port map(A => N_146, B => \cnt2[5]\, Y => \cnt2_2[5]\);
    
    \CLEAR_17\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_17);
    
    un3_activity_I_65 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \REG[466]\, C => 
        \REG[467]\, Y => N_22);
    
    un3_activity_I_13 : XOR2
      port map(A => N_60, B => \REG[460]\, Y => I_13_0);
    
    HWCLEARi : DFFC
      port map(CLK => CLK_c_c, D => \HWCLEARi_2\, CLR => 
        \HWRES_c_3\, Q => \NLBCLR_c\);
    
    HWRES_21_0 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_21_0);
    
    HWRES_17 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_17);
    
    cnt2_2_0_I_128 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[14]\, Y => N_71);
    
    \CLEAR_27\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_27);
    
    SOFT_PON_GENERATE_P_SoftPON_un7_stop2_i_12 : OR2
      port map(A => \cnt2_2_i_i[21]\, B => \cnt2_2[22]\, Y => 
        un7_stop2_i_12_i);
    
    LongSoftPON_0 : DFF
      port map(CLK => CLK_c_c, D => LongSoftPON_1_i, Q => 
        \TST_c_0[15]\);
    
    CLEAR_0_0 : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => CLEAR_0_net_1);
    
    SOFT_PON_GENERATE_cnt2_36 : MUX2H
      port map(A => \cnt2_2[28]\, B => \cnt2[28]\, S => stop2_0, 
        Y => cnt2_36);
    
    \CLEAR_8\ : OR3FTT
      port map(A => LOAD_RES_2, B => HWRES_c_0_1, C => CLEAR_0_i, 
        Y => CLEAR_8);
    
    \CLEAR_6\ : OR3FTT
      port map(A => LOAD_RES_2, B => \HWRES_c_0_2\, C => 
        CLEAR_0_i, Y => CLEAR_6);
    
    cnt2_2_0_I_55 : AND3
      port map(A => \DWACT_FINC_E_0[4]\, B => \cnt2[8]\, C => 
        \cnt2[9]\, Y => N_123);
    
    cnt2_2_0_I_176 : AND2
      port map(A => \cnt2[24]\, B => \cnt2[25]\, Y => 
        \DWACT_FINC_E[20]\);
    
    un3_activity_I_34 : AND3
      port map(A => \REG[460]\, B => \REG[461]\, C => \REG[462]\, 
        Y => \DWACT_FINC_E_0[2]\);
    
    TCNT2_2_I_33 : XOR2
      port map(A => \TCNT2[5]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => \TCNT2_2[5]\);
    
    cnt2_2_0_I_9 : XOR2
      port map(A => N_157, B => \cnt2[2]\, Y => \cnt2_2[2]\);
    
    \SOFT_PON_GENERATE_cnt2[18]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_26, Q => \cnt2[18]\);
    
    un3_activity_I_44 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E_0[2]\, 
        C => \DWACT_FINC_E_0[3]\, Y => N_37);
    
    HWRES_0_6_0 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_0_6_0);
    
    cnt2_2_0_I_56 : XOR2
      port map(A => N_123, B => \cnt2[10]\, Y => \cnt2_2[10]\);
    
    un1_cnt1_1_I_8 : AND2
      port map(A => \cnt1[1]\, B => \cnt1[0]\, Y => N_7);
    
    CLEAR_0_0_0 : NAND2
      port map(A => \NLBCLR_c\, B => RUN_c_0_0, Y => CLEAR_0_i_0);
    
    \SOFT_PON_GENERATE_cnt2[11]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_19, Q => \cnt2[11]\);
    
    cnt2_2 : MUX2H
      port map(A => \cnt2_0[1]\, B => N_254, S => \un4_ticki\, Y
         => \cnt2_2\);
    
    un3_activity_I_87 : AND3
      port map(A => \REG[469]\, B => \REG[470]\, C => \REG[471]\, 
        Y => \DWACT_FINC_E_0[9]\);
    
    \SOFT_PON_GENERATE_P_SoftPON_cnt1[2]\ : DFF
      port map(CLK => CLK_c_c, D => cnt1_5, Q => \cnt1[2]\);
    
    un3_activity_I_69 : AND3
      port map(A => \REG[466]\, B => \REG[467]\, C => \REG[468]\, 
        Y => \DWACT_FINC_E[7]\);
    
    TCNT3_2_I_30 : XOR2
      port map(A => \TCNT3[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, Y => \TCNT3_2[3]\);
    
    SOFT_PON_GENERATE_cnt2_19 : MUX2H
      port map(A => \cnt2_2[11]\, B => \cnt2[11]\, S => stop2, Y
         => cnt2_19);
    
    \TCNT2[4]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT2_2[4]\, Q => 
        \TCNT2_i_i[4]\);
    
    HWRES_36 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_36);
    
    \SOFT_PON_GENERATE_cnt2[14]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_22, Q => \cnt2[14]\);
    
    \TCNT3[6]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT3_2[6]\, Q => 
        \TCNT3_i_i[6]\);
    
    \SOFT_PON_GENERATE_cnt2[3]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_11, Q => \cnt2[3]\);
    
    cnt2_2_0_I_118 : AND3
      port map(A => \DWACT_FINC_E_0[7]\, B => \DWACT_FINC_E[9]\, 
        C => \DWACT_FINC_E[12]\, Y => \DWACT_FINC_E[13]\);
    
    \SOFT_PON_GENERATE_cnt2[19]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_27, Q => \cnt2[19]\);
    
    un6_tcnt1_i_0_2 : OR3
      port map(A => \TCNT1_i_i[1]\, B => \TCNT1_i_i[4]\, C => 
        \TCNT1[5]_net_1\, Y => un6_tcnt1_i_0_2_i);
    
    \ACTIVITY[4]\ : DFFC
      port map(CLK => ALICLK_c, D => I_20, CLR => \CLEAR_1\, Q
         => \REG[461]\);
    
    cnt2_2_0_I_224 : XOR2
      port map(A => N_4_1, B => \cnt2[31]\, Y => \cnt2_2_i_i[31]\);
    
    HWRES_29 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_29);
    
    cnt2_2_0_I_195 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[30]\, 
        C => \DWACT_FINC_E[23]\, Y => N_24);
    
    cnt2_2_0_I_94 : AND2
      port map(A => \DWACT_FINC_E_0[7]\, B => \DWACT_FINC_E[9]\, 
        Y => \DWACT_FINC_E[10]\);
    
    LongSoftPON_1 : DFF
      port map(CLK => CLK_c_c, D => LongSoftPON_1_i, Q => 
        \TST_c_1[15]\);
    
    cnt2_2_0_I_30 : AND3
      port map(A => \DWACT_FINC_E_0[0]\, B => \DWACT_FINC_E[1]\, 
        C => \cnt2[5]\, Y => N_141);
    
    TCNT2_2_I_28 : XOR2
      port map(A => \TCNT2_i_i[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => \TCNT2_2[4]\);
    
    EV_RESi : DFFC
      port map(CLK => ALICLK_c, D => \EV_RESi_1\, CLR => 
        un8_hwresi_i, Q => EV_RES_c);
    
    cnt2_2_0_I_19 : AND2
      port map(A => \cnt2[3]\, B => \DWACT_FINC_E_0[0]\, Y => 
        N_149);
    
    \CLEAR_18\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_18);
    
    HWRES_12 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_12);
    
    SOFT_PON_GENERATE_cnt2_15 : MUX2H
      port map(A => \cnt2_2[7]\, B => \cnt2[7]\, S => stop2, Y
         => cnt2_15);
    
    \CLEAR_28\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_28);
    
    un10_tcnt2_i_o3_2 : OR2
      port map(A => \TCNT2_i_i[2]\, B => \TCNT2[3]_net_1\, Y => 
        un10_tcnt2_i_o3_2_i);
    
    cnt2_2_0_I_132 : AND3
      port map(A => \cnt2[18]\, B => \cnt2[19]\, C => \cnt2[20]\, 
        Y => \DWACT_FINC_E[15]\);
    
    \SOFT_PON_GENERATE_cnt2[25]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_33, Q => \cnt2[25]\);
    
    BNC_RESi_0 : DFFC
      port map(CLK => ALICLK_c, D => \BNC_RESi_1\, CLR => 
        un8_hwresi_i, Q => LBSP_c_0(2));
    
    SOFT_PON_GENERATE_cnt2_29 : MUX2H
      port map(A => \cnt2_2_i_i[21]\, B => \cnt2[21]\, S => 
        stop2_1, Y => cnt2_29);
    
    SOFT_PON_GENERATE_cnt2_10 : MUX2H
      port map(A => \cnt2_2[2]\, B => \cnt2[2]\, S => stop2, Y
         => cnt2_10);
    
    HWRES_25 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_25);
    
    cnt2_2_0_I_69 : AND3
      port map(A => \cnt2[9]\, B => \cnt2[10]\, C => \cnt2[11]\, 
        Y => \DWACT_FINC_E_0[7]\);
    
    cnt2_2_0_I_121 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \cnt2[18]\, Y => N_76);
    
    TCNT4_2_I_18 : XOR2
      port map(A => \TCNT4_i_0_i[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, Y => \TCNT4_2[2]\);
    
    TCNT3_2_I_32 : XOR2
      port map(A => \TCNT3_i_i[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, Y => \TCNT3_2[2]\);
    
    HWRES_8 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_8);
    
    HWRES_32_0 : NAND3
      port map(A => N_259_1, B => NPWON_c_1, C => \TST_c_1[15]\, 
        Y => HWRES_c_32_0);
    
    un3_activity_I_90 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[7]\, C
         => \DWACT_FINC_E_0[9]\, Y => N_4_2);
    
    cnt2_2_0_I_37 : AND3
      port map(A => \DWACT_FINC_E_0[0]\, B => \DWACT_FINC_E[2]\, 
        C => \cnt2[6]\, Y => N_136);
    
    HWRES_11 : NAND3
      port map(A => N_259_3, B => NPWON_c_3, C => \TST_c_3[15]\, 
        Y => HWRES_c_11);
    
    cnt2_1 : XOR2
      port map(A => \cnt2_0[0]\, B => \un4_ticki\, Y => \cnt2_1\);
    
    un3_activity_I_80 : AND2
      port map(A => \REG[469]\, B => \REG[470]\, Y => 
        \DWACT_FINC_E_0[8]\);
    
    SOFT_PON_GENERATE_P_SoftPON_un3_stop2_i : NAND3
      port map(A => un3_stop2_i_0, B => I_9_1, C => I_13_2, Y => 
        un3_stop2_i);
    
    TCNT2_2_I_1 : AND2
      port map(A => \TCNT2_i_i[0]\, B => \TICK[0]\, Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    HWRES_0_4 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => HWRES_c_0_4);
    
    \CLEAR_15\ : OR3FTT
      port map(A => LOAD_RES_1, B => HWRES_c_0_1, C => 
        CLEAR_0_i_1, Y => CLEAR_15);
    
    \SOFT_PON_GENERATE_cnt2[8]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_16, Q => \cnt2[8]\);
    
    \CLEAR_25\ : OR3FTT
      port map(A => LOAD_RES_0, B => \HWRES_c_0_0\, C => 
        CLEAR_0_i_0, Y => CLEAR_25);
    
    \TICKi[0]\ : DFF
      port map(CLK => CLK_c_c, D => N_269_i_0, Q => \TICK[0]\);
    
    un11_tcnt3_i_0_1 : OR2
      port map(A => \TCNT3_i_i[4]\, B => \TCNT3[5]_net_1\, Y => 
        un11_tcnt3_i_0_1_i);
    
    stop : DFFC
      port map(CLK => CLK_c_c, D => \stop_7\, CLR => \HWRES_c_3\, 
        Q => \stop\);
    
    TCNT3_2_I_34 : XOR2
      port map(A => \TCNT3[7]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_2_0[0]\, Y => \TCNT3_2[7]\);
    
    TCNT4_2_I_21 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_1[0]\, B => 
        \TCNT4_i_0_i[2]\, Y => \DWACT_ADD_CI_0_g_array_12_3[0]\);
    
    SOFT_PON_GENERATE_cnt2_25 : MUX2H
      port map(A => \cnt2_2[17]\, B => \cnt2[17]\, S => stop2_1, 
        Y => cnt2_25);
    
    un3_activity_I_73 : XOR2
      port map(A => N_17, B => \REG[469]\, Y => I_73);
    
    un12_tcnt3_i : NOR2
      port map(A => \un11_tcnt3_i_0\, B => \un10_tcnt2_i_o3\, Y
         => \un12_tcnt3_i\);
    
    \SOFT_PON_GENERATE_cnt2[13]\ : DFF
      port map(CLK => CLK_c_c, D => cnt2_21, Q => \cnt2[13]\);
    
    SOFT_PON_GENERATE_P_SoftPON_stop2 : DFF
      port map(CLK => CLK_c_c, D => stop2_40_i_a3, Q => stop2);
    
    cnt2_2_0_I_172 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[19]\, Y => N_40);
    
    TCNT2_2_I_45 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11[0]\, B => 
        \TCNT2_i_i[6]\, Y => \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    \TCNT2[7]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT2_2[7]\, Q => 
        \TCNT2[7]_net_1\);
    
    HWRES_0_2 : NAND3
      port map(A => N_259_0, B => NPWON_c_0, C => \TST_c_0[15]\, 
        Y => \HWRES_c_0_2\);
    
    un2_hwresi : OR2
      port map(A => REG_0, B => SYSRESB_c, Y => N_259);
    
    SOFT_PON_GENERATE_P_SoftPON_cnt1_5 : MUX2H
      port map(A => I_9_1, B => \cnt1[2]\, S => \un1_stop2_1_0\, 
        Y => cnt1_5);
    
    SoftPON1 : DFF
      port map(CLK => CLK_c_c, D => \TST_c[14]\, Q => \TST_c[13]\);
    
    cnt2_2_0_I_8 : AND2
      port map(A => \cnt2[1]_net_1\, B => \cnt2[0]_net_1\, Y => 
        N_157);
    
    \TCNT3[5]\ : DFF
      port map(CLK => CLK_c_c, D => \TCNT3_2[5]\, Q => 
        \TCNT3[5]_net_1\);
    
    HWRES_24 : NAND3
      port map(A => N_259_2, B => NPWON_c_2, C => \TST_c_2[15]\, 
        Y => HWRES_c_24);
    
    SOFT_PON_GENERATE_P_SoftPON_un3_stop2_i_0 : AND2FT
      port map(A => \cnt1[0]\, B => I_5_1, Y => un3_stop2_i_0);
    
    SOFT_PON_GENERATE_cnt2_20 : MUX2H
      port map(A => \cnt2_2[12]\, B => \cnt2[12]\, S => stop2_1, 
        Y => cnt2_20);
    
    cnt2_2_0_I_139 : AND2
      port map(A => \DWACT_FINC_E[15]\, B => \cnt2[21]\, Y => 
        \DWACT_FINC_E[16]\);
    
    cnt2_2_0_I_111 : AND3
      port map(A => \DWACT_FINC_E_0[0]\, B => \DWACT_FINC_E[2]\, 
        C => \DWACT_FINC_E[5]\, Y => \DWACT_FINC_E[28]\);
    
    cnt2_2_0_I_73 : XOR2
      port map(A => N_111, B => \cnt2[12]\, Y => \cnt2_2[12]\);
    
    cnt2_2_0_I_217 : XOR2
      port map(A => N_9, B => \cnt2[30]\, Y => \cnt2_2[30]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity SPI_INTERF is

    port( CROMWDT        : out   std_logic_vector(7 downto 0);
          DACCFG_WDT     : out   std_logic_vector(13 downto 4);
          TICK           : in    std_logic_vector(1 to 1);
          FBOUT          : out   std_logic_vector(7 downto 0);
          REG_i_0        : in    std_logic_vector(80 to 80);
          REG_400        : out   std_logic;
          REG_398        : out   std_logic;
          REG_396        : out   std_logic;
          REG_393        : out   std_logic;
          REG_0          : in    std_logic;
          REG_1          : in    std_logic;
          REG_2          : in    std_logic;
          REG_3          : in    std_logic;
          REG_4          : in    std_logic;
          REG_5          : in    std_logic;
          REG_6          : in    std_logic;
          REG_7          : in    std_logic;
          REG_8          : in    std_logic;
          REG_399        : out   std_logic;
          REG_395        : out   std_logic;
          REG_397        : out   std_logic;
          REG_394        : out   std_logic;
          CROMWAD        : out   std_logic_vector(8 downto 0);
          sstate_0_2     : out   std_logic;
          PULSE_6        : in    std_logic;
          PULSE_0        : in    std_logic;
          PULSE_10       : in    std_logic;
          sstate_0_i_0   : in    std_logic_vector(2 to 2);
          HWRES_c_30     : in    std_logic;
          HWRES_c_23_0   : in    std_logic;
          HWRES_c_28     : in    std_logic;
          HWRES_c_31     : in    std_logic;
          HWRES_c_24     : in    std_logic;
          HWRES_c_25     : in    std_logic;
          DACCFG_nWR     : out   std_logic;
          PDLCFG_nWR     : out   std_logic;
          HWRES_c_32     : in    std_logic;
          WRCROM         : out   std_logic;
          HWRES_c_26     : in    std_logic;
          HWRES_c_27     : in    std_logic;
          NCYC_RELOAD_in : in    std_logic;
          HWRES_c_29     : in    std_logic;
          un1_drive_spi  : out   std_logic;
          F_SO_c         : in    std_logic;
          LOAD_RES       : out   std_logic;
          DRIVE_RELOAD   : out   std_logic;
          ISCK           : out   std_logic;
          FWIMG2LOAD     : in    std_logic;
          ISI            : out   std_logic;
          FCS_c          : out   std_logic;
          PON_LOAD_i     : in    std_logic;
          HWRES_c_32_0   : in    std_logic;
          LOAD_RES_0     : out   std_logic;
          LOAD_RES_1     : out   std_logic;
          LOAD_RES_2     : out   std_logic;
          CLK_c_c        : in    std_logic;
          HWRES_c_27_0   : in    std_logic;
          LOAD_RES_3     : out   std_logic
        );

end SPI_INTERF;

architecture DEF_ARCH of SPI_INTERF is 

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component AOI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_1038, \sstate_0[0]_net_1\, \sstate_0[3]_net_1\, 
        N_1054, N_412, N_1047, G_0_0_i, G_0_1_i, \G\, N_425, 
        \RESCNT_6[15]\, N_313_0, \G_5\, N_528_i_0_0, 
        \RESCNT[15]_net_1\, \G_4\, G_4_4_i, G_4_3_i, 
        \DWACT_ADD_CI_0_pog_array_2_1[0]\, \RESCNT[0]_net_1\, 
        \RESCNT[1]_net_1\, G_4_0_i, 
        \DWACT_ADD_CI_0_pog_array_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_5[0]\, \RESCNT[14]_net_1\, 
        \DWACT_ADD_CI_0_TMP[0]\, \DWACT_ADD_CI_0_g_array_11_2[0]\, 
        G_2_3_i, G_2_2_i, G_2_0, \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_g_array_10[0]\, G_2_i, G_1_i, 
        \DWACT_ADD_CI_0_g_array_2[0]\, \G_0_0\, 
        \DWACT_ADD_CI_0_g_array_3[0]\, G_1_1, \LOAD_RESi_1\, 
        \sstate_ns[0]\, \sstate_0[1]_net_1\, \sstate_ns[1]\, 
        N_846_i_0, N_1022_i_0, \sstate_0[4]_net_1\, 
        \sstate_ns[4]\, N_1078_2, N_1078_1, N_1078_0, N_313_7_i, 
        N_402_0, N_401, N_1041, \DWACT_ADD_CI_0_g_array_2_0[0]\, 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_3_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_2_0[0]\, 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_g_array_3_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_2_2[0]\, 
        \DWACT_ADD_CI_0_g_array_11_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_3[0]\, 
        \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_11_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1_1[0]\, 
        \DWACT_ADD_CI_0_TMP_0[0]\, \PAGECNT_i_0_i[1]\, 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, \PAGECNT[4]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12[0]\, \PAGECNT[2]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, \PAGECNT[6]_net_1\, 
        \DWACT_ADD_CI_0_g_array_11_3[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1_2[0]\, 
        \DWACT_ADD_CI_0_TMP_1[0]\, 
        \DWACT_ADD_CI_0_g_array_12_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, 
        \DWACT_ADD_CI_0_g_array_12_2_0[0]\, 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, 
        \DWACT_ADD_CI_0_TMP_2[0]\, \BITCNT[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, \RESCNT[2]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_2_1[0]\, \RESCNT[6]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_4[0]\, \RESCNT[10]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_5[0]\, \RESCNT[12]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_3_0[0]\, \RESCNT[8]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_1_1[0]\, \RESCNT[4]_net_1\, 
        \DWACT_ADD_CI_0_g_array_1_3[0]\, 
        \DWACT_ADD_CI_0_TMP_3[0]\, 
        \DWACT_ADD_CI_0_g_array_2_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\, 
        \DWACT_ADD_CI_0_g_array_11_4[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1_3[0]\, 
        \DWACT_ADD_CI_0_g_array_12_1_2[0]\, 
        \DWACT_ADD_CI_0_g_array_12_6[0]\, 
        \DWACT_ADD_CI_0_g_array_12_2_2[0]\, \RELOAD_EDGE_i\, 
        \RELOAD_EDGE\, N_363_1, \sstate_ns_1_iv_i_5[3]_net_1\, 
        N_295_i, \sstate_ns_1_iv_i_3_i[3]\, 
        \sstate_ns_1_iv_i_2_i[3]\, N_392, N_289, N_407, N_219, 
        N_394, N_1053, N_343_1, \sstate_ns_1_iv_i_1[3]_net_1\, 
        N_293, N_292_i, \sstate_0[2]_net_1\, N_414, 
        \sstate[4]_net_1\, \sstate_ns_1_iv_i_0_4[2]_net_1\, 
        N_1050, \sstate[2]_net_1\, N_7181_i, 
        \sstate_ns_1_iv_i_0_2_i[2]\, \sstate_ns_1_iv_i_0_1_i[2]\, 
        N_1039, \sstate_ns_1_iv_i_0_0[2]_net_1\, N_416, N_396_1, 
        N_426, \sstate[1]_net_1\, N_362, \sstate[3]_net_1\, N_423, 
        N_413, \NCS0\, \FCS_SEL\, \un1_sstate_26_0_0_i\, N_282, 
        N_283, N_354_1, N_237, \sstate[0]_net_1\, N_1058, N_361, 
        \sstate_ns_0_0_0_0[4]_net_1\, N_348, N_422, N_420, N_433, 
        N_1078, \LUT_5_i_0\, \LUT\, N_216, N_436_1, 
        \COMMAND_3_i_0\, \COMMAND\, N_7179_i, N_353_i, 
        \sstate_ns_1_iv_0_0_3_i[1]\, \sstate_ns_1_iv_0_0_1_i[1]\, 
        \sstate_ns_1_iv_0_0_0_i[1]\, N_7176_i, N_421, N_417, 
        \sstate_ns_1_iv_0_0_a3_4[1]_net_1\, N_418, N_1074, 
        \sstate_ns_1_iv_0_0_a3_2[1]_net_1\, 
        \sstate_ns_1_iv_0_0_a3_2_0[1]_net_1\, 
        \sstate_ns_1_iv_0_0_a3_0_i[1]\, \sstate_i_0[0]\, N_353_1, 
        N_406, N_382_i, N_1076, N_1047_i_0, N_1078_i_0, 
        \sstate_ns_1_iv_0_0_3_i[0]\, N_373_i, 
        \sstate_ns_1_iv_0_0_2_i[0]\, 
        \sstate_ns_1_iv_0_0_a3_3_0[0]_net_1\, 
        \sstate_ns_1_iv_0_0_1[0]_net_1\, N_424, N_1063, 
        \sstate_ns_1_iv_0_0_0[0]_net_1\, 
        \sstate_ns_1_iv_0_0_a3_4_1[0]_net_1\, 
        \sstate_ns_1_iv_0_0_0_tz_0[0]_net_1\, N_427_1, N_390, 
        \sstate_i_0[3]\, N_434, 
        \sstate_ns_1_iv_0_0_a3_1[0]_net_1\, \DACCfgValue_29\, 
        \DACCfgValue[13]_net_1\, N_1011, N_945, N_991, 
        \DACCfgValue_28\, \DACCfgValue[12]_net_1\, N_1012, 
        \DACCfgValue_27\, \DACCfgValue[11]_net_1\, 
        \DACCfgValue_9[11]\, N_276, N_275, N_402, 
        \DACCfgValue_26\, \DACCfgValue[10]_net_1\, 
        \DACCfgValue_9[10]\, N_274, N_273, \DACCfgValue_25\, 
        \DACCfgValue[9]_net_1\, \DACCfgValue_9[9]\, N_272, N_271, 
        \DACCfgValue_24\, \DACCfgValue[8]_net_1\, 
        \DACCfgValue_9[8]\, N_270, N_269, \DACCfgValue_23\, 
        \DACCfgValue[7]_net_1\, \DACCfgValue_9[7]\, N_268, N_267, 
        \DACCfgValue_22\, \DACCfgValue[6]_net_1\, 
        \DACCfgValue_9[6]\, N_266, N_265, \DACCfgValue_21\, 
        \DACCfgValue[5]_net_1\, \DACCfgValue_9[5]\, N_264, N_263, 
        \FBOUT[1]\, \DACCfgValue_20\, \DACCfgValue[4]_net_1\, 
        \DACCfgValue_9[4]\, N_317, N_261, N_260, \FBOUT[0]\, 
        \WRDACi_19\, \WRDACi\, N_946, un1_pulse_1, N_383_i, 
        N_384_i, N_395, \CROMWAD[6]\, N_1064, N_1042, \WRPDLi_18\, 
        \WRPDLi\, N_944, \WRPDLi_0_sqmuxa_1_i_0_a3_1\, N_435, 
        \CROMWAD_i_0[7]\, \CROMWAD[4]\, \WRCROMi_17\, \WRCROMi\, 
        N_943, N_315, N_1043, \WRCROMi_0_sqmuxa_1_i_0_a3_0\, 
        \CROMWAD[7]\, \CROMWAD[8]\, N_391, N_389, \ISI_16\, ISI_8, 
        un1_ISI_1_sqmuxa_1, un1_ISI_1_sqmuxa_1_0_1_0_i, N_350_i, 
        N_351, N_115_i, N_559, \un1_pulse_7_0_0_0_0\, N_248, 
        N_235, \FBOUT[7]\, \NCS0_15\, NCS0_6, un1_NCS0_2_sqmuxa, 
        N_344, \un1_NCS0_2_sqmuxa_0_0_0_0\, N_410, N_1033_i, 
        N_359, \SBYTE_14\, \SBYTE_7[7]\, un1_SBYTE_0_sqmuxa, 
        N_334, N_332, N_1075, \FBOUT[6]\, N_1046, \SBYTE_13\, 
        \SBYTE_7[6]\, N_331, N_330, \FBOUT[5]\, \SBYTE_12\, 
        \SBYTE_7[5]\, N_329, N_328, \FBOUT[4]\, \SBYTE_11\, 
        \SBYTE_7[4]\, N_325_i, N_324_i, \FBOUT[3]\, \SBYTE_10\, 
        \SBYTE_7[3]\, N_327, N_326, \FBOUT[2]\, \SBYTE_9\, 
        \SBYTE_7[2]\, N_323_i, N_322_i, \SBYTE_8\, \SBYTE_7[1]\, 
        N_321_i, N_320_i, \SBYTE_7\, \SBYTE_7[0]\, N_218_i_i, 
        N_432, N_319_i, N_318_i, \F_SO_maj\, N_1044, \FCS_SEL_6\, 
        un1_pulse_3, un1_FCS_SEL_0_sqmuxa, N_281_i, N_280_i, 
        N_405, N_1038_i_0, N_1050_i_0, \ISCK_4\, sstate_26_sqmuxa, 
        N_498, N_349_i, un1_ISCK_1_sqmuxa_i_0_0_2_i, 
        un1_ISCK_1_sqmuxa_i_0_0_1_i, N_347_i, 
        \un1_ISCK_1_sqmuxa_i_0_0_a3\, 
        un1_ISCK_1_sqmuxa_i_0_0_a3_1_0_i, N_247_i, \N_414_i\, 
        \DRIVE_RELOAD_2\, RESCNT_1_sqmuxa, un1_LOAD_RESi_0_sqmuxa, 
        \BYTECNT_9[8]\, N_437_i_0, I_36, \BYTECNT_9[7]\, I_34, 
        \BYTECNT_9[6]\, I_38_1, \BYTECNT_9[5]\, I_33, 
        \BYTECNT_9[4]\, I_30_0, \BYTECNT_9[3]\, N_312, I_37, 
        un1_pulse_9, \BYTECNT_9[2]\, I_35, \BYTECNT_9[1]\, I_32, 
        \BYTECNT_9[0]\, \DWACT_ADD_CI_0_partial_sum[0]\, N_351_1, 
        \un1_pulse_9_0_0_0\, N_399, \un1_pulse_9_0_0_a2_0_0\, 
        N_409, N_1059, N_408, N_398, \PAGECNT_9[8]\, N_436_i_0, 
        I_36_0, \PAGECNT_9[7]\, I_34_0, \PAGECNT_9[6]\, I_38_2, 
        \PAGECNT_9[5]\, I_33_0, \PAGECNT_9[4]\, I_30_1, 
        \PAGECNT_9[3]\, I_37_0, \PAGECNT_9[2]\, I_35_0, 
        \PAGECNT_9[1]\, I_32_0, \PAGECNT_9[0]\, 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, 
        un1_ISCK_1_sqmuxa_i_0_0_o2_0_i, 
        un1_ISCK_1_sqmuxa_i_0_0_o2_1_i, N_143_i_0, 
        \PAGECNT_i_0_i[3]\, N_1065, N_1045, N_1062, N_419, N_411, 
        LUT_5_i_0_a2_0_0_i, LUT_5_i_0_a2_0_1_i, 
        \sstate_ns_1_iv_0_a2_9_0_a2_i_2_i[0]\, \PAGECNT_i_i[7]\, 
        \PAGECNT[8]_net_1\, \PAGECNT_i_i[0]\, \PAGECNT_i_i[5]\, 
        \RESCNT_6[14]\, I_65, \RESCNT_6[13]\, I_60, 
        \RESCNT_6[12]\, I_58, \RESCNT_6[11]\, I_56_1, 
        \RESCNT_6[10]\, I_53, \RESCNT_6[9]\, I_52_1, 
        \RESCNT_6[8]\, I_63, \RESCNT_6[7]\, N_313, I_61, 
        N_528_i_0, \RESCNT_6[6]\, I_59, \RESCNT_6[5]\, I_57, 
        \RESCNT_6[4]\, I_55, \RESCNT_6[3]\, I_54, \RESCNT_6[2]\, 
        I_51, \RESCNT_6[1]\, I_64, \RESCNT_6[0]\, 
        \DWACT_ADD_CI_0_partial_sum_1[0]\, 
        \RESCNT_6_0_a3_7_12_i[0]\, \RESCNT_6_0_a3_7_8_i[0]\, 
        \RESCNT_6_0_a3_7_9_i[0]\, \RESCNT_6_0_a3_7_4[0]_net_1\, 
        \RESCNT[5]_net_1\, \RESCNT[7]_net_1\, 
        \RESCNT_6_0_a3_7_6[0]_net_1\, \RESCNT[3]_net_1\, 
        \RESCNT_6_0_a3_7_10_i[0]\, \RESCNT_6_0_a3_7_0_i[0]\, 
        \RESCNT_6_0_a3_7_1_i[0]\, \RESCNT[13]_net_1\, 
        \RESCNT_6_0_a3_7_2[0]_net_1\, \RESCNT[9]_net_1\, 
        \RESCNT[11]_net_1\, \BITCNT_8[2]\, I_14_0, N_562, 
        \BITCNT_8[1]\, I_13_4, \BITCNT_8[0]\, 
        \DWACT_ADD_CI_0_partial_sum_2[0]\, \ISI_8_iv_0_i_o2_0\, 
        \BITCNT[0]_net_1\, \BITCNT[2]_net_1\, N_415_i, N_7115_i, 
        F_SO_maj_2, N_342, N_700, \F_SO_sync1\, \F_SO_sync2\, 
        \F_SO_sync\, \un1_sstate_25_0_0_0\, 
        un1_sstate_25_0_0_0_1_i, un1_sstate_25_0_0_0_0_i, 
        \sstate_ns_1_iv_i_o2_0[3]_net_1\, \CROMWAD[3]\, 
        \CROMWAD[2]\, \CROMWAD[1]\, N_1040, 
        \un1_sstate_1_sqmuxa_0_0_0\, N_278, \CROMWAD[5]\, 
        F_SO_sync2_2, F_SO_sync1_2, F_SO_sync_2, un3_reload_edge, 
        RELOAD_EDGE_r_i_0, \LOAD_RES\, ISI_net_1, ISCK_net_1, 
        DRIVE_RELOAD_net_1, \CROMWAD[0]\, 
        \DWACT_ADD_CI_0_partial_sum_3[0]\, \REG[474]\, 
        \RELOAD_CNT_3[1]\, \REG[475]\, \RELOAD_CNT_3[2]\, 
        \RELOAD_CNT_3[3]\, \REG[477]\, \RELOAD_CNT_3[4]\, 
        \RELOAD_CNT_3[5]\, \REG[479]\, \RELOAD_CNT_3[6]\, 
        \RELOAD_CNT_3[7]\, \REG[478]\, \REG[476]\, \REG[480]\, 
        \REG[473]\, \DWACT_ADD_CI_0_pog_array_1_4[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_2_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_2_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_2_2[0]\, \GND\, \VCC\
         : std_logic;

begin 

    FBOUT(7) <= \FBOUT[7]\;
    FBOUT(6) <= \FBOUT[6]\;
    FBOUT(5) <= \FBOUT[5]\;
    FBOUT(4) <= \FBOUT[4]\;
    FBOUT(3) <= \FBOUT[3]\;
    FBOUT(2) <= \FBOUT[2]\;
    FBOUT(1) <= \FBOUT[1]\;
    FBOUT(0) <= \FBOUT[0]\;
    REG_400 <= \REG[480]\;
    REG_398 <= \REG[478]\;
    REG_396 <= \REG[476]\;
    REG_393 <= \REG[473]\;
    REG_399 <= \REG[479]\;
    REG_395 <= \REG[475]\;
    REG_397 <= \REG[477]\;
    REG_394 <= \REG[474]\;
    CROMWAD(8) <= \CROMWAD[8]\;
    CROMWAD(7) <= \CROMWAD[7]\;
    CROMWAD(6) <= \CROMWAD[6]\;
    CROMWAD(5) <= \CROMWAD[5]\;
    CROMWAD(4) <= \CROMWAD[4]\;
    CROMWAD(3) <= \CROMWAD[3]\;
    CROMWAD(2) <= \CROMWAD[2]\;
    CROMWAD(1) <= \CROMWAD[1]\;
    CROMWAD(0) <= \CROMWAD[0]\;
    sstate_0_2 <= \sstate_0[2]_net_1\;
    LOAD_RES <= \LOAD_RES\;
    DRIVE_RELOAD <= DRIVE_RELOAD_net_1;
    ISCK <= ISCK_net_1;
    ISI <= ISI_net_1;

    \sstate_ns_1_iv_0_0_a2_0[0]\ : AND2
      port map(A => \sstate_0[1]_net_1\, B => \sstate_0[2]_net_1\, 
        Y => N_424);
    
    \SBYTE[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_11\, CLR => HWRES_c_31, 
        Q => \FBOUT[4]\);
    
    \SBYTE_7_1_i_a3[6]\ : NOR2
      port map(A => N_1046, B => REG_7, Y => N_330);
    
    \BITCNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_8[0]\, CLR => 
        HWRES_c_23_0, Q => \BITCNT[0]_net_1\);
    
    un1_RESCNT_I_61 : XOR2
      port map(A => \RESCNT[7]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_2_1[0]\, Y => I_61);
    
    un1_FCS_SEL_0_sqmuxa_0_0_0_a3 : NOR2FT
      port map(A => PULSE_6, B => N_405, Y => N_280_i);
    
    \RESCNT[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[12]\, CLR => 
        HWRES_c_30, Q => \RESCNT[12]_net_1\);
    
    un1_RESCNT_G : AND3FFT
      port map(A => G_2_i, B => G_1_i, C => \G\, Y => 
        \DWACT_ADD_CI_0_g_array_10[0]\);
    
    \RELOAD_CNT[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \RELOAD_CNT_3[7]\, CLR => 
        HWRES_c_29, Q => \REG[480]\);
    
    LOAD_RESi_2 : DFFS
      port map(CLK => CLK_c_c, D => \LOAD_RESi_1\, SET => 
        HWRES_c_27_0, Q => LOAD_RES_2);
    
    \SBYTE_7_1_i_a3[3]\ : NOR2
      port map(A => N_1046, B => REG_4, Y => N_326);
    
    \sstate_ns_1_iv_0_0_a2[1]\ : NOR3FFT
      port map(A => N_1047_i_0, B => N_1078_i_0, C => N_414, Y
         => N_382_i);
    
    \sstate_ns_1_iv_0_0_3[1]\ : OR3
      port map(A => \sstate_ns_1_iv_0_0_1_i[1]\, B => 
        \sstate_ns_1_iv_0_0_0_i[1]\, C => N_7176_i, Y => 
        \sstate_ns_1_iv_0_0_3_i[1]\);
    
    WRPDLi_0_sqmuxa_1_i_0_o2 : NAND2
      port map(A => \CROMWAD[4]\, B => \CROMWAD[5]\, Y => N_1064);
    
    LUT_5_i_0_a2 : NAND2
      port map(A => N_389, B => N_411, Y => N_414);
    
    \DACCfgValue_9_i_a3_0[4]\ : NOR2
      port map(A => \FBOUT[0]\, B => N_402, Y => N_261);
    
    un1_RESCNT_I_54 : XOR2
      port map(A => \RESCNT[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, Y => I_54);
    
    \sstate_0[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns[4]\, CLR => 
        HWRES_c_32_0, Q => \sstate_0[4]_net_1\);
    
    \PAGECNT_9_0_a3[1]\ : AND2
      port map(A => N_436_i_0, B => I_32_0, Y => \PAGECNT_9[1]\);
    
    ISI_8_r : NOR3
      port map(A => N_115_i, B => N_559, C => 
        \un1_pulse_7_0_0_0_0\, Y => ISI_8);
    
    un1_PAGECNT_1_I_53 : AND2
      port map(A => \PAGECNT[4]_net_1\, B => \PAGECNT_i_i[5]\, Y
         => \DWACT_ADD_CI_0_pog_array_1_1_1[0]\);
    
    ISI_8_iv_0_i_o2_0_0 : AND2
      port map(A => \BITCNT[1]_net_1\, B => \BITCNT[2]_net_1\, Y
         => \ISI_8_iv_0_i_o2_0\);
    
    un1_PAGECNT_1_I_52 : AND2
      port map(A => \PAGECNT[2]_net_1\, B => \PAGECNT_i_0_i[3]\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_0[0]\);
    
    \sstate_ns_1_iv_i_o2_5[3]\ : OR2FT
      port map(A => \CROMWAD[0]\, B => \CROMWAD[7]\, Y => N_1040);
    
    \ISCK\ : DFFC
      port map(CLK => CLK_c_c, D => \ISCK_4\, CLR => HWRES_c_27, 
        Q => ISCK_net_1);
    
    \sstate_ns_1_iv_i_0_1[2]\ : OAI21
      port map(A => N_1039, B => \sstate_0[0]_net_1\, C => 
        \sstate_ns_1_iv_i_0_0[2]_net_1\, Y => 
        \sstate_ns_1_iv_i_0_1_i[2]\);
    
    SBYTE_9 : MUX2H
      port map(A => \FBOUT[2]\, B => \SBYTE_7[2]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_9\);
    
    \DACCfgValue[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_26\, CLR => 
        HWRES_c_25, Q => \DACCfgValue[10]_net_1\);
    
    \sstate_0[2]\ : DFFS
      port map(CLK => CLK_c_c, D => N_846_i_0, SET => 
        HWRES_c_32_0, Q => \sstate_0[2]_net_1\);
    
    LOAD_RESi_3 : DFFS
      port map(CLK => CLK_c_c, D => \LOAD_RESi_1\, SET => 
        HWRES_c_27_0, Q => LOAD_RES_3);
    
    \DACCFG_WDT_1[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[4]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(4));
    
    un1_pulse_6_i_0_i_a3 : OR2FT
      port map(A => N_1058, B => N_410, Y => N_359);
    
    F_SO_sync2 : DFFC
      port map(CLK => CLK_c_c, D => F_SO_sync2_2, CLR => 
        HWRES_c_27, Q => \F_SO_sync2\);
    
    F_SO_sync1 : DFFC
      port map(CLK => CLK_c_c, D => F_SO_sync1_2, CLR => 
        HWRES_c_27, Q => \F_SO_sync1\);
    
    \PDLCFG_WDT_1[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[7]\, CLR => HWRES_c_29, 
        Q => CROMWDT(7));
    
    un1_sstate_26_0_0_i_o2_0 : NOR2
      port map(A => N_1058, B => \sstate[2]_net_1\, Y => N_237);
    
    un1_FCS_SEL_0_sqmuxa_0_0_a2_1 : OR2FT
      port map(A => \sstate[1]_net_1\, B => \sstate_0[2]_net_1\, 
        Y => N_406);
    
    \SBYTE[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_9\, CLR => HWRES_c_31, 
        Q => \FBOUT[2]\);
    
    LUT_5_i_0_a2_0 : AND3FFT
      port map(A => LUT_5_i_0_a2_0_0_i, B => LUT_5_i_0_a2_0_1_i, 
        C => N_143_i_0, Y => N_389);
    
    un1_ISI_1_sqmuxa_1_0_1_a3 : NOR2FT
      port map(A => N_1053, B => N_1054, Y => N_350_i);
    
    \RESCNT_6_r[3]\ : OA21
      port map(A => N_313, B => I_54, C => N_528_i_0, Y => 
        \RESCNT_6[3]\);
    
    un1_PAGECNT_1_I_34 : XOR2
      port map(A => \PAGECNT_i_i[7]\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => I_34_0);
    
    \sstate_ns_1_iv_0_a2_9_0_a2_i_2[0]\ : OR3
      port map(A => \PAGECNT_i_i[0]\, B => \PAGECNT_i_i[5]\, C
         => \PAGECNT[6]_net_1\, Y => 
        \sstate_ns_1_iv_0_a2_9_0_a2_i_2_i[0]\);
    
    un1_sstate_25_0_0_0_1 : OR2
      port map(A => N_1065, B => N_419, Y => 
        un1_sstate_25_0_0_0_1_i);
    
    un1_RESCNT_I_97 : AND2
      port map(A => \RESCNT[12]_net_1\, B => \RESCNT[13]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_5[0]\);
    
    \sstate_ns_1_iv_i_a2_0[3]\ : NOR2FT
      port map(A => \sstate[2]_net_1\, B => \sstate[1]_net_1\, Y
         => N_407);
    
    \RESCNT_6_0_a3_7_0[0]\ : NAND2
      port map(A => \RESCNT[14]_net_1\, B => \RESCNT[15]_net_1\, 
        Y => \RESCNT_6_0_a3_7_0_i[0]\);
    
    \PDLCFG_WDT_1[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[2]\, CLR => HWRES_c_28, 
        Q => CROMWDT(2));
    
    \DACCfgValue_9_i_a3[9]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[9]_net_1\, Y => 
        N_271);
    
    WRPDLi_18 : MUX2H
      port map(A => \WRPDLi\, B => un1_pulse_1, S => N_944, Y => 
        \WRPDLi_18\);
    
    \DACCFG_WDT_1[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[8]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(8));
    
    un1_LOAD_RESi_1_sqmuxa_1_i_o2_0_0_a2 : AND2FT
      port map(A => N_413, B => \sstate[2]_net_1\, Y => N_419);
    
    WRPDLi : DFFS
      port map(CLK => CLK_c_c, D => \WRPDLi_18\, SET => 
        HWRES_c_32, Q => \WRPDLi\);
    
    \sstate_ns_1_iv_i_o2_1[3]\ : NOR2
      port map(A => N_1041, B => N_1043, Y => N_1045);
    
    SBYTE_8 : MUX2H
      port map(A => \FBOUT[1]\, B => \SBYTE_7[1]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_8\);
    
    \CROMWAD_i[7]\ : INV
      port map(A => \CROMWAD[7]\, Y => \CROMWAD_i_0[7]\);
    
    \BYTECNT_9_0_a3[7]\ : AND2
      port map(A => N_437_i_0, B => I_34, Y => \BYTECNT_9[7]\);
    
    \sstate_ns_1_iv_0_0_a3_4[1]\ : OR2
      port map(A => N_418, B => N_1074, Y => 
        \sstate_ns_1_iv_0_0_a3_4[1]_net_1\);
    
    \RELOAD_CNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \RELOAD_CNT_3[1]\, CLR => 
        HWRES_c_29, Q => \REG[474]\);
    
    un1_RESCNT_I_56 : XOR2
      port map(A => \RESCNT[11]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_4[0]\, Y => I_56_1);
    
    \sstate_ns_1_iv_i_0_i[2]\ : INV
      port map(A => N_1078, Y => N_1078_i_0);
    
    \sstate_ns_1_iv_i_0[2]\ : OA21FTT
      port map(A => N_363_1, B => \sstate[4]_net_1\, C => 
        \sstate_ns_1_iv_i_0_4[2]_net_1\, Y => N_846_i_0);
    
    un1_BYTECNT_3_I_43 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\);
    
    un1_BITCNT_I_9 : XOR2
      port map(A => \BITCNT[0]_net_1\, B => \un1_sstate_25_0_0_0\, 
        Y => \DWACT_ADD_CI_0_partial_sum_2[0]\);
    
    \RESCNT_6_r[9]\ : OA21
      port map(A => N_313_0, B => I_52_1, C => N_528_i_0_0, Y => 
        \RESCNT_6[9]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_44 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_3[0]\, B => 
        \REG[475]\, Y => \DWACT_ADD_CI_0_g_array_12_6[0]\);
    
    COMMAND_3_i_0 : AO21
      port map(A => \COMMAND\, B => N_216, C => N_1078, Y => 
        \COMMAND_3_i_0\);
    
    un1_RESCNT_G_6 : AND2
      port map(A => \RESCNT[0]_net_1\, B => \G\, Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    FCS_SEL_6 : MUX2H
      port map(A => \FCS_SEL\, B => un1_pulse_3, S => 
        un1_FCS_SEL_0_sqmuxa, Y => \FCS_SEL_6\);
    
    \DACCfgValue_9_r[7]\ : NOR3
      port map(A => N_1078_2, B => N_268, C => N_267, Y => 
        \DACCfgValue_9[7]\);
    
    un1_BITCNT_I_13 : XOR2
      port map(A => \BITCNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP_2[0]\, Y => I_13_4);
    
    \RELOAD_CNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \RELOAD_CNT_3[3]\, CLR => 
        HWRES_c_29, Q => \REG[476]\);
    
    G_0_0 : NAND2FT
      port map(A => sstate_0_i_0(2), B => PULSE_10, Y => G_0_0_i);
    
    \BYTECNT_9_r[0]\ : OA21FTT
      port map(A => N_312, B => \DWACT_ADD_CI_0_partial_sum[0]\, 
        C => un1_pulse_9, Y => \BYTECNT_9[0]\);
    
    \BYTECNT_9_0_o2[8]\ : AND2
      port map(A => N_312, B => un1_pulse_9, Y => N_437_i_0);
    
    FCS : MUX2H
      port map(A => REG_i_0(80), B => \NCS0\, S => \FCS_SEL\, Y
         => FCS_c);
    
    LUT_5_i_0_a2_0_i : NOR3
      port map(A => \sstate_ns_1_iv_0_a2_9_0_a2_i_2_i[0]\, B => 
        \PAGECNT_i_i[7]\, C => \PAGECNT[8]_net_1\, Y => N_143_i_0);
    
    un1_sstate_33_i_0_a2 : OAI21TTF
      port map(A => N_383_i, B => N_384_i, C => N_395, Y => N_401);
    
    un1_PAGECNT_1_I_43 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\);
    
    \DACCfgValue_9_i_a3[4]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[4]_net_1\, Y => 
        N_260);
    
    un1_PAGECNT_1_I_42 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_0[0]\);
    
    \sstate_ns_1_iv_0_0_a2_2[0]\ : OR2FT
      port map(A => \sstate[3]_net_1\, B => N_1074, Y => N_1076);
    
    SBYTE_13 : MUX2H
      port map(A => \FBOUT[6]\, B => \SBYTE_7[6]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_13\);
    
    \DACCfgValue[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_27\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[11]_net_1\);
    
    un1_BYTECNT_3_I_34 : XOR2
      port map(A => \CROMWAD[7]\, B => 
        \DWACT_ADD_CI_0_g_array_12_2_0[0]\, Y => I_34);
    
    \DACCfgValue_9_r[10]\ : NOR3
      port map(A => N_1078_2, B => N_274, C => N_273, Y => 
        \DACCfgValue_9[10]\);
    
    \DACCfgValue[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_20\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[4]_net_1\);
    
    \SBYTE_7_1_i_a3_0[5]\ : NOR2FT
      port map(A => N_1075, B => \FBOUT[4]\, Y => N_329);
    
    \sstate_ns_1_iv_i_o2_0[3]\ : NAND2
      port map(A => N_394, B => N_1053, Y => N_219);
    
    \DACCFG_WDT_1[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[7]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(7));
    
    SBYTE_11 : MUX2H
      port map(A => \FBOUT[4]\, B => \SBYTE_7[4]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_11\);
    
    N_1050_i : INV
      port map(A => N_1050, Y => N_1050_i_0);
    
    un1_RESCNT_G_2_0 : AND2
      port map(A => \RESCNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_pog_array_1_5[0]\, Y => G_2_0);
    
    un1_PAGECNT_1_I_1 : AND2
      port map(A => \PAGECNT_i_i[0]\, B => 
        \un1_sstate_1_sqmuxa_0_0_0\, Y => 
        \DWACT_ADD_CI_0_TMP_0[0]\);
    
    \RESCNT_6_r[10]\ : OA21
      port map(A => N_313_0, B => I_53, C => N_528_i_0_0, Y => 
        \RESCNT_6[10]\);
    
    \RESCNT_6_0_a3_7_9[0]\ : NAND3
      port map(A => \RESCNT_6_0_a3_7_4[0]_net_1\, B => 
        \RESCNT[4]_net_1\, C => \RESCNT[5]_net_1\, Y => 
        \RESCNT_6_0_a3_7_9_i[0]\);
    
    \sstate_ns_1_iv_0_0_a3_5[1]\ : NOR3
      port map(A => N_421, B => N_417, C => N_313_7_i, Y => 
        N_7176_i);
    
    un1_sstate_25_0_0_0_0 : OR2
      port map(A => N_7115_i, B => N_426, Y => 
        un1_sstate_25_0_0_0_0_i);
    
    un1_BYTECNT_3_I_47 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_1[0]\, B => 
        \CROMWAD[4]\, Y => \DWACT_ADD_CI_0_g_array_12_1_0[0]\);
    
    \SBYTE[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_12\, CLR => HWRES_c_31, 
        Q => \FBOUT[5]\);
    
    DACCfgValue_20 : MUX2H
      port map(A => \DACCfgValue[4]_net_1\, B => 
        \DACCfgValue_9[4]\, S => N_945, Y => \DACCfgValue_20\);
    
    \sstate_0[3]\ : DFFC
      port map(CLK => CLK_c_c, D => N_1022_i_0, CLR => 
        HWRES_c_32_0, Q => \sstate_0[3]_net_1\);
    
    \RESCNT_6_r[0]\ : OA21
      port map(A => N_313, B => \DWACT_ADD_CI_0_partial_sum_1[0]\, 
        C => N_528_i_0, Y => \RESCNT_6[0]\);
    
    \DACCfgValue[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_24\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[8]_net_1\);
    
    \SBYTE_7_1_i_a3_0[6]\ : NOR2FT
      port map(A => N_1075, B => \FBOUT[5]\, Y => N_331);
    
    un1_RESCNT_I_82 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11_1[0]\, B => 
        \RESCNT[10]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_4[0]\);
    
    DACCfgValue_26 : MUX2H
      port map(A => \DACCfgValue[10]_net_1\, B => 
        \DACCfgValue_9[10]\, S => N_945, Y => \DACCfgValue_26\);
    
    WRDACi : DFFS
      port map(CLK => CLK_c_c, D => \WRDACi_19\, SET => 
        HWRES_c_32, Q => \WRDACi\);
    
    \RESCNT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[4]\, CLR => 
        HWRES_c_30, Q => \RESCNT[4]_net_1\);
    
    \PAGECNT_9_0_a3[7]\ : AND2
      port map(A => N_436_i_0, B => I_34_0, Y => \PAGECNT_9[7]\);
    
    LUT : DFFC
      port map(CLK => CLK_c_c, D => \LUT_5_i_0\, CLR => 
        HWRES_c_27, Q => \LUT\);
    
    DACCfgValue_24 : MUX2H
      port map(A => \DACCfgValue[8]_net_1\, B => 
        \DACCfgValue_9[8]\, S => N_945, Y => \DACCfgValue_24\);
    
    \BYTECNT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[5]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[5]\);
    
    un1_pulse_3_0_0_0 : OR2FT
      port map(A => N_433, B => N_1078_1, Y => un1_pulse_3);
    
    \RELOAD_CNT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \RELOAD_CNT_3[4]\, CLR => 
        HWRES_c_29, Q => \REG[477]\);
    
    \BYTECNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[1]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[1]\);
    
    F_SO_maj_2_iv_0_0 : AO21
      port map(A => \F_SO_sync1\, B => \F_SO_sync2\, C => 
        \F_SO_sync\, Y => N_700);
    
    un1_sstate_26_0_0_i_a3 : NOR3
      port map(A => N_237, B => \sstate[1]_net_1\, C => 
        \sstate[0]_net_1\, Y => N_282);
    
    un1_BYTECNT_3_I_32 : XOR2
      port map(A => \CROMWAD[1]\, B => \DWACT_ADD_CI_0_TMP_1[0]\, 
        Y => I_32);
    
    \BYTECNT_9_0_a3[4]\ : AND2
      port map(A => N_437_i_0, B => I_30_0, Y => \BYTECNT_9[4]\);
    
    un1_RESCNT_I_51 : XOR2
      port map(A => \RESCNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_51);
    
    LUT_5_i_0_a2_0_1 : OR2
      port map(A => \PAGECNT_i_0_i[1]\, B => \PAGECNT[2]_net_1\, 
        Y => LUT_5_i_0_a2_0_1_i);
    
    un1_sstate_25_0_0_0 : NAND3FFT
      port map(A => un1_sstate_25_0_0_0_1_i, B => 
        un1_sstate_25_0_0_0_0_i, C => N_351, Y => 
        \un1_sstate_25_0_0_0\);
    
    \RESCNT_6_r[13]\ : OA21
      port map(A => N_313_0, B => I_60, C => N_528_i_0_0, Y => 
        \RESCNT_6[13]\);
    
    un1_BITCNT_I_1 : AND2
      port map(A => \BITCNT[0]_net_1\, B => \un1_sstate_25_0_0_0\, 
        Y => \DWACT_ADD_CI_0_TMP_2[0]\);
    
    \sstate_ns_1_iv_0_0_a3_1_1[1]\ : NAND2
      port map(A => \sstate[0]_net_1\, B => \sstate[2]_net_1\, Y
         => N_354_1);
    
    \PAGECNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[0]\, CLR => 
        HWRES_c_27_0, Q => \PAGECNT_i_i[0]\);
    
    un1_sstate_26_0_0_i_a3_0 : NOR2FT
      port map(A => N_1047, B => N_354_1, Y => N_283);
    
    \sstate_ns_1_iv_i_0_a3_4[2]\ : NOR2
      port map(A => N_413, B => N_414, Y => N_7181_i);
    
    un1_RESCNT_I_63 : XOR2
      port map(A => \RESCNT[8]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_3[0]\, Y => I_63);
    
    \sstate_ns_1_iv_0_0_0[1]\ : AO21TTF
      port map(A => N_420, B => N_423, C => 
        \sstate_ns_1_iv_0_0_a3_4[1]_net_1\, Y => 
        \sstate_ns_1_iv_0_0_0_i[1]\);
    
    \SBYTE_7_i_i_a2_0[0]\ : NOR2
      port map(A => N_394, B => N_1044, Y => N_1075);
    
    \WRCROM\ : DFFS
      port map(CLK => CLK_c_c, D => \WRCROMi\, SET => HWRES_c_32, 
        Q => WRCROM);
    
    F_SO_sync1_2_0_a2_0_a3 : NOR2FT
      port map(A => \F_SO_sync\, B => N_1078_0, Y => F_SO_sync1_2);
    
    \sstate_ns_1_iv_0_0_0_tz_0[0]\ : OAI21FTT
      port map(A => PULSE_10, B => N_427_1, C => N_392, Y => 
        \sstate_ns_1_iv_0_0_0_tz_0[0]_net_1\);
    
    \DACCfgValue_9_i_a3[10]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[10]_net_1\, Y => 
        N_273);
    
    DACCfgValue_22 : MUX2H
      port map(A => \DACCfgValue[6]_net_1\, B => 
        \DACCfgValue_9[6]\, S => N_945, Y => \DACCfgValue_22\);
    
    un1_sstate_25_0_0_0_o2 : NOR2FT
      port map(A => \sstate_0[1]_net_1\, B => N_1054, Y => N_1065);
    
    un1_ISI_1_sqmuxa_1_0_a3_0_1 : OR2
      port map(A => N_1050, B => \sstate_0[3]_net_1\, Y => 
        N_351_1);
    
    un1_ISCK_1_sqmuxa_i_0_0_a3 : AO21
      port map(A => N_406, B => N_417, C => N_1078, Y => 
        \un1_ISCK_1_sqmuxa_i_0_0_a3\);
    
    \SBYTE_7_1_i_a3_0[3]\ : NOR2FT
      port map(A => N_1075, B => \FBOUT[2]\, Y => N_327);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \sstate_ns_1_iv_i_a3[3]\ : OR3FFT
      port map(A => N_407, B => N_219, C => \sstate_0[0]_net_1\, 
        Y => N_289);
    
    \DACCFG_nWR\ : DFFS
      port map(CLK => CLK_c_c, D => \WRDACi\, SET => HWRES_c_25, 
        Q => DACCFG_nWR);
    
    \sstate_ns_1_iv_0_0_a2_1[1]\ : NOR2FT
      port map(A => \sstate_0[0]_net_1\, B => \sstate_0[2]_net_1\, 
        Y => N_423);
    
    \SBYTE_7_i_i_a3[2]\ : NOR2FT
      port map(A => REG_3, B => N_1046, Y => N_322_i);
    
    \RESCNT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[5]\, CLR => 
        HWRES_c_30, Q => \RESCNT[5]_net_1\);
    
    \PDLCFG_WDT_1[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[3]\, CLR => HWRES_c_28, 
        Q => CROMWDT(3));
    
    G_0_1 : OR2
      port map(A => \sstate_0[0]_net_1\, B => \sstate_0[3]_net_1\, 
        Y => G_0_1_i);
    
    \RESCNT_6_r[11]\ : OA21
      port map(A => N_313_0, B => I_56_1, C => N_528_i_0_0, Y => 
        \RESCNT_6[11]\);
    
    DACCfgValue_21 : MUX2H
      port map(A => \DACCfgValue[5]_net_1\, B => 
        \DACCfgValue_9[5]\, S => N_945, Y => \DACCfgValue_21\);
    
    un1_pulse_6_i_0_i_a2 : OR2
      port map(A => N_406, B => N_392, Y => N_418);
    
    N_400_1_i_i_i_o3_1 : NAND2FT
      port map(A => PULSE_0, B => PON_LOAD_i, Y => N_1078_1);
    
    \sstate_ns_1_iv_i_1[3]\ : NOR3FTT
      port map(A => N_293, B => N_1078_2, C => N_292_i, Y => 
        \sstate_ns_1_iv_i_1[3]_net_1\);
    
    \DACCfgValue_9_i_a3_0[7]\ : NOR2
      port map(A => \FBOUT[3]\, B => N_402, Y => N_268);
    
    \sstate_ns_1_iv_0_0_1[0]\ : AOI21TTF
      port map(A => N_420, B => N_1063, C => 
        \sstate_ns_1_iv_0_0_0[0]_net_1\, Y => 
        \sstate_ns_1_iv_0_0_1[0]_net_1\);
    
    \SBYTE[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_13\, CLR => HWRES_c_31, 
        Q => \FBOUT[6]\);
    
    \RESCNT[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[14]\, CLR => 
        HWRES_c_30, Q => \RESCNT[14]_net_1\);
    
    \DACCfgValue_9_i_a3[8]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[8]_net_1\, Y => 
        N_269);
    
    \sstate_ns_1_iv_i_a3_3[3]\ : OR2
      port map(A => \sstate_0[2]_net_1\, B => N_1038, Y => N_293);
    
    \BYTECNT_9_0_a3[8]\ : AND2
      port map(A => N_437_i_0, B => I_36, Y => \BYTECNT_9[8]\);
    
    un1_RESCNT_I_100 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_3[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_4[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2_1[0]\);
    
    un1_ISI_1_sqmuxa_1_0_1_0 : OR2FT
      port map(A => N_434, B => N_1078_1, Y => 
        un1_ISI_1_sqmuxa_1_0_1_0_i);
    
    \BITCNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_8[1]\, CLR => 
        HWRES_c_24, Q => \BITCNT[1]_net_1\);
    
    un1_ISCK_1_sqmuxa_i_0_0_2 : OAI21TTF
      port map(A => N_1074, B => N_247_i, C => N_348, Y => 
        un1_ISCK_1_sqmuxa_i_0_0_2_i);
    
    un1_ISCK_1_sqmuxa_i_0_0_a3_2 : NOR3FFT
      port map(A => \sstate_0[0]_net_1\, B => \sstate_0[4]_net_1\, 
        C => N_421, Y => N_348);
    
    \sstate_ns_0_0_0_a2[4]\ : NOR2
      port map(A => N_394, B => N_1078, Y => N_420);
    
    \RESCNT_6_r[4]\ : OA21
      port map(A => N_313, B => I_55, C => N_528_i_0, Y => 
        \RESCNT_6[4]\);
    
    \PAGECNT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[4]\, CLR => 
        HWRES_c_28, Q => \PAGECNT[4]_net_1\);
    
    un1_ISCK_1_sqmuxa_i_0_0_o2_1_0 : NAND2
      port map(A => \PAGECNT_i_0_i[1]\, B => \PAGECNT[2]_net_1\, 
        Y => un1_ISCK_1_sqmuxa_i_0_0_o2_1_i);
    
    un1_BYTECNT_3_I_49 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_1[0]\, B => 
        \CROMWAD[2]\, Y => \DWACT_ADD_CI_0_g_array_12_0[0]\);
    
    WRCROMi_0_sqmuxa_1_i_0_a2_0 : NOR2
      port map(A => \CROMWAD[8]\, B => N_395, Y => N_435);
    
    F_SO_sync_2_0_a2_0_a3 : NOR2FT
      port map(A => F_SO_c, B => N_1078_0, Y => F_SO_sync_2);
    
    \DACCfgValue[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_28\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[12]_net_1\);
    
    \RESCNT[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[9]\, CLR => 
        HWRES_c_31, Q => \RESCNT[9]_net_1\);
    
    WRCROMi : DFFS
      port map(CLK => CLK_c_c, D => \WRCROMi_17\, SET => 
        HWRES_c_32, Q => \WRCROMi\);
    
    un1_BYTECNT_3_I_46 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_2_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_3_1[0]\);
    
    ISI_8_iv_0_i_o2_0 : OR2FT
      port map(A => \sstate[2]_net_1\, B => REG_8, Y => N_235);
    
    un1_NCS0_2_sqmuxa_0_0_0 : NAND3
      port map(A => N_344, B => \un1_NCS0_2_sqmuxa_0_0_0_0\, C
         => N_410, Y => un1_NCS0_2_sqmuxa);
    
    \un1_drive_spi\ : OR2FT
      port map(A => \LOAD_RES\, B => REG_0, Y => un1_drive_spi);
    
    \sstate[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns[4]\, CLR => 
        HWRES_c_32_0, Q => \sstate[4]_net_1\);
    
    un1_sstate_26_0_0_i : NOR3
      port map(A => N_282, B => N_283, C => \sstate[3]_net_1\, Y
         => \un1_sstate_26_0_0_i\);
    
    \SBYTE_7_r[2]\ : OA21TTF
      port map(A => N_323_i, B => N_322_i, C => N_559, Y => 
        \SBYTE_7[2]\);
    
    \sstate_ns_1_iv_0_0_0[0]\ : OAI21TTF
      port map(A => \sstate_ns_1_iv_0_0_a3_4_1[0]_net_1\, B => 
        \sstate_ns_1_iv_0_0_0_tz_0[0]_net_1\, C => N_421, Y => 
        \sstate_ns_1_iv_0_0_0[0]_net_1\);
    
    \sstate_ns_1_iv_i_a2_i_0[3]\ : INV
      port map(A => \sstate[3]_net_1\, Y => \sstate_i_0[3]\);
    
    \sstate_0[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns[0]\, CLR => 
        HWRES_c_32_0, Q => \sstate_0[0]_net_1\);
    
    \RESCNT_6_0_a3_7_12[0]\ : OR3
      port map(A => \RESCNT_6_0_a3_7_10_i[0]\, B => 
        \RESCNT_6_0_a3_7_0_i[0]\, C => \RESCNT_6_0_a3_7_1_i[0]\, 
        Y => \RESCNT_6_0_a3_7_12_i[0]\);
    
    \SBYTE_7_i_i_a3[0]\ : NOR2FT
      port map(A => REG_1, B => N_1046, Y => N_318_i);
    
    \SBYTE[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_14\, CLR => HWRES_c_31, 
        Q => \FBOUT[7]\);
    
    un1_RESCNT_G_0 : AND3
      port map(A => \G\, B => \G_0_0\, C => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    LUT_5_i_0_o2 : NAND3
      port map(A => N_1065, B => N_1045, C => N_1062, Y => N_216);
    
    G_0 : OR3
      port map(A => N_1047, B => G_0_0_i, C => G_0_1_i, Y => 
        N_412);
    
    un1_PAGECNT_1_I_47 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \PAGECNT[4]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    un1_RESCNT_G_1_0 : NAND3
      port map(A => \DWACT_ADD_CI_0_pog_array_1[0]\, B => 
        \RESCNT[0]_net_1\, C => \RESCNT[1]_net_1\, Y => G_1_i);
    
    un1_PAGECNT_1_I_36 : XOR2
      port map(A => \PAGECNT[8]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_3_0[0]\, Y => I_36_0);
    
    \SBYTE_7_i_i_a3[4]\ : NOR2FT
      port map(A => REG_5, B => N_1046, Y => N_324_i);
    
    NCS0_15 : MUX2H
      port map(A => \NCS0\, B => NCS0_6, S => un1_NCS0_2_sqmuxa, 
        Y => \NCS0_15\);
    
    \DACCfgValue[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_23\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[7]_net_1\);
    
    \sstate_ns_1_iv_i_0_a3[2]\ : OAI21
      port map(A => N_1047, B => \sstate[3]_net_1\, C => N_423, Y
         => N_362);
    
    \SBYTE_7_r[7]\ : NOR3
      port map(A => N_559, B => N_334, C => N_332, Y => 
        \SBYTE_7[7]\);
    
    LUT_5_i_0_a2_0_0 : OR2
      port map(A => \PAGECNT_i_0_i[3]\, B => \PAGECNT[4]_net_1\, 
        Y => LUT_5_i_0_a2_0_0_i);
    
    COMMAND : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_3_i_0\, CLR => 
        HWRES_c_24, Q => \COMMAND\);
    
    \RESCNT[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[13]\, CLR => 
        HWRES_c_30, Q => \RESCNT[13]_net_1\);
    
    un1_ISCK_1_sqmuxa_i_0_0_a3_3 : NOR3FFT
      port map(A => \sstate[0]_net_1\, B => \N_414_i\, C => 
        N_1074, Y => N_349_i);
    
    RESCNT_1_sqmuxa_0_a2_0_a2_0_a3 : NOR2FT
      port map(A => PULSE_10, B => N_1078, Y => RESCNT_1_sqmuxa);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_45 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11_4[0]\, B => 
        \REG[479]\, Y => \DWACT_ADD_CI_0_g_array_12_2_2[0]\);
    
    WRDACi_19 : MUX2H
      port map(A => \WRDACi\, B => N_991, S => N_946, Y => 
        \WRDACi_19\);
    
    \sstate_ns_1_iv_0_0[1]\ : OR3
      port map(A => N_7179_i, B => N_353_i, C => 
        \sstate_ns_1_iv_0_0_3_i[1]\, Y => \sstate_ns[1]\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \sstate[3]\ : DFFC
      port map(CLK => CLK_c_c, D => N_1022_i_0, CLR => HWRES_c_32, 
        Q => \sstate[3]_net_1\);
    
    SBYTE_7 : MUX2H
      port map(A => \FBOUT[0]\, B => \SBYTE_7[0]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_7\);
    
    G_4 : OR3
      port map(A => \sstate_0[0]_net_1\, B => \sstate_0[3]_net_1\, 
        C => sstate_0_i_0(2), Y => N_1054);
    
    \DACCfgValue_9_i_a3[5]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[5]_net_1\, Y => 
        N_263);
    
    un1_PAGECNT_1_I_51 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_1_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_2_2[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2_0[0]\);
    
    \sstate_ns_1_iv_i_o2_3[3]\ : OR2
      port map(A => \CROMWAD[8]\, B => N_1040, Y => N_1041);
    
    \sstate_ns_1_iv_i_0_4[2]\ : NOR3
      port map(A => N_7181_i, B => \sstate_ns_1_iv_i_0_2_i[2]\, C
         => \sstate_ns_1_iv_i_0_1_i[2]\, Y => 
        \sstate_ns_1_iv_i_0_4[2]_net_1\);
    
    \sstate[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns[0]\, CLR => 
        HWRES_c_32, Q => \sstate[0]_net_1\);
    
    un1_NCS0_2_sqmuxa_0_0_0_a3_1 : NOR2
      port map(A => N_1038, B => N_1047, Y => N_343_1);
    
    N_400_1_i_i_i_o3_0 : NAND2FT
      port map(A => PULSE_0, B => PON_LOAD_i, Y => N_1078_0);
    
    DACCfgValue_29 : MUX2H
      port map(A => \DACCfgValue[13]_net_1\, B => N_1011, S => 
        N_945, Y => \DACCfgValue_29\);
    
    un1_ISCK_1_sqmuxa_i_0_0_a2_1 : OR2FT
      port map(A => N_407, B => N_1078_0, Y => N_421);
    
    \un1_BYTECNT_3_i_m_i_a3[1]\ : OR2
      port map(A => N_406, B => N_351_1, Y => N_312);
    
    \BYTECNT_9_0_a3[2]\ : AND2
      port map(A => N_437_i_0, B => I_35, Y => \BYTECNT_9[2]\);
    
    un1_RESCNT_I_92 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \RESCNT[4]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12_1_1[0]\);
    
    un1_LOAD_RESi_0_sqmuxa_0_0_0_a2 : OR2
      port map(A => N_1047, B => N_1054, Y => N_405);
    
    \sstate_ns_1_iv_0_0_a3_1[1]\ : AOI21FTT
      port map(A => N_382_i, B => N_1076, C => N_354_1, Y => 
        N_7179_i);
    
    DRIVE_RELOAD_2 : MUX2H
      port map(A => DRIVE_RELOAD_net_1, B => RESCNT_1_sqmuxa, S
         => un1_LOAD_RESi_0_sqmuxa, Y => \DRIVE_RELOAD_2\);
    
    \RESCNT_6_r_i_0[0]\ : NOR2FT
      port map(A => N_412, B => N_1078_0, Y => N_528_i_0_0);
    
    G : NAND2
      port map(A => N_412, B => N_425, Y => \G\);
    
    un1_FCS_SEL_0_sqmuxa_0_0_0 : NAND3FFT
      port map(A => N_281_i, B => N_280_i, C => N_528_i_0_0, Y
         => un1_FCS_SEL_0_sqmuxa);
    
    un1_RESCNT_I_86 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_10[0]\, B => 
        \RESCNT[12]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_5[0]\);
    
    \SBYTE_7_1_i_a3[7]\ : NOR2
      port map(A => N_1046, B => REG_8, Y => N_332);
    
    \DACCfgValue[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_25\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[9]_net_1\);
    
    \RESCNT_6_r[14]\ : OA21
      port map(A => N_313_0, B => I_65, C => N_528_i_0_0, Y => 
        \RESCNT_6[14]\);
    
    \sstate_ns_0_0_0_o2[4]\ : OR2
      port map(A => \sstate_0[2]_net_1\, B => \sstate_0[1]_net_1\, 
        Y => N_1039);
    
    un1_RESCNT_I_53 : XOR2
      port map(A => \RESCNT[10]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_11_1[0]\, Y => I_53);
    
    \RESCNT_6_r[1]\ : OA21
      port map(A => N_313, B => I_64, C => N_528_i_0, Y => 
        \RESCNT_6[1]\);
    
    un1_ISCK_1_sqmuxa_i_0_0_a3_1 : NOR3FTT
      port map(A => N_1058, B => N_1078_1, C => 
        un1_ISCK_1_sqmuxa_i_0_0_a3_1_0_i, Y => N_347_i);
    
    \RESCNT_6_0_a3_7_10[0]\ : NAND3
      port map(A => \RESCNT_6_0_a3_7_2[0]_net_1\, B => 
        \RESCNT[8]_net_1\, C => \RESCNT[9]_net_1\, Y => 
        \RESCNT_6_0_a3_7_10_i[0]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_32 : XOR2
      port map(A => \REG[475]\, B => 
        \DWACT_ADD_CI_0_g_array_1_3[0]\, Y => \RELOAD_CNT_3[2]\);
    
    un1_PAGECNT_1_I_54 : AND2
      port map(A => \PAGECNT[6]_net_1\, B => \PAGECNT_i_i[7]\, Y
         => \DWACT_ADD_CI_0_pog_array_1_2_2[0]\);
    
    un1_RESCNT_I_95 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_1_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_2_0[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2[0]\);
    
    un1_sstate_33_i_0_a2_1 : NOR2
      port map(A => \CROMWAD[6]\, B => N_1064, Y => N_384_i);
    
    \RESCNT[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[15]\, CLR => 
        HWRES_c_30, Q => \RESCNT[15]_net_1\);
    
    \BYTECNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[0]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[0]\);
    
    un1_BITCNT_I_14 : XOR2
      port map(A => \BITCNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, Y => I_14_0);
    
    \PAGECNT_9_0_a3[3]\ : AND2
      port map(A => N_436_i_0, B => I_37_0, Y => \PAGECNT_9[3]\);
    
    \BITCNT_8_r[1]\ : OA21
      port map(A => N_391, B => I_13_4, C => N_562, Y => 
        \BITCNT_8[1]\);
    
    \sstate_ns_1_iv_0_0_o2[0]\ : OR2FT
      port map(A => N_1039, B => N_424, Y => N_1063);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_47 : AND2
      port map(A => \REG[475]\, B => \REG[476]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\);
    
    \sstate_ns_0_0_0_a2_0[4]\ : NAND2
      port map(A => \sstate[3]_net_1\, B => \sstate[4]_net_1\, Y
         => N_394);
    
    WRCROMi_17 : MUX2H
      port map(A => \WRCROMi\, B => un1_pulse_1, S => N_943, Y
         => \WRCROMi_17\);
    
    \RESCNT_6_0_a3_7_2[0]\ : AND2
      port map(A => \RESCNT[10]_net_1\, B => \RESCNT[11]_net_1\, 
        Y => \RESCNT_6_0_a3_7_2[0]_net_1\);
    
    \DACCfgValue_9_r[6]\ : NOR3
      port map(A => N_1078_1, B => N_266, C => N_265, Y => 
        \DACCfgValue_9[6]\);
    
    un1_pulse_9_0_0_a2 : NOR3FTT
      port map(A => \sstate_0[2]_net_1\, B => N_409, C => N_1059, 
        Y => N_399);
    
    \sstate_ns_1_iv_0_0_a3_0[1]\ : NOR3FFT
      port map(A => \sstate_i_0[0]\, B => N_353_1, C => N_406, Y
         => N_353_i);
    
    un1_RESCNT_G_4_0 : NAND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_5[0]\, B => 
        \RESCNT[14]_net_1\, Y => G_4_0_i);
    
    \sstate_ns_0_0_0_a3_0[4]\ : NOR2
      port map(A => N_433, B => N_1078, Y => N_361);
    
    \BYTECNT_9_0_a3[6]\ : AND2
      port map(A => N_437_i_0, B => I_38_1, Y => \BYTECNT_9[6]\);
    
    \sstate[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns[1]\, CLR => 
        HWRES_c_32, Q => \sstate[1]_net_1\);
    
    F_SO_sync2_2_0_a2_0_a3 : NOR2FT
      port map(A => \F_SO_sync1\, B => N_1078_0, Y => 
        F_SO_sync2_2);
    
    \SBYTE[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_8\, CLR => HWRES_c_31, 
        Q => \FBOUT[1]\);
    
    DACCfgValue_28 : MUX2H
      port map(A => \DACCfgValue[12]_net_1\, B => N_1012, S => 
        N_945, Y => \DACCfgValue_28\);
    
    \PAGECNT_9_0_o2_1[8]\ : OA21FTF
      port map(A => N_419, B => N_414, C => N_1078, Y => N_436_1);
    
    \SBYTE_7_1_i_a3[5]\ : NOR2
      port map(A => N_1046, B => REG_6, Y => N_328);
    
    G_5 : OR2
      port map(A => \sstate_0[0]_net_1\, B => \sstate_0[3]_net_1\, 
        Y => N_1038);
    
    WRCROMi_0_sqmuxa_1_i_0_o3 : OAI21FTF
      port map(A => N_396_1, B => N_392, C => N_1078_2, Y => 
        un1_pulse_1);
    
    \RESCNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[2]\, CLR => 
        HWRES_c_30, Q => \RESCNT[2]_net_1\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_1 : AND2
      port map(A => \REG[473]\, B => un3_reload_edge, Y => 
        \DWACT_ADD_CI_0_TMP_3[0]\);
    
    un1_RESCNT_G_0_0 : AND2
      port map(A => \RESCNT[0]_net_1\, B => \RESCNT[1]_net_1\, Y
         => \G_0_0\);
    
    \RESCNT_6_0_a3_7_4[0]\ : AND2
      port map(A => \RESCNT[6]_net_1\, B => \RESCNT[7]_net_1\, Y
         => \RESCNT_6_0_a3_7_4[0]_net_1\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_33 : XOR2
      port map(A => \REG[478]\, B => 
        \DWACT_ADD_CI_0_g_array_12_1_2[0]\, Y => 
        \RELOAD_CNT_3[5]\);
    
    \DACCfgValue_9_r[4]\ : NOR3
      port map(A => N_1078_1, B => N_261, C => N_260, Y => 
        \DACCfgValue_9[4]\);
    
    \BYTECNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[2]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[2]\);
    
    un1_LOAD_RESi_1_sqmuxa_1_i_o2_0_0 : NOR2
      port map(A => N_218_i_i, B => N_419, Y => N_562);
    
    \sstate_ns_1_iv_0_0_a3_4_1[0]\ : NOR3FFT
      port map(A => N_390, B => \sstate_i_0[3]\, C => N_1053, Y
         => \sstate_ns_1_iv_0_0_a3_4_1[0]_net_1\);
    
    \PDLCFG_WDT_1[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[5]\, CLR => HWRES_c_28, 
        Q => CROMWDT(5));
    
    un1_ISCK_1_sqmuxa_i_0_0_o2_0 : NOR3
      port map(A => N_423, B => \sstate[1]_net_1\, C => 
        \sstate[3]_net_1\, Y => N_247_i);
    
    \RELOAD_CNT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \RELOAD_CNT_3[5]\, CLR => 
        HWRES_c_29, Q => \REG[478]\);
    
    \DACCfgValue_9_i_a3_0[10]\ : NOR2
      port map(A => \FBOUT[6]\, B => N_402, Y => N_274);
    
    \BITCNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_8[2]\, CLR => 
        HWRES_c_24, Q => \BITCNT[2]_net_1\);
    
    \RESCNT[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[11]\, CLR => 
        HWRES_c_30, Q => \RESCNT[11]_net_1\);
    
    \DACCfgValue[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_29\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[13]_net_1\);
    
    WRCROMi_0_sqmuxa_1_i_0_a3 : NOR3
      port map(A => N_395, B => N_1043, C => 
        \WRCROMi_0_sqmuxa_1_i_0_a3_0\, Y => N_315);
    
    un1_sstate_1_sqmuxa_0_0_0 : OAI21FTT
      port map(A => TICK(1), B => N_410, C => N_278, Y => 
        \un1_sstate_1_sqmuxa_0_0_0\);
    
    un1_LOAD_RESi_1_sqmuxa_1_i_o2_0_a2_0 : NOR2FT
      port map(A => N_7115_i, B => \sstate_0[4]_net_1\, Y => 
        N_415_i);
    
    \BITCNT_8_r[2]\ : OA21
      port map(A => N_391, B => I_14_0, C => N_562, Y => 
        \BITCNT_8[2]\);
    
    un1_RESCNT_I_98 : AND2
      port map(A => \RESCNT[2]_net_1\, B => \RESCNT[3]_net_1\, Y
         => \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    N_414_i : INV
      port map(A => N_414, Y => \N_414_i\);
    
    \DACCfgValue_9_i[12]\ : OA21TTF
      port map(A => \DACCfgValue[12]_net_1\, B => \FBOUT[0]\, C
         => N_991, Y => N_1012);
    
    un1_pulse_6_i_0_i : NOR3FFT
      port map(A => N_418, B => N_359, C => N_1078_1, Y => 
        N_1033_i);
    
    \RESCNT[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[7]\, CLR => 
        HWRES_c_31, Q => \RESCNT[7]_net_1\);
    
    F_SO_maj_2_r : NOR3FFT
      port map(A => N_342, B => N_700, C => N_1078_0, Y => 
        F_SO_maj_2);
    
    un1_PAGECNT_1_I_49 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_0[0]\, B => 
        \PAGECNT[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    un1_BYTECNT_3_I_53 : AND2
      port map(A => \CROMWAD[4]\, B => \CROMWAD[5]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1_2[0]\);
    
    N_400_1_i_i_i_o3_2 : NAND2FT
      port map(A => PULSE_0, B => PON_LOAD_i, Y => N_1078_2);
    
    un1_BYTECNT_3_I_51 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_1_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_2_1[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2_2[0]\);
    
    \sstate_ns_1_iv_0_0_a3_2_0[1]\ : NOR3
      port map(A => \sstate_ns_1_iv_0_0_a3_0_i[1]\, B => N_1053, 
        C => N_1078_2, Y => \sstate_ns_1_iv_0_0_a3_2[1]_net_1\);
    
    \PAGECNT_9_0_a3[2]\ : AND2
      port map(A => N_436_i_0, B => I_35_0, Y => \PAGECNT_9[2]\);
    
    \PAGECNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[2]\, CLR => 
        HWRES_c_27_0, Q => \PAGECNT[2]_net_1\);
    
    un1_pulse_9_0_0 : NOR3FTT
      port map(A => N_434, B => \un1_pulse_9_0_0_0\, C => N_399, 
        Y => un1_pulse_9);
    
    un1_PAGECNT_1_I_44 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_0[0]\, B => 
        \PAGECNT_i_0_i[1]\, Y => \DWACT_ADD_CI_0_g_array_1_0[0]\);
    
    un1_BYTECNT_3_I_44 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_1[0]\, B => \CROMWAD[1]\, 
        Y => \DWACT_ADD_CI_0_g_array_1_1[0]\);
    
    \sstate_ns_1_iv_i_0_0[2]\ : AOI21
      port map(A => N_416, B => N_396_1, C => N_1078_2, Y => 
        \sstate_ns_1_iv_i_0_0[2]_net_1\);
    
    \PAGECNT[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[7]\, CLR => 
        HWRES_c_28, Q => \PAGECNT_i_i[7]\);
    
    \BYTECNT[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[7]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[7]\);
    
    un1_pulse_9_0_0_a2_2 : NOR3FTT
      port map(A => \sstate_0[1]_net_1\, B => N_1038, C => N_1041, 
        Y => N_398);
    
    \sstate_ns_1_iv_0_0_2[0]\ : OAI21FTT
      port map(A => \sstate_ns_1_iv_0_0_a3_3_0[0]_net_1\, B => 
        N_1074, C => \sstate_ns_1_iv_0_0_1[0]_net_1\, Y => 
        \sstate_ns_1_iv_0_0_2_i[0]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_30 : XOR2
      port map(A => \REG[476]\, B => 
        \DWACT_ADD_CI_0_g_array_12_6[0]\, Y => \RELOAD_CNT_3[3]\);
    
    un1_RESCNT_I_78 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11[0]\, B => 
        \RESCNT[6]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12_2_1[0]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_27 : XOR2
      port map(A => \REG[479]\, B => 
        \DWACT_ADD_CI_0_g_array_11_4[0]\, Y => \RELOAD_CNT_3[6]\);
    
    un1_SBYTE_0_sqmuxa_0_0_0_a2 : NOR2FT
      port map(A => \sstate[4]_net_1\, B => N_1044, Y => N_432);
    
    un1_FCS_SEL_0_sqmuxa_0_0_a2_i_1 : INV
      port map(A => N_1047, Y => N_1047_i_0);
    
    \sstate_ns_1_iv_i_0_2[2]\ : AO21TTF
      port map(A => N_426, B => \sstate[1]_net_1\, C => N_362, Y
         => \sstate_ns_1_iv_i_0_2_i[2]\);
    
    ISI_8_iv_0_i_m3 : MUX2H
      port map(A => N_235, B => \FBOUT[7]\, S => 
        \sstate[4]_net_1\, Y => N_248);
    
    un1_RESCNT_I_57 : XOR2
      port map(A => \RESCNT[5]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_1_1[0]\, Y => I_57);
    
    \sstate_ns_1_iv_i_a2[3]\ : OR2FT
      port map(A => \sstate_0[0]_net_1\, B => \sstate_0[3]_net_1\, 
        Y => N_392);
    
    \PAGECNT[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[8]\, CLR => 
        HWRES_c_28, Q => \PAGECNT[8]_net_1\);
    
    \RESCNT_6_0_a3_7_6[0]\ : AND2
      port map(A => \RESCNT[2]_net_1\, B => \RESCNT[3]_net_1\, Y
         => \RESCNT_6_0_a3_7_6[0]_net_1\);
    
    ISI_8_iv_0_i_o2 : NAND3
      port map(A => \sstate[4]_net_1\, B => \ISI_8_iv_0_i_o2_0\, 
        C => \BITCNT[0]_net_1\, Y => N_1053);
    
    \DACCFG_WDT_1[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[5]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(5));
    
    \DACCFG_WDT_1[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[10]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(10));
    
    un1_BYTECNT_3_I_21 : XOR2
      port map(A => \CROMWAD[0]\, B => \un1_sstate_26_0_0_i\, Y
         => \DWACT_ADD_CI_0_partial_sum[0]\);
    
    un1_RESCNT_G_5 : XOR2
      port map(A => \RESCNT[15]_net_1\, B => \G_4\, Y => \G_5\);
    
    NCS0_6_s : OAI21FTT
      port map(A => FWIMG2LOAD, B => N_412, C => N_1033_i, Y => 
        NCS0_6);
    
    \DACCfgValue[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_21\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[5]_net_1\);
    
    RELOAD_EDGE_i : INV
      port map(A => \RELOAD_EDGE\, Y => \RELOAD_EDGE_i\);
    
    un1_RESCNT_G_4 : AND3FFT
      port map(A => G_4_4_i, B => G_4_3_i, C => \G\, Y => \G_4\);
    
    un1_PAGECNT_1_I_35 : XOR2
      port map(A => \PAGECNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, Y => I_35_0);
    
    \PDLCFG_WDT_1[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[6]\, CLR => HWRES_c_28, 
        Q => CROMWDT(6));
    
    un1_RESCNT_G_2_5 : NAND2
      port map(A => \DWACT_ADD_CI_0_pog_array_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_2_1[0]\, Y => G_2_i);
    
    un1_ISCK_1_sqmuxa_i_0_0_a2 : OR2FT
      port map(A => N_416, B => N_1078_0, Y => N_422);
    
    \sstate_ns_1_iv_i_3[3]\ : OAI21FTT
      port map(A => N_343_1, B => PULSE_6, C => 
        \sstate_ns_1_iv_i_1[3]_net_1\, Y => 
        \sstate_ns_1_iv_i_3_i[3]\);
    
    \DACCfgValue_9_i_a3[11]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[11]_net_1\, Y => 
        N_275);
    
    un1_RESCNT_I_94 : AND2
      port map(A => \RESCNT[8]_net_1\, B => \RESCNT[9]_net_1\, Y
         => \DWACT_ADD_CI_0_pog_array_1_3[0]\);
    
    un1_ISI_1_sqmuxa_1_0_1 : NAND3FFT
      port map(A => un1_ISI_1_sqmuxa_1_0_1_0_i, B => N_350_i, C
         => N_351, Y => un1_ISI_1_sqmuxa_1);
    
    \DACCfgValue_9_i[13]\ : OA21TTF
      port map(A => \DACCfgValue[13]_net_1\, B => \FBOUT[1]\, C
         => N_991, Y => N_1011);
    
    \BYTECNT_9_0_a3[1]\ : AND2
      port map(A => N_437_i_0, B => I_32, Y => \BYTECNT_9[1]\);
    
    \RELOAD_CNT[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \RELOAD_CNT_3[6]\, CLR => 
        HWRES_c_29, Q => \REG[479]\);
    
    un1_RESCNT_I_70 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_3[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_1[0]\);
    
    un1_LOAD_RESi_0_sqmuxa_0_0_0 : OR2FT
      port map(A => N_405, B => N_1078_0, Y => 
        un1_LOAD_RESi_0_sqmuxa);
    
    \RESCNT_6_r[5]\ : OA21
      port map(A => N_313, B => I_57, C => N_528_i_0, Y => 
        \RESCNT_6[5]\);
    
    \sstate_ns_1_iv_0_0_a2_0[1]\ : OR2FT
      port map(A => \sstate[4]_net_1\, B => N_392, Y => N_417);
    
    \RESCNT_6_r[2]\ : OA21
      port map(A => N_313, B => I_51, C => N_528_i_0, Y => 
        \RESCNT_6[2]\);
    
    un1_BYTECNT_3_I_42 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_3[0]\);
    
    \DACCFG_WDT_1[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[12]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(12));
    
    \sstate_ns_1_iv_0_0_3[0]\ : OAI21
      port map(A => N_1074, B => N_434, C => 
        \sstate_ns_1_iv_0_0_a3_1[0]_net_1\, Y => 
        \sstate_ns_1_iv_0_0_3_i[0]\);
    
    \SBYTE[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_7\, CLR => HWRES_c_31, 
        Q => \FBOUT[0]\);
    
    WRPDLi_0_sqmuxa_1_i_0_a3_1 : NOR3FFT
      port map(A => \CROMWAD_i_0[7]\, B => N_1064, C => 
        \CROMWAD[6]\, Y => \WRPDLi_0_sqmuxa_1_i_0_a3_1\);
    
    \RESCNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[0]\, CLR => 
        HWRES_c_30, Q => \RESCNT[0]_net_1\);
    
    \PAGECNT_9_0_a3[8]\ : AND2
      port map(A => N_436_i_0, B => I_36_0, Y => \PAGECNT_9[8]\);
    
    un1_PAGECNT_1_I_30 : XOR2
      port map(A => \PAGECNT[4]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\, Y => I_30_1);
    
    DACCfgValue_25 : MUX2H
      port map(A => \DACCfgValue[9]_net_1\, B => 
        \DACCfgValue_9[9]\, S => N_945, Y => \DACCfgValue_25\);
    
    \sstate_ns_1_iv_0_0_a2[0]\ : NOR2FT
      port map(A => \LUT\, B => \COMMAND\, Y => N_390);
    
    un1_RESCNT_I_74 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \RESCNT[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_3[0]\);
    
    un1_sstate_33_i_0 : OR2FT
      port map(A => N_317, B => N_1078_1, Y => N_945);
    
    \sstate_ns_0_0_0_0[4]\ : OAI21TTF
      port map(A => N_422, B => N_1039, C => N_420, Y => 
        \sstate_ns_0_0_0_0[4]_net_1\);
    
    un1_ISCK_1_sqmuxa_i_0_0_o2 : NAND3FFT
      port map(A => un1_ISCK_1_sqmuxa_i_0_0_o2_0_i, B => 
        un1_ISCK_1_sqmuxa_i_0_0_o2_1_i, C => N_143_i_0, Y => 
        N_1058);
    
    \RESCNT_6_r[12]\ : OA21
      port map(A => N_313_0, B => I_58, C => N_528_i_0_0, Y => 
        \RESCNT_6[12]\);
    
    \SBYTE_7_r[0]\ : OA21TTF
      port map(A => N_319_i, B => N_318_i, C => N_559, Y => 
        \SBYTE_7[0]\);
    
    \DACCfgValue_9_i_a3_0[9]\ : NOR2
      port map(A => \FBOUT[5]\, B => N_402, Y => N_272);
    
    un1_PAGECNT_1_I_38 : XOR2
      port map(A => \PAGECNT[6]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_11_0[0]\, Y => I_38_2);
    
    un1_BYTECNT_3_I_35 : XOR2
      port map(A => \CROMWAD[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, Y => I_35);
    
    \DACCfgValue_9_i_a3_0[6]\ : NOR2
      port map(A => \FBOUT[2]\, B => N_402, Y => N_266);
    
    un1_ISCK_1_sqmuxa_i_0_0_a3_1_0 : OR2
      port map(A => \sstate_0[2]_net_1\, B => \sstate_0[0]_net_1\, 
        Y => un1_ISCK_1_sqmuxa_i_0_0_a3_1_0_i);
    
    \SBYTE_7_i_i_a3_0[0]\ : AND2
      port map(A => \F_SO_maj\, B => N_1075, Y => N_319_i);
    
    DACCfgValue_23 : MUX2H
      port map(A => \DACCfgValue[7]_net_1\, B => 
        \DACCfgValue_9[7]\, S => N_945, Y => \DACCfgValue_23\);
    
    un1_NCS0_2_sqmuxa_0_0_0_0 : AOI21
      port map(A => PULSE_10, B => N_343_1, C => N_1078_1, Y => 
        \un1_NCS0_2_sqmuxa_0_0_0_0\);
    
    un1_sstate_33_i_0_a2_0 : AND2
      port map(A => \CROMWAD[6]\, B => N_1042, Y => N_383_i);
    
    LOAD_RESi_1 : MUX2H
      port map(A => \LOAD_RES\, B => N_1078_i_0, S => 
        un1_LOAD_RESi_0_sqmuxa, Y => \LOAD_RESi_1\);
    
    \DACCFG_WDT_1[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[11]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(11));
    
    \DACCfgValue_9_r[8]\ : NOR3
      port map(A => N_1078_2, B => N_270, C => N_269, Y => 
        \DACCfgValue_9[8]\);
    
    un1_PAGECNT_1_I_21 : XOR2
      port map(A => \PAGECNT_i_i[0]\, B => 
        \un1_sstate_1_sqmuxa_0_0_0\, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\);
    
    \RESCNT[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[6]\, CLR => 
        HWRES_c_31, Q => \RESCNT[6]_net_1\);
    
    \PDLCFG_WDT_1[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[4]\, CLR => HWRES_c_28, 
        Q => CROMWDT(4));
    
    un1_pulse_7_0_0_0_o3 : OR2
      port map(A => N_1065, B => N_1078_2, Y => N_559);
    
    un1_sstate_25_0_0_0_a2 : NOR2FT
      port map(A => \sstate_0[4]_net_1\, B => N_1038, Y => N_426);
    
    un1_RESCNT_I_96 : AND2
      port map(A => \RESCNT[4]_net_1\, B => \RESCNT[5]_net_1\, Y
         => \DWACT_ADD_CI_0_pog_array_1_1_0[0]\);
    
    \SBYTE_7_r[5]\ : NOR3
      port map(A => N_559, B => N_329, C => N_328, Y => 
        \SBYTE_7[5]\);
    
    \SBYTE_7_r[1]\ : OA21TTF
      port map(A => N_321_i, B => N_320_i, C => N_559, Y => 
        \SBYTE_7[1]\);
    
    \DRIVE_RELOAD\ : DFFC
      port map(CLK => CLK_c_c, D => \DRIVE_RELOAD_2\, CLR => 
        HWRES_c_26, Q => DRIVE_RELOAD_net_1);
    
    un1_BYTECNT_3_I_1 : AND2
      port map(A => \CROMWAD[0]\, B => \un1_sstate_26_0_0_i\, Y
         => \DWACT_ADD_CI_0_TMP_1[0]\);
    
    DACCfgValue_27 : MUX2H
      port map(A => \DACCfgValue[11]_net_1\, B => 
        \DACCfgValue_9[11]\, S => N_945, Y => \DACCfgValue_27\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_48 : AND2
      port map(A => \REG[477]\, B => \REG[478]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1_3[0]\);
    
    LOAD_RESi : DFFS
      port map(CLK => CLK_c_c, D => \LOAD_RESi_1\, SET => 
        HWRES_c_27, Q => \LOAD_RES\);
    
    un1_pulse_9_0_0_a2_3 : NAND2FT
      port map(A => N_1043, B => N_1062, Y => N_409);
    
    \sstate_ns_1_iv_0_0_a3_2[1]\ : OR2FT
      port map(A => \sstate_0[1]_net_1\, B => N_422, Y => 
        \sstate_ns_1_iv_0_0_a3_2_0[1]_net_1\);
    
    \RESCNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[3]\, CLR => 
        HWRES_c_30, Q => \RESCNT[3]_net_1\);
    
    \sstate_ns_1_iv_0_0_a3_0_0[1]\ : OAI21TTF
      port map(A => \COMMAND\, B => \LUT\, C => 
        \sstate_0[1]_net_1\, Y => \sstate_ns_1_iv_0_0_a3_0_i[1]\);
    
    \sstate_ns_1_iv_0_0_1[1]\ : OAI21FTT
      port map(A => \sstate_ns_1_iv_0_0_a3_2[1]_net_1\, B => 
        N_1054, C => \sstate_ns_1_iv_0_0_a3_2_0[1]_net_1\, Y => 
        \sstate_ns_1_iv_0_0_1_i[1]\);
    
    un1_LOAD_RESi_1_sqmuxa_1_i_o2_0_0_o3 : OR3FTT
      port map(A => N_351, B => N_559, C => N_415_i, Y => 
        N_218_i_i);
    
    \sstate_ns_1_iv_i[3]\ : OA21FTT
      port map(A => N_363_1, B => \sstate_0[3]_net_1\, C => 
        \sstate_ns_1_iv_i_5[3]_net_1\, Y => N_1022_i_0);
    
    \RESCNT_6_0_a3_0[0]\ : NOR2
      port map(A => N_313_7_i, B => N_425, Y => N_313_0);
    
    \DACCfgValue_9_r[5]\ : NOR3
      port map(A => N_1078_1, B => N_264, C => N_263, Y => 
        \DACCfgValue_9[5]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_19 : XOR2
      port map(A => \REG[473]\, B => un3_reload_edge, Y => 
        \DWACT_ADD_CI_0_partial_sum_3[0]\);
    
    \PAGECNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[1]\, CLR => 
        HWRES_c_27_0, Q => \PAGECNT_i_0_i[1]\);
    
    \DACCFG_WDT_1[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[13]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(13));
    
    WRCROMi_0_sqmuxa_1_i_0_o2 : OR2FT
      port map(A => N_1042, B => \CROMWAD[6]\, Y => N_1043);
    
    un1_SBYTE_0_sqmuxa_0_0_0 : OR2
      port map(A => N_218_i_i, B => N_432, Y => 
        un1_SBYTE_0_sqmuxa);
    
    un1_pulse_7_0_0_0_a2 : OR2
      port map(A => N_410, B => N_1058, Y => N_434);
    
    WRPDLi_0_sqmuxa_1_i_0 : AO21
      port map(A => \WRPDLi_0_sqmuxa_1_i_0_a3_1\, B => N_435, C
         => un1_pulse_1, Y => N_944);
    
    un1_PAGECNT_1_I_33 : XOR2
      port map(A => \PAGECNT_i_i[5]\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => I_33_0);
    
    \DACCfgValue_9_i_a3_0[5]\ : NOR2
      port map(A => \FBOUT[1]\, B => N_402, Y => N_264);
    
    un1_PAGECNT_1_I_32 : XOR2
      port map(A => \PAGECNT_i_0_i[1]\, B => 
        \DWACT_ADD_CI_0_TMP_0[0]\, Y => I_32_0);
    
    un1_RESCNT_G_3 : AND3
      port map(A => \G\, B => \RESCNT[0]_net_1\, C => 
        \RESCNT[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \SBYTE_7_i_i_a3_0[2]\ : AND2
      port map(A => \FBOUT[1]\, B => N_1075, Y => N_323_i);
    
    \sstate_ns_1_iv_i_0_a3_0_1[2]\ : NOR2FT
      port map(A => N_1050, B => \sstate[2]_net_1\, Y => N_363_1);
    
    RELOAD_EDGE_r : DFFS
      port map(CLK => CLK_c_c, D => \RELOAD_EDGE_i\, SET => 
        HWRES_c_29, Q => RELOAD_EDGE_r_i_0);
    
    \PAGECNT_9_0_a3[4]\ : AND2
      port map(A => N_436_i_0, B => I_30_1, Y => \PAGECNT_9[4]\);
    
    un1_RESCNT_I_65 : XOR2
      port map(A => \RESCNT[14]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_11_2[0]\, Y => I_65);
    
    un1_pulse_9_0_0_0 : OAI21TTF
      port map(A => N_1050, B => \un1_pulse_9_0_0_a2_0_0\, C => 
        N_1078, Y => \un1_pulse_9_0_0_0\);
    
    LOAD_RESi_1_0 : DFFS
      port map(CLK => CLK_c_c, D => \LOAD_RESi_1\, SET => 
        HWRES_c_27_0, Q => LOAD_RES_1);
    
    \DACCfgValue_9_i_a3[7]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[7]_net_1\, Y => 
        N_267);
    
    \RESCNT_6_0_a3_7_1[0]\ : NAND2
      port map(A => \RESCNT[12]_net_1\, B => \RESCNT[13]_net_1\, 
        Y => \RESCNT_6_0_a3_7_1_i[0]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_36 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_3[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_2[0]\);
    
    \RELOAD_CNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => 
        \DWACT_ADD_CI_0_partial_sum_3[0]\, CLR => HWRES_c_29, Q
         => \REG[473]\);
    
    un1_sstate_33_i_0_a3 : OR3
      port map(A => N_401, B => \CROMWAD[7]\, C => \CROMWAD[8]\, 
        Y => N_317);
    
    un1_pulse_9_0_0_a2_0_0 : OR2
      port map(A => N_392, B => \sstate[2]_net_1\, Y => 
        \un1_pulse_9_0_0_a2_0_0\);
    
    \DACCFG_WDT_1[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[6]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(6));
    
    WRDACi_0_sqmuxa_1_i_0 : OR2FT
      port map(A => N_317, B => un1_pulse_1, Y => N_946);
    
    un1_BYTECNT_3_I_50 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11_3[0]\, B => 
        \CROMWAD[6]\, Y => \DWACT_ADD_CI_0_g_array_12_2_0[0]\);
    
    \SBYTE_7_i_i_a3[1]\ : NOR2FT
      port map(A => REG_2, B => N_1046, Y => N_320_i);
    
    \RESCNT[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[10]\, CLR => 
        HWRES_c_30, Q => \RESCNT[10]_net_1\);
    
    \PDLCFG_nWR\ : DFFS
      port map(CLK => CLK_c_c, D => \WRPDLi\, SET => HWRES_c_29, 
        Q => PDLCFG_nWR);
    
    \RESCNT_6_r[8]\ : OA21
      port map(A => N_313_0, B => I_63, C => N_528_i_0_0, Y => 
        \RESCNT_6[8]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_34 : XOR2
      port map(A => \REG[480]\, B => 
        \DWACT_ADD_CI_0_g_array_12_2_2[0]\, Y => 
        \RELOAD_CNT_3[7]\);
    
    G_3 : OA21
      port map(A => N_313_0, B => \G_5\, C => N_528_i_0_0, Y => 
        \RESCNT_6[15]\);
    
    \DACCfgValue_9_i_a3_0[8]\ : NOR2
      port map(A => \FBOUT[4]\, B => N_402, Y => N_270);
    
    un1_RESCNT_G_4_4 : NAND3FTT
      port map(A => G_4_0_i, B => \DWACT_ADD_CI_0_pog_array_2[0]\, 
        C => \DWACT_ADD_CI_0_pog_array_1[0]\, Y => G_4_4_i);
    
    \PAGECNT_9_0_o2[8]\ : AND3
      port map(A => N_436_1, B => N_216, C => N_434, Y => 
        N_436_i_0);
    
    ISCK_4 : MUX2H
      port map(A => sstate_26_sqmuxa, B => ISCK_net_1, S => N_498, 
        Y => \ISCK_4\);
    
    un1_ISCK_1_sqmuxa_i_0_0 : OR3
      port map(A => N_349_i, B => un1_ISCK_1_sqmuxa_i_0_0_2_i, C
         => un1_ISCK_1_sqmuxa_i_0_0_1_i, Y => N_498);
    
    un1_BYTECNT_3_I_33 : XOR2
      port map(A => \CROMWAD[5]\, B => 
        \DWACT_ADD_CI_0_g_array_12_1_0[0]\, Y => I_33);
    
    \sstate_ns_1_iv_i_a3_5[3]\ : NOR2
      port map(A => N_414, B => N_392, Y => N_295_i);
    
    ISI_8_iv_0_i_o3_i_0 : INV
      port map(A => \sstate[0]_net_1\, Y => \sstate_i_0[0]\);
    
    un1_sstate_26_0_0_i_o2 : OR2
      port map(A => \sstate_0[4]_net_1\, B => \sstate[1]_net_1\, 
        Y => N_1047);
    
    WRDACi_7_i_a2_0_a3 : OR2FT
      port map(A => N_402_0, B => N_1078_1, Y => N_991);
    
    \sstate_ns_1_iv_i_o2_0_0[3]\ : NOR2
      port map(A => \CROMWAD[2]\, B => \CROMWAD[1]\, Y => 
        \sstate_ns_1_iv_i_o2_0[3]_net_1\);
    
    \sstate_0[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns[1]\, CLR => 
        HWRES_c_32_0, Q => \sstate_0[1]_net_1\);
    
    \RESCNT[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[8]\, CLR => 
        HWRES_c_31, Q => \RESCNT[8]_net_1\);
    
    NCS0 : DFFS
      port map(CLK => CLK_c_c, D => \NCS0_15\, SET => HWRES_c_27, 
        Q => \NCS0\);
    
    \DACCfgValue_9_i_a3[6]\ : NOR2FT
      port map(A => N_402_0, B => \DACCfgValue[6]_net_1\, Y => 
        N_265);
    
    \PAGECNT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[5]\, CLR => 
        HWRES_c_28, Q => \PAGECNT_i_i[5]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_28 : XOR2
      port map(A => \REG[477]\, B => 
        \DWACT_ADD_CI_0_g_array_2_2[0]\, Y => \RELOAD_CNT_3[4]\);
    
    un1_RESCNT_I_91 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_3[0]\, B => 
        \RESCNT[8]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12_3_0[0]\);
    
    \sstate[2]\ : DFFS
      port map(CLK => CLK_c_c, D => N_846_i_0, SET => HWRES_c_32, 
        Q => \sstate[2]_net_1\);
    
    \SBYTE_7_i_i_a3_0[1]\ : AND2
      port map(A => \FBOUT[0]\, B => N_1075, Y => N_321_i);
    
    un1_sstate_25_0_0_a2_0 : NOR2FT
      port map(A => PULSE_6, B => N_1054, Y => N_7115_i);
    
    \sstate_ns_1_iv_i_0_a2_0[2]\ : NOR2FT
      port map(A => \sstate_0[3]_net_1\, B => \sstate[0]_net_1\, 
        Y => N_416);
    
    \ISI\ : DFFC
      port map(CLK => CLK_c_c, D => \ISI_16\, CLR => HWRES_c_27, 
        Q => ISI_net_1);
    
    un1_RESCNT_G_1_1 : AND3
      port map(A => \DWACT_ADD_CI_0_pog_array_1[0]\, B => 
        \RESCNT[0]_net_1\, C => \RESCNT[1]_net_1\, Y => G_1_1);
    
    un1_pulse_7_0_0_0_o2_i : INV
      port map(A => N_1038, Y => N_1038_i_0);
    
    \sstate_ns_1_iv_i_o2[3]\ : NAND3
      port map(A => N_1045, B => \sstate_ns_1_iv_i_o2_0[3]_net_1\, 
        C => \CROMWAD[3]\, Y => N_1050);
    
    \BYTECNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[3]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[3]\);
    
    \sstate_ns_1_iv_0_0_a3_2[0]\ : NOR2FT
      port map(A => N_353_1, B => N_392, Y => N_373_i);
    
    un1_RESCNT_G_2_2 : NAND2
      port map(A => \DWACT_ADD_CI_0_pog_array_2_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => G_2_2_i);
    
    un1_NCS0_2_sqmuxa_0_0_0_a2 : OR2
      port map(A => N_1039, B => N_1038, Y => N_410);
    
    \SBYTE_7_1_i_a3_0[7]\ : NOR2FT
      port map(A => N_1075, B => \FBOUT[6]\, Y => N_334);
    
    LUT_5_i_0 : AOI21FTF
      port map(A => \LUT\, B => N_216, C => N_436_1, Y => 
        \LUT_5_i_0\);
    
    un1_sstate_1_sqmuxa_0_0_0_a2 : NOR2
      port map(A => N_408, B => N_409, Y => N_411);
    
    un1_ISI_1_sqmuxa_1_0_1_o2 : OR2FT
      port map(A => \sstate[0]_net_1\, B => N_1039, Y => N_1044);
    
    \PAGECNT_9_0_a3[5]\ : AND2
      port map(A => N_436_i_0, B => I_33_0, Y => \PAGECNT_9[5]\);
    
    \BYTECNT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[4]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[4]\);
    
    \un1_BITCNT_i_m_i_s_0_a2[1]\ : NOR2
      port map(A => N_1053, B => N_1038, Y => N_391);
    
    un1_BYTECNT_3_I_37 : XOR2
      port map(A => \CROMWAD[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, Y => I_37);
    
    un1_RESCNT_G_4_3 : NAND3
      port map(A => \DWACT_ADD_CI_0_pog_array_2_1[0]\, B => 
        \RESCNT[0]_net_1\, C => \RESCNT[1]_net_1\, Y => G_4_3_i);
    
    un1_ISCK_1_sqmuxa_i_0_0_a2_0 : OR2
      port map(A => \sstate_0[4]_net_1\, B => N_1078, Y => N_1074);
    
    un1_BITCNT_I_15 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_2[0]\, B => 
        \BITCNT[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1_2[0]\);
    
    \sstate_ns_1_iv_0_0_a2_1_1[0]\ : OR2
      port map(A => PULSE_6, B => \sstate[4]_net_1\, Y => N_427_1);
    
    \PAGECNT[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[6]\, CLR => 
        HWRES_c_28, Q => \PAGECNT[6]_net_1\);
    
    WRCROMi_0_sqmuxa_1_i_0_a2_1_0 : NOR2FT
      port map(A => \sstate_0[1]_net_1\, B => \sstate_0[4]_net_1\, 
        Y => N_396_1);
    
    WRCROMi_0_sqmuxa_1_i_0_o2_0 : NOR2
      port map(A => \CROMWAD[4]\, B => \CROMWAD[5]\, Y => N_1042);
    
    un1_RESCNT_I_60 : XOR2
      port map(A => \RESCNT[13]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_5[0]\, Y => I_60);
    
    un1_RESCNT_I_40 : XOR2
      port map(A => \RESCNT[0]_net_1\, B => \G\, Y => 
        \DWACT_ADD_CI_0_partial_sum_1[0]\);
    
    un1_PAGECNT_1_I_46 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_2_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_3_0[0]\);
    
    un1_pulse_3_0_0_0_a2 : OR2
      port map(A => N_412, B => PULSE_6, Y => N_433);
    
    un1_BYTECNT_3_I_38 : XOR2
      port map(A => \CROMWAD[6]\, B => 
        \DWACT_ADD_CI_0_g_array_11_3[0]\, Y => I_38_1);
    
    LOAD_RESi_0 : DFFS
      port map(CLK => CLK_c_c, D => \LOAD_RESi_1\, SET => 
        HWRES_c_27_0, Q => LOAD_RES_0);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_42 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_2[0]\, B => 
        \REG[477]\, Y => \DWACT_ADD_CI_0_g_array_12_1_2[0]\);
    
    \PAGECNT_9_0_a3[0]\ : AND2
      port map(A => N_436_i_0, B => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, Y => \PAGECNT_9[0]\);
    
    \RESCNT_6_0_a3_7[0]\ : OR3
      port map(A => \RESCNT_6_0_a3_7_12_i[0]\, B => 
        \RESCNT_6_0_a3_7_8_i[0]\, C => \RESCNT_6_0_a3_7_9_i[0]\, 
        Y => N_313_7_i);
    
    \SBYTE_7_r[4]\ : OA21TTF
      port map(A => N_325_i, B => N_324_i, C => N_559, Y => 
        \SBYTE_7[4]\);
    
    \DACCfgValue_9_i_a2[4]\ : NOR2
      port map(A => N_401, B => N_1041, Y => N_402);
    
    \BITCNT_8_r[0]\ : OA21
      port map(A => N_391, B => \DWACT_ADD_CI_0_partial_sum_2[0]\, 
        C => N_562, Y => \BITCNT_8[0]\);
    
    un1_RESCNT_I_64 : XOR2
      port map(A => \RESCNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_64);
    
    F_SO_sync : DFFC
      port map(CLK => CLK_c_c, D => F_SO_sync_2, CLR => 
        HWRES_c_27, Q => \F_SO_sync\);
    
    F_SO_maj : DFFC
      port map(CLK => CLK_c_c, D => F_SO_maj_2, CLR => HWRES_c_26, 
        Q => \F_SO_maj\);
    
    FCS_SEL : DFFS
      port map(CLK => CLK_c_c, D => \FCS_SEL_6\, SET => 
        HWRES_c_26, Q => \FCS_SEL\);
    
    \sstate_ns_1_iv_i_0_a2[2]\ : OR2
      port map(A => N_392, B => N_1047, Y => N_413);
    
    \BYTECNT_9_0_a3[5]\ : AND2
      port map(A => N_437_i_0, B => I_33, Y => \BYTECNT_9[5]\);
    
    un1_RESCNT_G_1 : AND3
      port map(A => \G\, B => G_1_1, C => 
        \DWACT_ADD_CI_0_pog_array_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_3[0]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_31 : XOR2
      port map(A => \REG[474]\, B => \DWACT_ADD_CI_0_TMP_3[0]\, Y
         => \RELOAD_CNT_3[1]\);
    
    \PAGECNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PAGECNT_9[3]\, CLR => 
        HWRES_c_27_0, Q => \PAGECNT_i_0_i[3]\);
    
    \DACCFG_WDT_1[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue[9]_net_1\, CLR
         => HWRES_c_25, Q => DACCFG_WDT(9));
    
    un1_RESCNT_G_2 : AND3FFT
      port map(A => G_2_3_i, B => G_2_2_i, C => \G\, Y => 
        \DWACT_ADD_CI_0_g_array_11_2[0]\);
    
    \sstate_ns_0_0_0[4]\ : OR3
      port map(A => N_361, B => \sstate_ns_0_0_0_0[4]_net_1\, C
         => N_348, Y => \sstate_ns[4]\);
    
    N_400_1_i_i_i_o3 : NAND2FT
      port map(A => PULSE_0, B => PON_LOAD_i, Y => N_1078);
    
    un1_ISCK_1_sqmuxa_i_0_0_1 : NAND3FTT
      port map(A => N_347_i, B => \un1_ISCK_1_sqmuxa_i_0_0_a3\, C
         => N_422, Y => un1_ISCK_1_sqmuxa_i_0_0_1_i);
    
    \SBYTE[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_10\, CLR => HWRES_c_31, 
        Q => \FBOUT[3]\);
    
    un1_RESCNT_I_87 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    \sstate_ns_1_iv_i_5[3]\ : NOR3
      port map(A => N_295_i, B => \sstate_ns_1_iv_i_3_i[3]\, C
         => \sstate_ns_1_iv_i_2_i[3]\, Y => 
        \sstate_ns_1_iv_i_5[3]_net_1\);
    
    un1_FCS_SEL_0_sqmuxa_0_0_a3_0 : NOR3FFT
      port map(A => N_1038_i_0, B => N_1050_i_0, C => N_406, Y
         => N_281_i);
    
    ISI_8_iv_0_i : NOR3FTT
      port map(A => N_1053, B => N_1038, C => N_248, Y => N_115_i);
    
    RELOAD_EDGE : DFFC
      port map(CLK => CLK_c_c, D => NCYC_RELOAD_in, CLR => 
        HWRES_c_29, Q => \RELOAD_EDGE\);
    
    \sstate_ns_1_iv_i_a3_2[3]\ : NOR3FFT
      port map(A => \sstate_0[4]_net_1\, B => \sstate_0[1]_net_1\, 
        C => \sstate_0[3]_net_1\, Y => N_292_i);
    
    un1_RESCNT_I_52 : XOR2
      port map(A => \RESCNT[9]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_3_0[0]\, Y => I_52_1);
    
    SBYTE_14 : MUX2H
      port map(A => \FBOUT[7]\, B => \SBYTE_7[7]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_14\);
    
    \RESCNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \RESCNT_6[1]\, CLR => 
        HWRES_c_30, Q => \RESCNT[1]_net_1\);
    
    \sstate_ns_1_iv_0_0_a3_3_0[0]\ : NOR2FT
      port map(A => N_424, B => \sstate_0[3]_net_1\, Y => 
        \sstate_ns_1_iv_0_0_a3_3_0[0]_net_1\);
    
    \BYTECNT[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[8]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[8]\);
    
    \sstate_ns_1_iv_i_2[3]\ : OAI21FTT
      port map(A => N_1047, B => N_392, C => N_289, Y => 
        \sstate_ns_1_iv_i_2_i[3]\);
    
    \RELOAD_CNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \RELOAD_CNT_3[2]\, CLR => 
        HWRES_c_29, Q => \REG[475]\);
    
    \PAGECNT_9_0_a3[6]\ : AND2
      port map(A => N_436_i_0, B => I_38_2, Y => \PAGECNT_9[6]\);
    
    \DACCfgValue_9_i_a3_0[11]\ : NOR2
      port map(A => \FBOUT[7]\, B => N_402, Y => N_276);
    
    \SBYTE_7_i_i_o2[0]\ : OA21FTF
      port map(A => \sstate[3]_net_1\, B => \sstate[4]_net_1\, C
         => N_1044, Y => N_1046);
    
    \BYTECNT_9_r[3]\ : OA21FTT
      port map(A => N_312, B => I_37, C => un1_pulse_9, Y => 
        \BYTECNT_9[3]\);
    
    un1_RESCNT_I_55 : XOR2
      port map(A => \RESCNT[4]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => I_55);
    
    un1_ISCK_1_sqmuxa_i_0_0_o2_0_0 : NAND2
      port map(A => \PAGECNT_i_0_i[3]\, B => \PAGECNT[4]_net_1\, 
        Y => un1_ISCK_1_sqmuxa_i_0_0_o2_0_i);
    
    \DACCfgValue_9_r[9]\ : NOR3
      port map(A => N_1078_2, B => N_272, C => N_271, Y => 
        \DACCfgValue_9[9]\);
    
    \RESCNT_6_0_a3_7_8[0]\ : NAND3
      port map(A => \RESCNT_6_0_a3_7_6[0]_net_1\, B => 
        \RESCNT[0]_net_1\, C => \RESCNT[1]_net_1\, Y => 
        \RESCNT_6_0_a3_7_8_i[0]\);
    
    \SBYTE_7_i_i_a3_0[4]\ : AND2
      port map(A => \FBOUT[3]\, B => N_1075, Y => N_325_i);
    
    ISI_16 : MUX2H
      port map(A => ISI_net_1, B => ISI_8, S => 
        un1_ISI_1_sqmuxa_1, Y => \ISI_16\);
    
    un1_PAGECNT_1_I_37 : XOR2
      port map(A => \PAGECNT_i_0_i[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_37_0);
    
    un1_NCS0_2_sqmuxa_0_0_a3_0 : OR2
      port map(A => N_418, B => N_1050, Y => N_344);
    
    \RESCNT_6_r[7]\ : OA21
      port map(A => N_313, B => I_61, C => N_528_i_0, Y => 
        \RESCNT_6[7]\);
    
    WRCROMi_0_sqmuxa_1_i_0_a3_0 : OR2
      port map(A => \CROMWAD[3]\, B => \CROMWAD[7]\, Y => 
        \WRCROMi_0_sqmuxa_1_i_0_a3_0\);
    
    un1_BYTECNT_3_I_54 : AND2
      port map(A => \CROMWAD[6]\, B => \CROMWAD[7]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_2_1[0]\);
    
    LUT_5_i_0_o2_1 : NOR3FFT
      port map(A => \CROMWAD[1]\, B => \CROMWAD[2]\, C => 
        \CROMWAD[3]\, Y => N_1062);
    
    \DACCfgValue_9_r[11]\ : NOR3
      port map(A => N_1078_2, B => N_276, C => N_275, Y => 
        \DACCfgValue_9[11]\);
    
    sstate_26_sqmuxa_0_a2_1_a2_0_a3 : NOR2FT
      port map(A => N_432, B => N_1078_0, Y => sstate_26_sqmuxa);
    
    un1_sstate_1_sqmuxa_0_0_0_a3 : NAND2
      port map(A => N_411, B => N_419, Y => N_278);
    
    un1_pulse_7_0_0_0_0 : OAI21
      port map(A => N_1054, B => N_427_1, C => N_434, Y => 
        \un1_pulse_7_0_0_0_0\);
    
    \SBYTE_7_r[3]\ : NOR3
      port map(A => N_559, B => N_327, C => N_326, Y => 
        \SBYTE_7[3]\);
    
    un1_BYTECNT_3_I_30 : XOR2
      port map(A => \CROMWAD[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, Y => I_30_0);
    
    \RESCNT_6_r_i[0]\ : NOR2FT
      port map(A => N_412, B => N_1078_0, Y => N_528_i_0);
    
    un1_pulse_5_0_0_a3 : OR2
      port map(A => \F_SO_sync1\, B => \F_SO_sync2\, Y => N_342);
    
    WRCROMi_0_sqmuxa_1_i_0_a2_1 : NAND3
      port map(A => N_391, B => N_389, C => N_390, Y => N_395);
    
    un1_BYTECNT_3_I_36 : XOR2
      port map(A => \CROMWAD[8]\, B => 
        \DWACT_ADD_CI_0_g_array_3_1[0]\, Y => I_36);
    
    un1_RESCNT_I_102 : AND2
      port map(A => \RESCNT[10]_net_1\, B => \RESCNT[11]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_4[0]\);
    
    un1_PAGECNT_1_I_50 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11_0[0]\, B => 
        \PAGECNT[6]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    WRCROMi_0_sqmuxa_1_i_0 : OR3
      port map(A => N_435, B => N_315, C => un1_pulse_1, Y => 
        N_943);
    
    SBYTE_12 : MUX2H
      port map(A => \FBOUT[5]\, B => \SBYTE_7[5]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_12\);
    
    \DACCfgValue[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACCfgValue_22\, CLR => 
        HWRES_c_26, Q => \DACCfgValue[6]_net_1\);
    
    un1_pulse_9_0_0_o2_0 : OA21TTF
      port map(A => N_408, B => N_413, C => N_398, Y => N_1059);
    
    un1_sstate_1_sqmuxa_0_0_a2_1 : NAND2FT
      port map(A => N_1040, B => \CROMWAD[8]\, Y => N_408);
    
    un1_RESCNT_I_93 : AND2
      port map(A => \RESCNT[6]_net_1\, B => \RESCNT[7]_net_1\, Y
         => \DWACT_ADD_CI_0_pog_array_1_2_0[0]\);
    
    un1_ISI_1_sqmuxa_1_0_a3_0 : OR2
      port map(A => N_351_1, B => N_1044, Y => N_351);
    
    \SBYTE_7_r[6]\ : NOR3
      port map(A => N_559, B => N_331, C => N_330, Y => 
        \SBYTE_7[6]\);
    
    un1_RESCNT_I_58 : XOR2
      port map(A => \RESCNT[12]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_10[0]\, Y => I_58);
    
    SBYTE_10 : MUX2H
      port map(A => \FBOUT[3]\, B => \SBYTE_7[3]\, S => 
        un1_SBYTE_0_sqmuxa, Y => \SBYTE_10\);
    
    P_RELOAD_COUNT_un3_reload_edge : NOR2
      port map(A => \RELOAD_EDGE\, B => RELOAD_EDGE_r_i_0, Y => 
        un3_reload_edge);
    
    un1_RESCNT_I_59 : XOR2
      port map(A => \RESCNT[6]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => I_59);
    
    \sstate_ns_1_iv_0_0_a3_1[0]\ : OR2
      port map(A => N_1063, B => N_1076, Y => 
        \sstate_ns_1_iv_0_0_a3_1[0]_net_1\);
    
    \PDLCFG_WDT_1[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[1]\, CLR => HWRES_c_28, 
        Q => CROMWDT(1));
    
    \sstate_ns_1_iv_0_0[0]\ : OR3
      port map(A => \sstate_ns_1_iv_0_0_3_i[0]\, B => N_373_i, C
         => \sstate_ns_1_iv_0_0_2_i[0]\, Y => \sstate_ns[0]\);
    
    \sstate_ns_1_iv_0_0_a3_0_1[1]\ : NOR2FT
      port map(A => N_1050, B => N_1074, Y => N_353_1);
    
    \RESCNT_6_r[6]\ : OA21
      port map(A => N_313, B => I_59, C => N_528_i_0, Y => 
        \RESCNT_6[6]\);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_39 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_4[0]\);
    
    un1_sstate_17_0_0_0_a2 : OR3FTT
      port map(A => \sstate_0[4]_net_1\, B => N_392, C => 
        \sstate[1]_net_1\, Y => N_425);
    
    un1_BYTECNT_3_I_52 : AND2
      port map(A => \CROMWAD[2]\, B => \CROMWAD[3]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    un1_RESCNT_G_2_3 : NAND3
      port map(A => \DWACT_ADD_CI_0_pog_array_2[0]\, B => G_2_0, 
        C => \RESCNT[0]_net_1\, Y => G_2_3_i);
    
    \DACCfgValue_9_i_a2_0[4]\ : NOR2
      port map(A => N_401, B => N_1041, Y => N_402_0);
    
    \BYTECNT[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \BYTECNT_9[6]\, CLR => 
        HWRES_c_24, Q => \CROMWAD[6]\);
    
    \RESCNT_6_0_a3[0]\ : NOR2
      port map(A => N_313_7_i, B => N_425, Y => N_313);
    
    P_RELOAD_COUNT_RELOAD_CNT_3_I_35 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_3[0]\, B => \REG[474]\, Y
         => \DWACT_ADD_CI_0_g_array_1_3[0]\);
    
    \PDLCFG_WDT_1[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \FBOUT[0]\, CLR => HWRES_c_28, 
        Q => CROMWDT(0));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity event_fifo is

    port( FID       : in    std_logic_vector(31 downto 0);
          DPR       : out   std_logic_vector(31 downto 0);
          WRB       : in    std_logic;
          CLEAR_i_0 : in    std_logic;
          NRDMEB    : in    std_logic;
          CLK_c_c   : in    std_logic;
          FF_c      : out   std_logic;
          EF        : out   std_logic
        );

end event_fifo;

architecture DEF_ARCH of event_fifo is 

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component FIFO256x9SST
    port( DO8    : out   std_logic;
          DO7    : out   std_logic;
          DO6    : out   std_logic;
          DO5    : out   std_logic;
          DO4    : out   std_logic;
          DO3    : out   std_logic;
          DO2    : out   std_logic;
          DO1    : out   std_logic;
          DO0    : out   std_logic;
          FULL   : out   std_logic;
          EMPTY  : out   std_logic;
          EQTH   : out   std_logic;
          GEQTH  : out   std_logic;
          WPE    : out   std_logic;
          RPE    : out   std_logic;
          DOS    : out   std_logic;
          LGDEP2 : in    std_logic := 'U';
          LGDEP1 : in    std_logic := 'U';
          LGDEP0 : in    std_logic := 'U';
          RESET  : in    std_logic := 'U';
          LEVEL7 : in    std_logic := 'U';
          LEVEL6 : in    std_logic := 'U';
          LEVEL5 : in    std_logic := 'U';
          LEVEL4 : in    std_logic := 'U';
          LEVEL3 : in    std_logic := 'U';
          LEVEL2 : in    std_logic := 'U';
          LEVEL1 : in    std_logic := 'U';
          LEVEL0 : in    std_logic := 'U';
          DI8    : in    std_logic := 'U';
          DI7    : in    std_logic := 'U';
          DI6    : in    std_logic := 'U';
          DI5    : in    std_logic := 'U';
          DI4    : in    std_logic := 'U';
          DI3    : in    std_logic := 'U';
          DI2    : in    std_logic := 'U';
          DI1    : in    std_logic := 'U';
          DI0    : in    std_logic := 'U';
          WRB    : in    std_logic := 'U';
          RDB    : in    std_logic := 'U';
          WBLKB  : in    std_logic := 'U';
          RBLKB  : in    std_logic := 'U';
          PARODD : in    std_logic := 'U';
          WCLKS  : in    std_logic := 'U';
          RCLKS  : in    std_logic := 'U';
          DIS    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal net00011, net00012, net00010, net00009, net00008, 
        net00006, net00007, net00005, net00004, net00003, 
        net00068, net00067, net00066, net00065, net00069, 
        net00016, net00021, net00071, net00070, \GND\, \VCC\, 
        net00062, net00015, net00020, net00064, net00063, 
        net00059, net00014, net00019, net00061, net00060, 
        net00056, net00013, net00018, net00058, net00057
         : std_logic;

begin 


    U5 : OR3
      port map(A => net00010, B => net00009, C => net00008, Y => 
        net00012);
    
    U4 : OR2
      port map(A => net00006, B => net00007, Y => FF_c);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    M1 : FIFO256x9SST
      port map(DO8 => DPR(17), DO7 => DPR(16), DO6 => DPR(15), 
        DO5 => DPR(14), DO4 => DPR(13), DO3 => DPR(12), DO2 => 
        DPR(11), DO1 => DPR(10), DO0 => DPR(9), FULL => net00004, 
        EMPTY => net00009, EQTH => net00014, GEQTH => net00019, 
        WPE => net00060, RPE => net00061, DOS => net00059, LGDEP2
         => \VCC\, LGDEP1 => \VCC\, LGDEP0 => \VCC\, RESET => 
        CLEAR_i_0, LEVEL7 => \GND\, LEVEL6 => \GND\, LEVEL5 => 
        \GND\, LEVEL4 => \GND\, LEVEL3 => \GND\, LEVEL2 => \GND\, 
        LEVEL1 => \GND\, LEVEL0 => \VCC\, DI8 => FID(17), DI7 => 
        FID(16), DI6 => FID(15), DI5 => FID(14), DI4 => FID(13), 
        DI3 => FID(12), DI2 => FID(11), DI1 => FID(10), DI0 => 
        FID(9), WRB => WRB, RDB => NRDMEB, WBLKB => \GND\, RBLKB
         => \GND\, PARODD => \GND\, WCLKS => CLK_c_c, RCLKS => 
        CLK_c_c, DIS => \GND\);
    
    M0 : FIFO256x9SST
      port map(DO8 => DPR(8), DO7 => DPR(7), DO6 => DPR(6), DO5
         => DPR(5), DO4 => DPR(4), DO3 => DPR(3), DO2 => DPR(2), 
        DO1 => DPR(1), DO0 => DPR(0), FULL => net00003, EMPTY => 
        net00008, EQTH => net00013, GEQTH => net00018, WPE => 
        net00057, RPE => net00058, DOS => net00056, LGDEP2 => 
        \VCC\, LGDEP1 => \VCC\, LGDEP0 => \VCC\, RESET => 
        CLEAR_i_0, LEVEL7 => \GND\, LEVEL6 => \GND\, LEVEL5 => 
        \GND\, LEVEL4 => \GND\, LEVEL3 => \GND\, LEVEL2 => \GND\, 
        LEVEL1 => \GND\, LEVEL0 => \VCC\, DI8 => FID(8), DI7 => 
        FID(7), DI6 => FID(6), DI5 => FID(5), DI4 => FID(4), DI3
         => FID(3), DI2 => FID(2), DI1 => FID(1), DI0 => FID(0), 
        WRB => WRB, RDB => NRDMEB, WBLKB => \GND\, RBLKB => \GND\, 
        PARODD => \GND\, WCLKS => CLK_c_c, RCLKS => CLK_c_c, DIS
         => \GND\);
    
    U3 : OR3
      port map(A => net00005, B => net00004, C => net00003, Y => 
        net00007);
    
    M2 : FIFO256x9SST
      port map(DO8 => DPR(26), DO7 => DPR(25), DO6 => DPR(24), 
        DO5 => DPR(23), DO4 => DPR(22), DO3 => DPR(21), DO2 => 
        DPR(20), DO1 => DPR(19), DO0 => DPR(18), FULL => net00005, 
        EMPTY => net00010, EQTH => net00015, GEQTH => net00020, 
        WPE => net00063, RPE => net00064, DOS => net00062, LGDEP2
         => \VCC\, LGDEP1 => \VCC\, LGDEP0 => \VCC\, RESET => 
        CLEAR_i_0, LEVEL7 => \GND\, LEVEL6 => \GND\, LEVEL5 => 
        \GND\, LEVEL4 => \GND\, LEVEL3 => \GND\, LEVEL2 => \GND\, 
        LEVEL1 => \GND\, LEVEL0 => \VCC\, DI8 => FID(26), DI7 => 
        FID(25), DI6 => FID(24), DI5 => FID(23), DI4 => FID(22), 
        DI3 => FID(21), DI2 => FID(20), DI1 => FID(19), DI0 => 
        FID(18), WRB => WRB, RDB => NRDMEB, WBLKB => \GND\, RBLKB
         => \GND\, PARODD => \GND\, WCLKS => CLK_c_c, RCLKS => 
        CLK_c_c, DIS => \GND\);
    
    U6 : OR2
      port map(A => net00011, B => net00012, Y => EF);
    
    M3 : FIFO256x9SST
      port map(DO8 => net00065, DO7 => net00066, DO6 => net00067, 
        DO5 => net00068, DO4 => DPR(31), DO3 => DPR(30), DO2 => 
        DPR(29), DO1 => DPR(28), DO0 => DPR(27), FULL => net00006, 
        EMPTY => net00011, EQTH => net00016, GEQTH => net00021, 
        WPE => net00070, RPE => net00071, DOS => net00069, LGDEP2
         => \VCC\, LGDEP1 => \VCC\, LGDEP0 => \VCC\, RESET => 
        CLEAR_i_0, LEVEL7 => \GND\, LEVEL6 => \GND\, LEVEL5 => 
        \GND\, LEVEL4 => \GND\, LEVEL3 => \GND\, LEVEL2 => \GND\, 
        LEVEL1 => \GND\, LEVEL0 => \VCC\, DI8 => \GND\, DI7 => 
        \GND\, DI6 => \GND\, DI5 => \GND\, DI4 => FID(31), DI3
         => FID(30), DI2 => FID(29), DI1 => FID(28), DI0 => 
        FID(27), WRB => WRB, RDB => NRDMEB, WBLKB => \GND\, RBLKB
         => \GND\, PARODD => \GND\, WCLKS => CLK_c_c, RCLKS => 
        CLK_c_c, DIS => \GND\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity ROC32 is

    port( DPR          : out   std_logic_vector(31 downto 0);
          un2_evread_0 : out   std_logic;
          CHANNEL      : out   std_logic_vector(2 downto 0);
          CHIP_ADDR    : out   std_logic_vector(2 downto 0);
          I2C_RDATA    : in    std_logic_vector(9 downto 0);
          OR_RDATA     : in    std_logic_vector(9 downto 0);
          PDL_RDATA    : in    std_logic_vector(7 downto 0);
          GA_c         : in    std_logic_vector(3 downto 0);
          OR_RADDR     : out   std_logic_vector(5 downto 0);
          PDL_RADDR    : out   std_logic_vector(5 downto 0);
          LBSP_c       : in    std_logic_vector(2 to 2);
          LBSP_c_1     : in    std_logic_vector(2 to 2);
          LBSP_c_0     : in    std_logic_vector(2 to 2);
          PULSE        : in    std_logic_vector(3 downto 2);
          REG_i_0      : in    std_logic_vector(5 to 5);
          REG_c        : in    std_logic_vector(23 downto 21);
          REG_330      : out   std_logic;
          REG_329      : out   std_logic;
          REG_328      : out   std_logic;
          REG_408      : in    std_logic;
          REG_410      : in    std_logic;
          REG_432      : in    std_logic;
          REG_415      : in    std_logic;
          REG_406      : in    std_logic;
          REG_418      : in    std_logic;
          REG_421      : in    std_logic;
          REG_430      : in    std_logic;
          REG_433      : in    std_logic;
          REG_424      : in    std_logic;
          REG_427      : in    std_logic;
          REG_416      : in    std_logic;
          REG_419      : in    std_logic;
          REG_412      : in    std_logic;
          REG_413      : in    std_logic;
          REG_428      : in    std_logic;
          REG_431      : in    std_logic;
          REG_422      : in    std_logic;
          REG_425      : in    std_logic;
          REG_414      : in    std_logic;
          REG_417      : in    std_logic;
          REG_409      : in    std_logic;
          REG_411      : in    std_logic;
          REG_426      : in    std_logic;
          REG_429      : in    std_logic;
          REG_420      : in    std_logic;
          REG_423      : in    std_logic;
          REG_407      : in    std_logic;
          REG_434      : in    std_logic;
          REG_435      : in    std_logic;
          REG_404      : in    std_logic;
          REG_405      : in    std_logic;
          REG_43       : in    std_logic;
          REG_44       : in    std_logic;
          REG_45       : in    std_logic;
          REG_46       : in    std_logic;
          REG_47       : in    std_logic;
          REG_48       : in    std_logic;
          REG_49       : in    std_logic;
          REG_50       : in    std_logic;
          REG_51       : in    std_logic;
          REG_52       : in    std_logic;
          REG_53       : in    std_logic;
          REG_54       : in    std_logic;
          REG_55       : in    std_logic;
          REG_56       : in    std_logic;
          REG_57       : in    std_logic;
          REG_58       : in    std_logic;
          REG_59       : in    std_logic;
          REG_60       : in    std_logic;
          REG_61       : in    std_logic;
          REG_62       : in    std_logic;
          REG_63       : in    std_logic;
          REG_64       : in    std_logic;
          REG_65       : in    std_logic;
          REG_66       : in    std_logic;
          REG_67       : in    std_logic;
          REG_68       : in    std_logic;
          REG_69       : in    std_logic;
          REG_70       : in    std_logic;
          REG_71       : in    std_logic;
          REG_72       : in    std_logic;
          REG_73       : in    std_logic;
          REG_74       : in    std_logic;
          REG_41       : out   std_logic;
          REG_42       : out   std_logic;
          REG_0        : in    std_logic;
          REG_15       : out   std_logic;
          REG_27       : out   std_logic;
          REG_28       : out   std_logic;
          REG_30       : out   std_logic;
          REG_29       : out   std_logic;
          REG_39       : out   std_logic;
          REG_37       : out   std_logic;
          REG_36       : out   std_logic;
          REG_34       : out   std_logic;
          REG_33       : out   std_logic;
          REG_38       : out   std_logic;
          REG_35       : out   std_logic;
          REG_40       : out   std_logic;
          REG_31       : out   std_logic;
          REG_32       : out   std_logic;
          EF           : out   std_logic;
          FF_c         : out   std_logic;
          NRDMEB       : in    std_logic;
          CLEAR_i_0    : in    std_logic;
          CLEAR_14     : in    std_logic;
          CLEAR_13     : in    std_logic;
          CLEAR_4      : in    std_logic;
          CLEAR_3      : in    std_logic;
          CLEAR_2      : in    std_logic;
          CLEAR_8      : in    std_logic;
          CLEAR_7      : in    std_logic;
          CLEAR_6      : in    std_logic;
          CLEAR_11     : in    std_logic;
          CLEAR_10     : in    std_logic;
          CLEAR_19     : in    std_logic;
          CLEAR_9      : in    std_logic;
          CLEAR_18     : in    std_logic;
          CLEAR_12     : in    std_logic;
          CLEAR_15     : in    std_logic;
          CLEAR_20     : in    std_logic;
          CLEAR_5      : in    std_logic;
          PDL_RACK     : in    std_logic;
          CLEAR_17     : in    std_logic;
          OR_RACK      : in    std_logic;
          CLEAR_16     : in    std_logic;
          L2R_c_c      : in    std_logic;
          L2A_c_c      : in    std_logic;
          HWRES_c_12   : in    std_logic;
          L1A_c_c      : in    std_logic;
          ALICLK_c     : in    std_logic;
          HWRES_c_11   : in    std_logic;
          DTEST_FIFO   : out   std_logic;
          I2C_CHAIN    : out   std_logic;
          PDL_RREQ     : out   std_logic;
          I2C_RREQ     : out   std_logic;
          EVRDY_c      : out   std_logic;
          OR_RREQ      : out   std_logic;
          I2C_RACK     : in    std_logic;
          EVNT_TRG     : out   std_logic;
          EVREAD       : in    std_logic;
          CLK_c_c      : in    std_logic;
          CLEAR_0      : in    std_logic;
          I_8          : in    std_logic;
          I_16         : in    std_logic
        );

end ROC32;

architecture DEF_ARCH of ROC32 is 

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component AND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NAND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component event_fifo
    port( FID       : in    std_logic_vector(31 downto 0) := (others => 'U');
          DPR       : out   std_logic_vector(31 downto 0);
          WRB       : in    std_logic := 'U';
          CLEAR_i_0 : in    std_logic := 'U';
          NRDMEB    : in    std_logic := 'U';
          CLK_c_c   : in    std_logic := 'U';
          FF_c      : out   std_logic;
          EF        : out   std_logic
        );
  end component;

  component MUX2L
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \DWACT_ADD_CI_0_TMP[0]\, \CNT[0]_net_1\, 
        \un1_EVENT_DWORD_0_sqmuxa_0_0\, I_26, \CNT[5]_net_1\, 
        I_30, N_176, \STATE1_0[2]_net_1\, \STATE1_0[1]_net_1\, 
        N_1762, N_195, N_234, N_1593, N_215, N_1454_0, N_520, 
        ADD_16x16_slow_I5_CO1_0_a0_0, \CNT_8_i[5]_net_1\, N_185_i, 
        \DWACT_ADD_CI_0_g_array_2[0]\, \CNT[4]_net_1\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, \CNT_0[1]_net_1\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, \OR_RACK_sync\, G_0_x2, 
        ADD_16x16_slow_I14_S_0, G_0_o2, I12_un1_CO1, 
        ADD_16x16_slow_I13_CO1_0, I8_un4_CO1, N220, I11_un3_CO1, 
        I10_un1_CO1, I6_un4_CO1, G_8_0_a2_2, G_8_0_x2, N_19, 
        \FIFO_END_EVNT\, G_6, N_7210_i, I6_un1_CO1_i_0_i, N_55, 
        N_54, I7_un3_CO1, ADD_16x16_slow_I7_CO1_0, I8_un1_CO1, 
        ADD_16x16_slow_I8_un1_CO1_0, N224, 
        ADD_16x16_slow_I9_CO1_0, G_11_0_a2_0, \REG[42]\, N228, 
        ADD_16x16_slow_I11_CO1_0_m5_0, 
        ADD_16x16_slow_I12_un1_CO1_0, un5_evread_7, G_6_0, 
        ADD_16x16_slow_I3_CO1_1_0_i_i, 
        ADD_16x16_slow_I6_un1_CO1_0, N_43, 
        ADD_16x16_slow_I2_un1_CO1_0_a0_0, 
        ADD_16x16_slow_I6_un1_CO1_0_a0_2, 
        ADD_16x16_slow_I5_CO1_0_a0_3, 
        ADD_16x16_slow_I6_un4_CO1_5_tz, N_176_0, N_1585_0, 
        \STATE1[0]_net_1\, \STATE1[3]_net_1\, \CNT_0[0]_net_1\, 
        \CNT_8_i[0]_net_1\, \CNT_8_i[1]_net_1\, \CNT_0[2]_net_1\, 
        N_78, \CNT_0[3]_net_1\, N_81, \CNT_0[4]_net_1\, N_84, 
        \CNT_0[5]_net_1\, \STATE1_0[0]_net_1\, \STATE1_ns[0]\, 
        \STATE1_ns_i_0[1]_net_1\, \STATE1_ns[2]\, 
        \STATE1_0[3]_net_1\, \STATE1_ns[3]\, N_205_1, N_1587, 
        N_522, N_253, N_205_0, N_532_3_8, N_532_3_7, N_532_3_6, 
        N_532_3_5, N_532_3_4, N_532_3_3, N_532_3_2, N_532_3_1, 
        N_1585, N_532_3_0, N_1574_1, N_1574_0, N_620_4_1, N_1573, 
        N_221, N_620_4_0, N_1575_1, N_1575_0, \un2_evread_1[14]\, 
        \un2_evread_0[14]\, N_105_i_0_1, N_105_i_0_0, 
        un4_bnc_res_i_1, un4_bnc_res_NE_29_i, un4_bnc_res_NE_25_i, 
        un4_bnc_res_NE_24_i, un4_bnc_res_i_0, un1_STATE1_18_1, 
        N_1673_i, N_1672, un1_STATE1_18_0, N_1469_1, N_1469_0, 
        N_1229_i_1, N_180, N_1755_i, N_1229_i_0, N_190_i_0, 
        N_1768_i, N_701_i_0_0, N_193, N_252, 
        \DWACT_ADD_CI_0_g_array_3[0]\, 
        \DWACT_ADD_CI_0_g_array_2_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_2[0]\, 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\, 
        \DWACT_ADD_CI_0_g_array_11_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_3[0]\, 
        \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_TMP_0[0]\, \EVNT_NUM[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, \EVNT_NUM[4]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, \EVNT_NUM[6]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, \EVNT_NUM[8]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_4[0]\, \EVNT_NUM[10]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12[0]\, \EVNT_NUM[2]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, N_157, 
        \BNC_CNT[1]_net_1\, \BNC_CNT[0]_net_1\, N_149, 
        \BNC_CNT[3]_net_1\, \DWACT_FINC_E[0]\, N_126, 
        \BNC_CNT[8]_net_1\, \DWACT_FINC_E[4]\, N_111, 
        \DWACT_FINC_E[7]\, \DWACT_FINC_E[6]\, 
        \FAULT_STROBE_0_2_i\, \CLEAR_PSM_FLAGS\, N_701_i_0, 
        \REG_1_20_127_i_a2\, N_226_i_0, I_24_2, I_23, I_22_0, 
        I_21_0, \DWACT_ADD_CI_0_partial_sum[0]\, N_183, N_192, 
        N_1600, N_1759_i, N_1758_1, N_199, N_1757, N_120_i, N_188, 
        \STATE2_ns_i_i_a2_i[1]_net_1\, \STATE2[2]_net_1\, 
        \TRIGGER_sync\, N_161_i_0, N_1569_i, 
        \STATE1_ns_i_0_5_i[1]\, N_7189_i, 
        \STATE1_ns_i_0_4[1]_net_1\, \STATE1_ns_i_0_2[1]_net_1\, 
        N_1564, N_242, \STATE1_ns_i_0_1[1]_net_1\, N_1562_i, 
        N_1568_i, N_1563_i, \READ_PDL_FLAG\, \READ_ADC_FLAG\, 
        N_1576_1, N_1470, N_166, N_289, N_1195_1, 
        \RDY_CNT_8_i_0[1]_net_1\, N_267, I_10, 
        \RDY_CNT_8_i_0[0]_net_1\, 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, N_1583, N_1582, N_222, 
        \PDL_RACK_sync\, N_243, N_1733_i, 
        \STATE1_ns_0_0_0_2_i[3]\, STATE1_1_sqmuxa_1, 
        \STATE1_ns_0_0_0_0_i[3]\, N_1734, 
        \STATE1_ns_0_0_0_i_0[3]_net_1\, N_207, N_1731, N_230, 
        N_1601, N_1771, \STATE1_d[7]\, N_1733_1, N_620_4, 
        \STATE2_ns[0]\, \STATE2[1]_net_1\, \STATE2_ns[2]\, 
        \READ_OR_FLAG_91_i_0\, N_1539, N_1540, N_258_i_0, 
        \STATE1[1]_net_1\, \READ_OR_FLAG\, \STATE1_d[9]\, N_1777, 
        \STATE1[2]_net_1\, \STATE1_ns_1_iv_0_0_7[2]_net_1\, 
        N_1559_i, \STATE1_ns_1_iv_0_0_5_i[2]\, 
        \STATE1_ns_1_iv_0_0_2_i[2]\, 
        \STATE1_ns_1_iv_0_0_3[2]_net_1\, N_1586, N_1558_i, 
        N_215_i_0, \STATE1_ns_1_iv_0_0_a2_4_1[2]_net_1\, 
        \STATE1_ns_1_iv_0_0_1[2]_net_1\, EVNT_TRG_net_1, 
        \STATE1_ns_1_iv_0_0_0[2]_net_1\, 
        \STATE1_ns_1_iv_0_0_a2_3_1[2]_net_1\, N_1557, 
        \STATE1_i_0[2]\, \STATE1_i_0[3]\, 
        \STATE1_ns_1_iv_0_0_a2_0[0]_net_1\, N_1614, N_1778, 
        N_1752_1, \STATE1_ns_1_iv_0_0_o3_4[0]_net_1\, 
        \STATE1_ns_1_iv_0_0_o3_2_i[0]\, 
        \STATE1_ns_1_iv_0_0_o3_1_i[0]\, N_1575, N_1613, N_7200_i, 
        N_1470_i_0, \L2ASS\, \STATE1_ns_1_iv_0_0_a3_0_1[0]_net_1\, 
        \STATE1_ns_1_iv_0_0_o3_0[0]_net_1\, \RDY_CNT[0]_net_1\, 
        \RDY_CNT[1]_net_1\, N_1750, N_1183_i, N_1744, N_1746, 
        \STATE1_ns_1_iv_0_1_o2_3_o3_0[0]_net_1\, N_237, 
        \BNC_CNT_247\, \BNC_CNT[31]_net_1\, \BNC_CNT_3[31]_net_1\, 
        I_224, \BNC_CNT_246\, \BNC_CNT[30]_net_1\, 
        \BNC_CNT_3[30]_net_1\, I_217, \BNC_CNT_245\, 
        \BNC_CNT[29]_net_1\, \BNC_CNT_3[29]_net_1\, I_210, 
        \BNC_CNT_244\, \BNC_CNT[28]_net_1\, \BNC_CNT_3[28]_net_1\, 
        I_203, \BNC_CNT_243\, \BNC_CNT[27]_net_1\, 
        \BNC_CNT_3[27]_net_1\, I_196, \BNC_CNT_242\, 
        \BNC_CNT[26]_net_1\, \BNC_CNT_3[26]_net_1\, I_186, 
        \BNC_CNT_241\, \BNC_CNT[25]_net_1\, \BNC_CNT_3[25]_net_1\, 
        I_173, \BNC_CNT_240\, \BNC_CNT[24]_net_1\, 
        \BNC_CNT_3[24]_net_1\, I_166, \BNC_CNT_239\, 
        \BNC_CNT[23]_net_1\, \BNC_CNT_3[23]_net_1\, I_156, 
        \BNC_CNT_238\, \BNC_CNT[22]_net_1\, \BNC_CNT_3[22]_net_1\, 
        I_143, \BNC_CNT_237\, \BNC_CNT[21]_net_1\, 
        \BNC_CNT_3[21]_net_1\, I_136, \BNC_CNT_236\, 
        \BNC_CNT[20]_net_1\, \BNC_CNT_3[20]_net_1\, I_129, 
        \BNC_CNT_235\, \BNC_CNT[19]_net_1\, \BNC_CNT_3[19]_net_1\, 
        I_122, \BNC_CNT_234\, \BNC_CNT[18]_net_1\, 
        \BNC_CNT_3[18]_net_1\, I_115, \BNC_CNT_233\, 
        \BNC_CNT[17]_net_1\, \BNC_CNT_3[17]_net_1\, I_105, 
        \BNC_CNT_232\, \BNC_CNT[16]_net_1\, \BNC_CNT_3[16]_net_1\, 
        I_98, \BNC_CNT_231\, \BNC_CNT[15]_net_1\, 
        \BNC_CNT_3[15]_net_1\, I_91_0, \BNC_CNT_230\, 
        \BNC_CNT[14]_net_1\, \BNC_CNT_3[14]_net_1\, I_84_0, 
        \BNC_CNT_229\, \BNC_CNT[13]_net_1\, \BNC_CNT_3[13]_net_1\, 
        I_77_0, \BNC_CNT_228\, \BNC_CNT[12]_net_1\, 
        \BNC_CNT_3[12]_net_1\, I_73_0, \BNC_CNT_227\, 
        \BNC_CNT[11]_net_1\, \BNC_CNT_3[11]_net_1\, I_66_0, 
        \BNC_CNT_226\, \BNC_CNT[10]_net_1\, \BNC_CNT_3[10]_net_1\, 
        I_56_0, un4_bnc_res_i, \BNC_CNT_225\, \BNC_CNT[9]_net_1\, 
        \BNC_CNT_3[9]_net_1\, I_52_0, \BNC_CNT_224\, 
        \BNC_CNT_3[8]_net_1\, I_45_0, \BNC_CNT_223\, 
        \BNC_CNT[7]_net_1\, \BNC_CNT_3[7]_net_1\, I_38_0, 
        \BNC_CNT_222\, \BNC_CNT[6]_net_1\, \BNC_CNT_3[6]_net_1\, 
        I_31_0, \BNC_CNT_221\, \BNC_CNT[5]_net_1\, 
        \BNC_CNT_3[5]_net_1\, I_24_1, \BNC_CNT_220\, 
        \BNC_CNT[4]_net_1\, \BNC_CNT_3[4]_net_1\, I_20_1, 
        \BNC_CNT_219\, \BNC_CNT_3[3]_net_1\, I_13_3, 
        \BNC_CNT_218\, \BNC_CNT[2]_net_1\, \BNC_CNT_3[2]_net_1\, 
        I_9_2, \BNC_CNT_217\, \BNC_CNT_3[1]_net_1\, I_5_2, 
        \BNC_CNT_216\, \BNC_CNT_3[0]_net_1\, \PDL_RADDR_215\, 
        \PDL_RADDR_214\, \PDL_RADDR_213\, \CNT[3]_net_1\, 
        \PDL_RADDR_212\, \CNT[2]_net_1\, \PDL_RADDR_211\, 
        \CNT[1]_net_1\, \PDL_RADDR_210\, \OR_RADDR_209\, N_679, 
        N_248, \OR_RADDR_208\, N_681, \OR_RADDR_207\, N_683, 
        \OR_RADDR_206\, N_685, \OR_RADDR_205\, N_687, 
        \OR_RADDR_204\, N_689, \OR_RREQ_203\, N_252_i_0, N_203, 
        N_1454, \un1_STATE1_24_i_i_a2_1\, N_1205_i_i_o2_2_i, 
        \ORATETMO_i_i[3]\, \ORATETMO[4]_net_1\, \ORATETMO_i_i[0]\, 
        \ORATETMO_i_i[1]\, \ORATETMO[2]_net_1\, \EVRDYi_202\, 
        EVREAD_i_0, \un1_reg154\, un5_evread_i_0, 
        \un2_evread[15]_net_1\, un5_evread_11_i, un5_evread_8_i, 
        un5_evread_7_0_i, \un5_evread_4\, \REG[45]\, \REG[38]\, 
        \REG[41]\, \un5_evread_5\, \REG[43]\, \REG[44]\, 
        \REG[39]\, \un5_evread_1\, un5_evread_6_i, \REG[37]\, 
        \REG[40]\, \REG[36]\, \FID_201\, \FID[31]_net_1\, 
        \FID_6[31]\, N_1497_i, N_1498_i, \EVENT_DWORD[31]_net_1\, 
        N_1574, \FID_200\, \FID[30]_net_1\, \FID_6[30]\, N_1515, 
        N_1516, \EVENT_DWORD[30]_net_1\, \FID_199\, 
        \FID[29]_net_1\, \FID_6[29]\, N_1545_i, N_1546_i, 
        \EVENT_DWORD[29]_net_1\, \FID_198\, \FID[28]_net_1\, 
        \FID_6[28]\, N_1536_i, \FID_6_iv_0_0_0_i[28]\, 
        \EVENT_DWORD[28]_net_1\, \FID_197\, \FID[27]_net_1\, 
        \FID_6[27]\, N_1544_i, \FID_6_iv_0_0_i[27]\, 
        \EVNT_NUM[11]_net_1\, N_1543, \EVENT_DWORD[27]_net_1\, 
        \FID_196\, \FID[26]_net_1\, \FID_6[26]\, N_1496_i, 
        \FID_6_iv_0_0_0_i[26]\, N_1495, \EVENT_DWORD[26]_net_1\, 
        \FID_195\, \FID[25]_net_1\, \FID_6[25]\, N_1493_i, 
        \FID_6_iv_0_0_0_i[25]\, \EVNT_NUM[9]_net_1\, N_1492, 
        \EVENT_DWORD[25]_net_1\, \FID_194\, \FID[24]_net_1\, 
        \FID_6[24]\, N_1490_i, \FID_6_iv_0_0_0_i[24]\, N_1489, 
        \EVENT_DWORD[24]_net_1\, \FID_193\, \FID[23]_net_1\, 
        \FID_6[23]\, N_1487_i, \FID_6_iv_0_0_0_i[23]\, 
        \EVNT_NUM[7]_net_1\, N_1486, \EVENT_DWORD[23]_net_1\, 
        \FID_192\, \FID[22]_net_1\, \FID_6[22]\, N_1514_i, 
        \FID_6_iv_0_0_0_i[22]\, N_1513, \EVENT_DWORD[22]_net_1\, 
        \FID_191\, \FID[21]_net_1\, \FID_6[21]\, N_1484_i, 
        \FID_6_iv_0_0_0_i[21]\, \EVNT_NUM[5]_net_1\, N_1483, 
        \EVENT_DWORD[21]_net_1\, \FID_190\, \FID[20]_net_1\, 
        \FID_6[20]\, N_1481_i, \FID_6_iv_0_0_0_i[20]\, N_1480, 
        \EVENT_DWORD[20]_net_1\, \FID_189\, \FID[19]_net_1\, 
        \FID_6[19]\, N_324_i, \FID_6_iv_0_0_i[19]\, 
        \EVNT_NUM[3]_net_1\, N_323, \EVENT_DWORD[19]_net_1\, 
        \FID_188\, \FID[18]_net_1\, \FID_6[18]\, N_1550_i, 
        \FID_6_iv_0_0_1_i[18]\, \FID_6_iv_0_0_0[18]_net_1\, 
        \FAULT_STAT\, N_1547, \EVENT_DWORD[18]_net_1\, \FID_187\, 
        \FID[17]_net_1\, \FID_6[17]\, N_1555_i, 
        \FID_6_iv_0_0_1_i[17]\, \FID_6_iv_0_0_0[17]_net_1\, 
        \CYC_STAT\, N_1552, \EVENT_DWORD[17]_net_1\, \FID_186\, 
        \FID[16]_net_1\, \FID_6[16]\, N_1534_i, 
        \FID_6_iv_0_0_0_i[16]\, \EVNT_NUM[0]_net_1\, N_1533, 
        \EVENT_DWORD[16]_net_1\, \FID_185\, \FID[15]_net_1\, 
        \FID_6[15]\, N_1478_i, \FID_6_iv_0_0_0_i[15]\, N_57_i_0_i, 
        N_1477, \CRC32[11]_net_1\, \CRC32[23]_net_1\, 
        \EVENT_DWORD[15]_net_1\, \FID_184\, \FID[14]_net_1\, 
        \FID_6[14]\, N_1511_i, \FID_6_iv_0_0_0_i[14]\, 
        N_270_i_0_i, N_1510, \CRC32[10]_net_1\, \CRC32[22]_net_1\, 
        \EVENT_DWORD[14]_net_1\, \FID_183\, \FID[13]_net_1\, 
        \FID_6[13]\, N_1531_i, \FID_6_iv_0_0_0_i[13]\, 
        N_269_i_0_i, N_1530, \CRC32[9]_net_1\, \CRC32[21]_net_1\, 
        \EVENT_DWORD[13]_net_1\, \FID_182\, \FID[12]_net_1\, 
        \FID_6[12]\, N_1508_i, \FID_6_iv_0_0_0_i[12]\, 
        N_271_i_0_i, N_1507, \CRC32[8]_net_1\, \CRC32[20]_net_1\, 
        \EVENT_DWORD[12]_net_1\, \FID_181\, \FID[11]_net_1\, 
        \FID_6[11]\, N_1475_i, \FID_6_iv_0_0_0_i[11]\, 
        \FID_2_i[11]\, N_1474, \CRC32[7]_net_1\, 
        \FID_2_0[11]_net_1\, \CRC32[19]_net_1\, \CRC32[31]_net_1\, 
        \EVENT_DWORD[11]_net_1\, \FID_180\, \FID[10]_net_1\, 
        \FID_6[10]\, N_1472_i, \FID_6_iv_0_0_0_i[10]\, 
        \FID_2_i[10]\, N_1471, \CRC32[6]_net_1\, 
        \FID_2_0[10]_net_1\, \CRC32[18]_net_1\, \CRC32[30]_net_1\, 
        \EVENT_DWORD[10]_net_1\, \FID_179\, \FID[9]_net_1\, 
        \FID_6[9]\, N_205, N_1528, \FID_6_iv_0_0_0[9]_net_1\, 
        N_1526, \FID_2[9]_net_1\, \CRC32[5]_net_1\, 
        \FID_2_0[9]_net_1\, \CRC32[17]_net_1\, \CRC32[29]_net_1\, 
        \EVENT_DWORD[9]_net_1\, \FID_178\, \FID[8]_net_1\, 
        \FID_6[8]\, N_1525, \FID_6_iv_0_0_0[8]_net_1\, N_1523, 
        \FID_2[8]_net_1\, \CRC32[4]_net_1\, \FID_2_0[8]_net_1\, 
        \CRC32[16]_net_1\, \CRC32[28]_net_1\, 
        \EVENT_DWORD[8]_net_1\, \FID_177\, \FID[7]_net_1\, 
        \FID_6[7]\, N_320_i, \FID_6_iv_0_0_0_i[7]\, \FID_2_i[7]\, 
        N_319, \CRC32[3]_net_1\, \FID_2_0[7]_net_1\, 
        \CRC32[15]_net_1\, \CRC32[27]_net_1\, 
        \EVENT_DWORD[7]_net_1\, \FID_176\, \FID[6]_net_1\, 
        \FID_6[6]\, N_317_i, \FID_6_iv_0_0_0_i[6]\, \FID_2_i[6]\, 
        N_316, \CRC32[2]_net_1\, \FID_2_0[6]_net_1\, 
        \CRC32[14]_net_1\, \CRC32[26]_net_1\, 
        \EVENT_DWORD[6]_net_1\, \FID_175\, \FID[5]_net_1\, 
        \FID_6[5]\, N_1522, \FID_6_iv_0_0_0[5]_net_1\, N_1520, 
        \FID_2[5]_net_1\, \CRC32[1]_net_1\, \FID_2_0[5]_net_1\, 
        \CRC32[13]_net_1\, \CRC32[25]_net_1\, 
        \EVENT_DWORD[5]_net_1\, \FID_174\, \FID[4]_net_1\, 
        \FID_6[4]\, N_343_i, \FID_6_iv_0_0_0_i[4]\, \FID_2_i[4]\, 
        N_342, \CRC32[0]_net_1\, \FID_2_0[4]_net_1\, 
        \CRC32[12]_net_1\, \CRC32[24]_net_1\, 
        \EVENT_DWORD[4]_net_1\, \FID_173\, \FID[3]_net_1\, 
        \FID_6[3]\, N_309_i, \FID_6_0_iv_0_0_0_i[3]\, N_311, 
        \EVENT_DWORD[3]_net_1\, N_235, \FID_172\, \FID[2]_net_1\, 
        \FID_6[2]\, N_1517_i, \FID_6_0_iv_0_0_0_i[2]\, N_1519, 
        \EVENT_DWORD[2]_net_1\, \FID_171\, \FID[1]_net_1\, 
        \FID_6[1]\, N_1503_i, \FID_6_0_iv_0_0_0_i[1]\, N_1505, 
        \EVENT_DWORD[1]_net_1\, \FID_170\, \FID[0]_net_1\, 
        \FID_6[0]\, N_1500_i, \FID_6_0_iv_0_0_0_i[0]\, N_1502, 
        \EVENT_DWORD[0]_net_1\, \EVENT_DWORD_169\, 
        \EVENT_DWORD_17[31]\, N_1590, \EVENT_DWORD_168\, 
        \EVENT_DWORD_17[30]\, \EVENT_DWORD_167\, 
        \EVENT_DWORD_17[29]\, N_1683, 
        \EVENT_DWORD_17_i_1[29]_net_1\, 
        \EVENT_DWORD_17_i_0[29]_net_1\, N_1682, \EVENT_DWORD_166\, 
        \EVENT_DWORD_17[28]\, N_1694, 
        \EVENT_DWORD_17_i_0_1[28]_net_1\, 
        \EVENT_DWORD_17_i_0_0[28]_net_1\, N_1695, 
        \EVENT_DWORD_165\, \EVENT_DWORD_17[27]\, N_1679, 
        \EVENT_DWORD_17_i_1[27]_net_1\, 
        \EVENT_DWORD_17_i_0[27]_net_1\, N_1678, \EVENT_DWORD_164\, 
        \EVENT_DWORD_17[26]\, N_1698, 
        \EVENT_DWORD_17_i_0_1[26]_net_1\, 
        \EVENT_DWORD_17_i_0_0[26]_net_1\, N_1699, 
        \EVENT_DWORD_163\, \EVENT_DWORD_17[25]\, N_1737, 
        \EVENT_DWORD_17_i_0_1[25]_net_1\, 
        \EVENT_DWORD_17_i_0_0[25]_net_1\, N_1736, 
        \EVENT_DWORD_162\, \EVENT_DWORD_17[24]\, N_1706, 
        \EVENT_DWORD_17_i_0_1[24]_net_1\, 
        \EVENT_DWORD_17_i_0_0[24]_net_1\, N_1707, 
        \EVENT_DWORD_161\, \EVENT_DWORD_17[23]\, N_1714, 
        \EVENT_DWORD_17_i_0_1[23]_net_1\, 
        \EVENT_DWORD_17_i_0_0[23]_net_1\, N_1715, 
        \EVENT_DWORD_160\, \EVENT_DWORD_17[22]\, N_1710, 
        \EVENT_DWORD_17_i_0_1[22]_net_1\, 
        \EVENT_DWORD_17_i_0_0[22]_net_1\, N_1711, 
        \EVENT_DWORD_159\, \EVENT_DWORD_17[21]\, N_1718, 
        \EVENT_DWORD_17_i_0_1[21]_net_1\, 
        \EVENT_DWORD_17_i_0_0[21]_net_1\, N_1719, 
        \EVENT_DWORD_158\, \EVENT_DWORD_17[20]\, N_1702, 
        \EVENT_DWORD_17_i_0_1[20]_net_1\, 
        \EVENT_DWORD_17_i_0_0[20]_net_1\, N_1703, 
        \EVENT_DWORD_157\, \EVENT_DWORD_17[19]\, N_1676, 
        \EVENT_DWORD_17_i_0[19]_net_1\, N_1675, \EVENT_DWORD_156\, 
        \EVENT_DWORD_17[18]\, N_1666, 
        \EVENT_DWORD_17_i_0_0[18]_net_1\, N_1667, 
        \EVENT_DWORD_155\, \EVENT_DWORD_17[17]\, N_292, 
        \EVENT_DWORD_17_i_0_0[17]_net_1\, N_291, 
        \EVENT_DWORD_154\, \EVENT_DWORD_17[16]\, N_1660, 
        \EVENT_DWORD_17_i_0_0[16]_net_1\, N_1661, 
        \EVENT_DWORD_153\, \EVENT_DWORD_17[15]\, N_1624, 
        \EVENT_DWORD_17_i_0_0[15]_net_1\, N_1623, 
        \EVENT_DWORD_152\, \EVENT_DWORD_17[14]\, N_1657, 
        \EVENT_DWORD_17_i_0_0[14]_net_1\, N_1658, 
        \EVENT_DWORD_151\, \EVENT_DWORD_17[13]\, N_339, 
        \EVENT_DWORD_17_i_0_0[13]_net_1\, N_338, 
        \EVENT_DWORD_150\, \EVENT_DWORD_17[12]\, N_1654, 
        \EVENT_DWORD_17_i_0_0[12]_net_1\, N_1655, 
        \EVENT_DWORD_149\, \EVENT_DWORD_17[11]\, N_336, 
        \EVENT_DWORD_17_i_0_0[11]_net_1\, N_335, 
        \EVENT_DWORD_148\, \EVENT_DWORD_17[10]\, N_1651, 
        \EVENT_DWORD_17_i_0_0[10]_net_1\, N_1652, 
        \EVENT_DWORD_147\, \EVENT_DWORD_17[9]\, un1_STATE1_18, 
        N_295, \EVENT_DWORD_17_i_0[9]_net_1\, N_294, N_190_i, 
        N_1229_i, \EVENT_DWORD_146\, \EVENT_DWORD_17[8]\, N_1663, 
        \EVENT_DWORD_17_i_0_0[8]_net_1\, N_1664, 
        \EVENT_DWORD_145\, \EVENT_DWORD_17[7]\, N_1621, 
        \EVENT_DWORD_17_i_0_0[7]_net_1\, N_105_i_0, N_1620, 
        \EVENT_DWORD_144\, \EVENT_DWORD_17[6]\, N_1648, 
        \EVENT_DWORD_17_i_0_0[6]_net_1\, N_1649, 
        \EVENT_DWORD_143\, \EVENT_DWORD_17[5]\, N_333, 
        \EVENT_DWORD_17_i_0_0[5]_net_1\, N_332, \EVENT_DWORD_142\, 
        \EVENT_DWORD_17[4]\, N_326, 
        \EVENT_DWORD_17_i_0_0[4]_net_1\, N_327, \EVENT_DWORD_141\, 
        \EVENT_DWORD_17[3]\, N_1618, 
        \EVENT_DWORD_17_i_0_0[3]_net_1\, N_1616, 
        \EVENT_DWORD_140\, \EVENT_DWORD_17[2]\, N_1644, 
        \EVENT_DWORD_17_i_0_0[2]_net_1\, N_1645, 
        \EVENT_DWORD_139\, \EVENT_DWORD_17[1]\, N_330, 
        \EVENT_DWORD_17_i_0_0[1]_net_1\, N_329, \EVENT_DWORD_138\, 
        \EVENT_DWORD_17[0]\, N_1641, 
        \EVENT_DWORD_17_i_0_0[0]_net_1\, N_1642, N_1753, N_304, 
        \I2C_RREQ_137\, \STATE1_d_i[7]_net_1\, 
        un1_I2C_RREQ_1_sqmuxa, N_293, N_1592, \PDL_RREQ_136\, 
        un1_STATE1_1_sqmuxa, \CHIP_ADDR_135\, N_96, 
        I2C_RREQ_1_sqmuxa, N_7192_i, \un2_i2c_chain_0_0_0_2_i[3]\, 
        \un2_i2c_chain_0_0_0_1_i[3]\, N_1691_1, N_312, N_312_1, 
        N_1633, \un2_i2c_chain_0_0_0_a2_4[3]_net_1\, N_300, 
        N_1769, N_216, N_1603, N_186, N_219, N_1770, 
        \un2_i2c_chain_0_0_0_a2_1_0[3]_net_1\, N_194, N_1775, 
        \CHIP_ADDR_134\, N_721_i_0, \un2_i2c_chain_0_i_0_3_i[2]\, 
        N_298_i, \un2_i2c_chain_0_i_0_2_i[2]\, 
        \un2_i2c_chain_0_i_0_0[2]_net_1\, N_1629_1, N_1774, N_213, 
        N_1763, N_202_i_i_0, \un2_i2c_chain_0_i_0_1[2]_net_1\, 
        N_1765, N_189, N_1766, N_1773, \CHIP_ADDR_133\, N_94, 
        \un2_i2c_chain_0_0_0_3_i[1]\, 
        \un2_i2c_chain_0_0_0_0_i[1]\, N_1776, N_218, N_1630_i, 
        N_1638_1, \un2_i2c_chain_0_0_0_1[1]_net_1\, N_1631, 
        N_1764, \CHANNEL_132\, N_99, \un2_i2c_chain_0_0_0_0_i[6]\, 
        N_1637_i, N_1639_i, N_1612, N_1640, N_197, \CHANNEL_131\, 
        N_98, \un2_i2c_chain_0_0_0_0_3_i[5]\, 
        \un2_i2c_chain_0_0_0_0_0_i[5]\, N_1725_i, N_265_i_i_0_i, 
        \un2_i2c_chain_0_0_0_a2_11[5]_net_1\, 
        \un2_i2c_chain_0_0_0_0_1_tz[5]_net_1\, 
        \un2_i2c_chain_0_0_0_1_0_i[5]\, 
        \un2_i2c_chain_0_0_0_a2_9_0[5]_net_1\, N_1767, N_1724, 
        \CHANNEL_130\, N_97, \un2_i2c_chain_0_0_0_3_i[4]\, 
        \un2_i2c_chain_0_0_0_2_i[4]\, 
        \un2_i2c_chain_0_0_0_1_i[4]\, 
        \un2_i2c_chain_0_0_0_a2_1[4]_net_1\, N_1615_i, 
        \un2_i2c_chain_0_0_0_a2_0_i[4]\, N_1688_i, 
        \un2_i2c_chain_0_0_0_0[4]_net_1\, N_1692, \WRB_129\, 
        N_182, \WRB\, N_697, N_305, N_306, N_1541_i, 
        \I2C_CHAIN_128\, N_93, N_1674, \FAULT_STAT_126\, 
        \FAULT_STAT_3\, \FAULT_STAT_1_sqmuxa\, \FAULT_STROBE\, 
        FAULT_STROBE_0_i, \EVNT_TRG_125\, N_1147, 
        \STATE2[0]_net_1\, \CRC32_124\, N_1222, N_276_i_i_0, 
        \CRC32_123\, N_1294, N_260_i_i_0, \CRC32_122\, N_1594, 
        N_248_i_i_0, \CRC32_121\, N_1385, N_264_i_i_0, 
        \CRC32_120\, N_1142, N_242_i_i_0, \CRC32_119\, N_1384, 
        N_287_i_i_0, \CRC32_118\, N_1141, N_1780_i_0, \CRC32_117\, 
        N_1293, N_279_i_i_0, \CRC32_116\, N_1221, N_1781_i_0, 
        \CRC32_115\, N_1292, N_1782_i_0, \CRC32_114\, N_1220, 
        N_275_i_i_0, \CRC32_113\, N_1383, N_286_i_i_0, 
        \CRC32_112\, N_1468, N_273_i_i_0, \CRC32_111\, N_1382, 
        N_285_i_i_0, \CRC32_110\, N_1140, N_1779_i_0, \CRC32_109\, 
        N_1381, N_1783_i_0, \CRC32_108\, N_1219, N_251_i_i_0, 
        \CRC32_107\, N_1291, N_257_i_i_0, \CRC32_106\, N_1380, 
        N_284_i_i_0, \CRC32_105\, N_1290, N_256_i_i_0, 
        \CRC32_104\, N_1218, N_250_i_i_0, \CRC32_103\, N_1289, 
        N_278_i_i_0, \CRC32_102\, N_1379, N_1469, N_283_i_i_0, 
        \CRC32_101\, N_1378, N_282_i_i_0, \CRC32_100\, N_1596, 
        N_249_i_i_0, \CRC32_99\, N_1377, N_281_i_i_0, \CRC32_98\, 
        N_1376, N_280_i_i_0, \CRC32_97\, N_1216, N_274_i_i_0, 
        \CRC32_96\, N_1123, N_272_i_i_0, \CRC32_95\, N_1375, 
        N_261_i_i_0, \CRC32_94\, N_1288, N_277_i_i_0, \CRC32_93\, 
        N_1287, N_532_3, N_254_i_i_0, \READ_PDL_FLAG_92_0_0\, 
        N_1671, \READ_PDL_FLAG_92_0_0_0\, N_1669_i, N_266, 
        \READ_ADC_FLAG_90_0_0\, N_288_i, N_268_i_0, \CYC_STAT_89\, 
        CLEAR_PSM_FLAGS_i_0, \CYC_STAT_1_sqmuxa\, \CYC_STAT_1\, 
        \FIFO_END_EVNT_88\, un1_STATE1_5, \DTEST_FIFO_87\, N_795, 
        ADD_16x16_slow_I15_Y, ADD_16x16_slow_I15_Y_0, 
        I14_un1_CO1_i_0_i, \REG[47]\, \un2_evread_i_0[14]\, 
        ADD_16x16_slow_I14_un1_CO1_N_16_i_i, 
        ADD_16x16_slow_I14_un1_CO1_N_18, 
        ADD_16x16_slow_I14_un1_CO1_N_17, \un2_evread[14]\, 
        ADD_16x16_slow_I14_un1_CO1_m14_3_i, 
        ADD_16x16_slow_I14_un1_CO1_m14_2_0_i, \REG[46]\, 
        ADD_16x16_slow_I14_un1_CO1_m14_2, 
        ADD_16x16_slow_I14_un1_CO1_m7_4_i, 
        ADD_16x16_slow_I14_un1_CO1_m7_3_i, 
        ADD_16x16_slow_I14_un1_CO1_m7_1, 
        ADD_16x16_slow_I13_CO1_0_a0_5, 
        ADD_16x16_slow_I13_CO1_0_a0_2_i, 
        ADD_16x16_slow_I13_CO1_0_a0_3_i, 
        ADD_16x16_slow_I13_CO1_0_a0_0, ADD_16x16_slow_I13_S, 
        ADD_16x16_slow_I13_S_0, ADD_16x16_slow_I12_un1_CO1_0_tz_0, 
        ADD_16x16_slow_I12_S, ADD_16x16_slow_I12_S_0, 
        ADD_16x16_slow_I11_CO1_0_m5_0_a4_0, 
        ADD_16x16_slow_I11_CO1_0_m5_0_a4, 
        ADD_16x16_slow_I11_CO1_0tt_m3_0_a2, 
        ADD_16x16_slow_I11_CO1_0_m5_0_a4_0_0, 
        ADD_16x16_slow_I11_S, ADD_16x16_slow_I11_S_0, 
        ADD_16x16_slow_I10_S, ADD_16x16_slow_I10_S_0, 
        ADD_16x16_slow_I9_CO1_0_tz_0, ADD_16x16_slow_I9_S, 
        ADD_16x16_slow_I9_S_0, ADD_16x16_slow_I8_un1_CO1_0_tz_0, 
        ADD_16x16_slow_I8_S, ADD_16x16_slow_I8_S_0, 
        ADD_16x16_slow_I7_CO1_0_a0_2_i, 
        ADD_16x16_slow_I7_CO1_0_a0_3_i, \REG[32]\, \REG[33]\, 
        ADD_16x16_slow_I7_S, ADD_16x16_slow_I7_S_0, \REG[34]\, 
        ADD_16x16_slow_I6_un4_CO1_6_tz_0, \REG[35]\, 
        ADD_16x16_slow_I6_un1_CO1_0_a0_0, 
        ADD_16x16_slow_I4_un1_CO1_0_a0_0, ADD_16x16_slow_I6_S, 
        N216, ADD_16x16_slow_I6_S_0, I4_un1_CO1, 
        ADD_16x16_slow_I5_CO1_0, ADD_16x16_slow_I3_CO1_0_a0_1, 
        ADD_16x16_slow_I5_S, ADD_16x16_slow_I5_S_0, N212, 
        ADD_16x16_slow_I4_un1_CO1_0, 
        ADD_16x16_slow_I4_un1_CO1_0_a0_0_0_i, 
        ADD_16x16_slow_I4_un1_CO1_0_a0_1_i, ADD_16x16_slow_I4_S, 
        ADD_16x16_slow_I4_S_0, I2_un1_CO1, 
        ADD_16x16_slow_I3_CO1_0, ADD_16x16_slow_I3_S, 
        ADD_16x16_slow_I3_S_0, N208, ADD_16x16_slow_I2_un1_CO1_0, 
        ADD_16x16_slow_I2_S, ADD_16x16_slow_I2_S_0, 
        ADD_16x16_slow_I1_un3_CO1_0, ADD_16x16_slow_I1_CO1_0, 
        ADD_16x16_slow_I1_S, I0_un1_CO1, ADD_16x16_slow_I1_S_0, 
        ADD_16x16_slow_I0_S, \ORATETMO_7[4]\, N_233, I_22, 
        \ORATETMO_7[3]\, I_21, \ORATETMO_7[2]\, I_20_2, 
        \ORATETMO_7[1]\, I_19, \ORATETMO_7[0]\, 
        \DWACT_ADD_CI_0_partial_sum_1[0]\, N_1576_i, 
        \ORATETMO_7_0_0_a2_0[0]_net_1\, \BNC_LIMIT_2\, 
        un4_bnc_res_NE_16_i, un4_bnc_res_0_i_i, un4_bnc_res_1_i_i, 
        un4_bnc_res_3_i_i, un4_bnc_res_30_i_i, un4_bnc_res_31_i_i, 
        un4_bnc_res_NE_18_i, un4_bnc_res_NE_5_i, 
        un4_bnc_res_NE_6_i, un4_bnc_res_16_i_i, 
        un4_bnc_res_19_i_i, un4_bnc_res_22_i_i, 
        un4_bnc_res_25_i_i, un4_bnc_res_NE_7_i, un4_bnc_res_5_i_i, 
        un4_bnc_res_7_i_i, un4_bnc_res_10_i_i, un4_bnc_res_13_i_i, 
        un4_bnc_res_NE_27_i, un4_bnc_res_NE_21_i, 
        un4_bnc_res_NE_22_i, un4_bnc_res_NE_9_i, 
        un4_bnc_res_18_i_i, un4_bnc_res_21_i_i, 
        un4_bnc_res_24_i_i, un4_bnc_res_27_i_i, 
        un4_bnc_res_NE_11_i, un4_bnc_res_8_i_i, un4_bnc_res_9_i_i, 
        un4_bnc_res_12_i_i, un4_bnc_res_15_i_i, 
        un4_bnc_res_NE_20_i, un4_bnc_res_NE_14_i, 
        un4_bnc_res_NE_15_i, un4_bnc_res_NE_1_i, 
        un4_bnc_res_20_i_i, un4_bnc_res_23_i_i, 
        un4_bnc_res_26_i_i, un4_bnc_res_29_i_i, un4_bnc_res_2_i_i, 
        un4_bnc_res_14_i_i, un4_bnc_res_17_i_i, 
        un4_bnc_res_NE_13_i, un4_bnc_res_28_i_i, 
        un4_bnc_res_11_i_i, un4_bnc_res_4_i_i, un4_bnc_res_6_i_i, 
        \FAULT_STROBE_2\, \CYC_STAT_1_2\, \CYC_STAT_0\, 
        \CYC_STAT_0_2\, \BNC_LIMIT_stretched_1\, \BNC_LIMIT\, 
        \BNC_LIMIT_r\, \L2RS_1\, \L2RF1\, \L2RF2\, \L2RF3\, 
        \L2AS_1\, \L2AF1\, \L2AF2\, \L2AF3\, \L1AS_1\, \L1AF1\, 
        \L1AF2\, \L1AF3\, \BNC_LIMIT_stretched\, \REG[334]\, 
        OR_RREQ_net_1, \EVRDY_c\, I2C_RREQ_net_1, PDL_RREQ_net_1, 
        I2C_CHAIN_net_1, \REG[20]\, DTEST_FIFO_net_1, 
        \CHIP_ADDR[0]_net_1\, \CHIP_ADDR[1]_net_1\, 
        \CHIP_ADDR[2]_net_1\, \CHANNEL[0]_net_1\, 
        \CHANNEL[1]_net_1\, \CHANNEL[2]_net_1\, 
        \PDL_RADDR[0]_net_1\, \PDL_RADDR[1]_net_1\, 
        \PDL_RADDR[2]_net_1\, \PDL_RADDR[3]_net_1\, 
        \PDL_RADDR[4]_net_1\, \PDL_RADDR[5]_net_1\, 
        \OR_RADDR[0]_net_1\, \OR_RADDR[1]_net_1\, 
        \OR_RADDR[2]_net_1\, \OR_RADDR[3]_net_1\, 
        \OR_RADDR[4]_net_1\, \OR_RADDR[5]_net_1\, 
        \DWACT_ADD_CI_0_partial_sum_2[0]\, \EVNT_NUM_2[1]\, 
        \EVNT_NUM_2[2]\, \EVNT_NUM_2[3]\, \EVNT_NUM_2[4]\, 
        \EVNT_NUM_2[5]\, \EVNT_NUM_2[6]\, \EVNT_NUM_2[7]\, 
        \EVNT_NUM_2[8]\, \EVNT_NUM_2[9]\, \EVNT_NUM_2[10]\, 
        \EVNT_NUM_2[11]\, \DWACT_ADD_CI_0_TMP_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\, N_4, 
        \DWACT_FINC_E[24]\, \DWACT_FINC_E[23]\, 
        \DWACT_FINC_E[27]\, \DWACT_FINC_E[26]\, N_9, N_14, 
        \DWACT_FINC_E[25]\, N_19_0, \DWACT_FINC_E[29]\, 
        \DWACT_FINC_E[30]\, N_24, \DWACT_FINC_E[15]\, 
        \DWACT_FINC_E[17]\, \DWACT_FINC_E[22]\, N_31, 
        \DWACT_FINC_E[21]\, \DWACT_FINC_E[9]\, \DWACT_FINC_E[12]\, 
        \DWACT_FINC_E[20]\, N_40, \DWACT_FINC_E[13]\, 
        \DWACT_FINC_E[19]\, N_45, \DWACT_FINC_E[18]\, N_52, 
        \DWACT_FINC_E[33]\, \DWACT_FINC_E[34]\, \DWACT_FINC_E[2]\, 
        \DWACT_FINC_E[5]\, N_61, \DWACT_FINC_E[28]\, 
        \DWACT_FINC_E[16]\, N_66, N_71, \DWACT_FINC_E[14]\, N_76, 
        N_81_0, \DWACT_FINC_E[10]\, N_88, \DWACT_FINC_E[11]\, 
        N_93_0, N_98_0, N_103, \DWACT_FINC_E[8]\, N_108, N_116, 
        N_123, \DWACT_FINC_E[3]\, N_131, N_136, N_141, 
        \DWACT_FINC_E[1]\, N_146, N_154, 
        \DWACT_ADD_CI_0_pog_array_1_4[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\, 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, 
        \DWACT_ADD_CI_0_g_array_1_1_0[0]\, 
        \DWACT_ADD_CI_0_pog_array_0[0]\, 
        \DWACT_ADD_CI_0_TMP_2[0]\, 
        \DWACT_ADD_CI_0_g_array_0_1[0]\, 
        \DWACT_ADD_CI_0_g_array_12_5[0]\, 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, 
        \DWACT_ADD_CI_0_g_array_0_3[0]\, 
        \DWACT_ADD_CI_0_partial_sum[4]\, 
        \DWACT_ADD_CI_0_partial_sum[3]\, 
        \DWACT_ADD_CI_0_partial_sum[2]\, 
        \DWACT_ADD_CI_0_partial_sum[1]\, \GND\, \VCC\
         : std_logic;

    for all : event_fifo
	Use entity work.event_fifo(DEF_ARCH);
begin 

    un2_evread_0 <= \un2_evread[14]\;
    CHANNEL(2) <= \CHANNEL[2]_net_1\;
    CHANNEL(1) <= \CHANNEL[1]_net_1\;
    CHANNEL(0) <= \CHANNEL[0]_net_1\;
    CHIP_ADDR(2) <= \CHIP_ADDR[2]_net_1\;
    CHIP_ADDR(1) <= \CHIP_ADDR[1]_net_1\;
    CHIP_ADDR(0) <= \CHIP_ADDR[0]_net_1\;
    OR_RADDR(5) <= \OR_RADDR[5]_net_1\;
    OR_RADDR(4) <= \OR_RADDR[4]_net_1\;
    OR_RADDR(3) <= \OR_RADDR[3]_net_1\;
    OR_RADDR(2) <= \OR_RADDR[2]_net_1\;
    OR_RADDR(1) <= \OR_RADDR[1]_net_1\;
    OR_RADDR(0) <= \OR_RADDR[0]_net_1\;
    PDL_RADDR(5) <= \PDL_RADDR[5]_net_1\;
    PDL_RADDR(4) <= \PDL_RADDR[4]_net_1\;
    PDL_RADDR(3) <= \PDL_RADDR[3]_net_1\;
    PDL_RADDR(2) <= \PDL_RADDR[2]_net_1\;
    PDL_RADDR(1) <= \PDL_RADDR[1]_net_1\;
    PDL_RADDR(0) <= \PDL_RADDR[0]_net_1\;
    REG_329 <= \REG[334]\;
    REG_41 <= \REG[46]\;
    REG_42 <= \REG[47]\;
    REG_15 <= \REG[20]\;
    REG_27 <= \REG[32]\;
    REG_28 <= \REG[33]\;
    REG_30 <= \REG[35]\;
    REG_29 <= \REG[34]\;
    REG_39 <= \REG[44]\;
    REG_37 <= \REG[42]\;
    REG_36 <= \REG[41]\;
    REG_34 <= \REG[39]\;
    REG_33 <= \REG[38]\;
    REG_38 <= \REG[43]\;
    REG_35 <= \REG[40]\;
    REG_40 <= \REG[45]\;
    REG_31 <= \REG[36]\;
    REG_32 <= \REG[37]\;
    DTEST_FIFO <= DTEST_FIFO_net_1;
    I2C_CHAIN <= I2C_CHAIN_net_1;
    PDL_RREQ <= PDL_RREQ_net_1;
    I2C_RREQ <= I2C_RREQ_net_1;
    EVRDY_c <= \EVRDY_c\;
    OR_RREQ <= OR_RREQ_net_1;
    EVNT_TRG <= EVNT_TRG_net_1;

    \FID[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_188\, CLR => CLEAR_13, Q
         => \FID[18]_net_1\);
    
    \CNT_8_i[4]\ : AND2
      port map(A => N_185_i, B => I_24_2, Y => N_84);
    
    \CNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_8_i[0]_net_1\, CLR => 
        CLEAR_5, Q => \CNT[0]_net_1\);
    
    \FID[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_182\, CLR => CLEAR_13, Q
         => \FID[12]_net_1\);
    
    STATE1_tr9_i_o3_1_i_a2_0_a2_0_a2 : NOR2FT
      port map(A => \STATE1_0[1]_net_1\, B => \STATE1_0[2]_net_1\, 
        Y => N_166);
    
    \FID_6_0_iv_0_0_a2[30]\ : NOR2
      port map(A => N_1574, B => REG_73, Y => N_1515);
    
    \STATE1_ns_i_0_1[1]\ : NOR3
      port map(A => N_1562_i, B => N_1568_i, C => N_1563_i, Y => 
        \STATE1_ns_i_0_1[1]_net_1\);
    
    \EVENT_DWORD_17_r[19]\ : AND3FFT
      port map(A => N_1676, B => \EVENT_DWORD_17_i_0[19]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[19]\);
    
    un1_EVENT_DWORD_0_sqmuxa_0_0_a2_1 : AND2
      port map(A => I2C_RACK, B => \STATE1[0]_net_1\, Y => N_1593);
    
    \EVENT_DWORD_17_r[25]\ : AND3FFT
      port map(A => N_1737, B => \EVENT_DWORD_17_i_0_1[25]_net_1\, 
        C => N_532_3_6, Y => \EVENT_DWORD_17[25]\);
    
    \EVENT_DWORD_17_r[10]\ : AND3FFT
      port map(A => N_1651, B => \EVENT_DWORD_17_i_0_0[10]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[10]\);
    
    \CRC32_2_i_0_x2[27]\ : XOR2FT
      port map(A => \CRC32[27]_net_1\, B => 
        \EVENT_DWORD[27]_net_1\, Y => N_242_i_i_0);
    
    \BNC_CNT[28]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_244\, CLR => 
        CLEAR_4, Q => \BNC_CNT[28]_net_1\);
    
    \BNC_CNT_3[4]\ : AND2
      port map(A => I_20_1, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[4]_net_1\);
    
    \CRC32_2_i_0_x2[20]\ : XOR2FT
      port map(A => \CRC32[20]_net_1\, B => 
        \EVENT_DWORD[20]_net_1\, Y => N_286_i_i_0);
    
    \un2_i2c_chain_0_0_0_a2[0]\ : NOR3FFT
      port map(A => \CNT_0[4]_net_1\, B => \CNT_0[5]_net_1\, C
         => N_1766, Y => N_1674);
    
    \ORATETMO_7_0_0_o2[0]\ : NAND3FTT
      port map(A => N_1576_i, B => N_1564, C => N_532_3, Y => 
        N_233);
    
    FID_175 : MUX2H
      port map(A => \FID[5]_net_1\, B => \FID_6[5]\, S => N_205, 
        Y => \FID_175\);
    
    un2_bnc_cnt_I_23 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \BNC_CNT[3]_net_1\, C
         => \BNC_CNT[4]_net_1\, Y => N_146);
    
    \CRC32[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_101\, CLR => CLEAR_8, 
        Q => \CRC32[8]_net_1\);
    
    \BNC_CNT_3[25]\ : AND2
      port map(A => I_173, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[25]_net_1\);
    
    \FID[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_189\, CLR => CLEAR_13, Q
         => \FID[19]_net_1\);
    
    \FID_6_iv_0_0_a2_0[4]\ : OR2FT
      port map(A => REG_47, B => N_1574_0, Y => N_342);
    
    \FID_6_iv_0_0_0[11]\ : OAI21
      port map(A => N_1575_0, B => \FID_2_i[11]\, C => N_1474, Y
         => \FID_6_iv_0_0_0_i[11]\);
    
    \EVNT_NUM[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[8]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[8]_net_1\);
    
    EVENT_DWORD_139 : MUX2H
      port map(A => \EVENT_DWORD[1]_net_1\, B => 
        \EVENT_DWORD_17[1]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_139\);
    
    CYC_STAT_0_2 : NOR2FT
      port map(A => REG_c(21), B => \CLEAR_PSM_FLAGS\, Y => 
        \CYC_STAT_0_2\);
    
    \un2_i2c_chain_0_0_0_a2_2[6]\ : OR3FFT
      port map(A => N_1764, B => N_194, C => \CNT_0[0]_net_1\, Y
         => N_1640);
    
    un1_REG_1_ADD_16x16_slow_I6_un1_CO1_0_a0_2_0 : NOR3FFT
      port map(A => ADD_16x16_slow_I6_un1_CO1_0_a0_0, B => 
        ADD_16x16_slow_I4_un1_CO1_0_a0_0, C => \REG[33]\, Y => 
        ADD_16x16_slow_I6_un1_CO1_0_a0_2);
    
    \STATE1_ns_1_iv_0_m2_i_m2[0]\ : MUX2H
      port map(A => PULSE(3), B => N_1470_i_0, S => 
        \STATE1[1]_net_1\, Y => N_1613);
    
    \EVENT_DWORD_17_i_o2_1_a3[7]\ : OR2FT
      port map(A => N_304, B => \OR_RACK_sync\, Y => N_1753);
    
    EVENT_DWORD_160 : MUX2H
      port map(A => \EVENT_DWORD[22]_net_1\, B => 
        \EVENT_DWORD_17[22]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_160\);
    
    \EVENT_DWORD_17_i_0_a2[12]\ : NOR2
      port map(A => \EVENT_DWORD[12]_net_1\, B => N_1229_i_1, Y
         => N_1654);
    
    \BNC_CNT[12]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_228\, CLR => 
        CLEAR_2, Q => \BNC_CNT[12]_net_1\);
    
    \un2_i2c_chain_0_0_0_0[5]\ : OR3
      port map(A => \un2_i2c_chain_0_0_0_0_3_i[5]\, B => 
        \un2_i2c_chain_0_0_0_0_0_i[5]\, C => N_1725_i, Y => N_98);
    
    PDL_RADDR_214 : MUX2H
      port map(A => \CNT[4]_net_1\, B => \PDL_RADDR[4]_net_1\, S
         => STATE1_1_sqmuxa_1, Y => \PDL_RADDR_214\);
    
    \EVENT_DWORD[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_169\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[31]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I1_S : XOR2FT
      port map(A => I0_un1_CO1, B => ADD_16x16_slow_I1_S_0, Y => 
        ADD_16x16_slow_I1_S);
    
    un1_REG_1_G_11_0_a2_0 : OAI21
      port map(A => I_8, B => \REG[42]\, C => N224, Y => 
        G_11_0_a2_0);
    
    \OR_RADDR_3_i_0[5]\ : AND2
      port map(A => N_532_3_3, B => \CNT_0[5]_net_1\, Y => N_679);
    
    \CRC32_2_i_0_x2[16]\ : XOR2FT
      port map(A => \CRC32[16]_net_1\, B => 
        \EVENT_DWORD[16]_net_1\, Y => N_1783_i_0);
    
    \un2_i2c_chain_0_0_0_1[3]\ : OAI21FTT
      port map(A => N_1691_1, B => N_199, C => N_312, Y => 
        \un2_i2c_chain_0_0_0_1_i[3]\);
    
    L2AF1 : DFFC
      port map(CLK => ALICLK_c, D => L2A_c_c, CLR => HWRES_c_12, 
        Q => \L2AF1\);
    
    un1_REG_1_ADD_16x16_slow_I1_CO1 : OAI21FTT
      port map(A => ADD_16x16_slow_I1_un3_CO1_0, B => 
        \un2_evread[15]_net_1\, C => ADD_16x16_slow_I1_CO1_0, Y
         => N208);
    
    un1_ORATETMO_1_I_5 : AND2
      port map(A => \ORATETMO_i_i[1]\, B => N_701_i_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_1[0]\);
    
    \EVENT_DWORD_17_i_0_1[26]\ : OAI21FTF
      port map(A => N_1454, B => OR_RDATA(6), C => 
        \EVENT_DWORD_17_i_0_0[26]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[26]_net_1\);
    
    \FID_6_iv_0_0_a2_0[12]\ : OR2FT
      port map(A => REG_55, B => N_1574_0, Y => N_1507);
    
    \FID_6_0_iv_0_a2_2_0_a2[3]\ : OR2
      port map(A => \STATE1_0[3]_net_1\, B => N_176, Y => N_1574);
    
    \CRC32_2_i_0_x2[13]\ : XOR2FT
      port map(A => \CRC32[13]_net_1\, B => 
        \EVENT_DWORD[13]_net_1\, Y => N_284_i_i_0);
    
    un1_REG_1_ADD_16x16_slow_I7_CO1_0_a0_2 : OR3
      port map(A => ADD_16x16_slow_I5_CO1_0_a0_0, B => \REG[39]\, 
        C => \REG[38]\, Y => ADD_16x16_slow_I7_CO1_0_a0_2_i);
    
    un1_ORATETMO_1_I_17 : XOR2
      port map(A => \ORATETMO_i_i[0]\, B => N_701_i_0, Y => 
        \DWACT_ADD_CI_0_partial_sum_1[0]\);
    
    \FID[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_197\, CLR => CLEAR_14, Q
         => \FID[27]_net_1\);
    
    \ORATETMO[4]\ : DFFS
      port map(CLK => CLK_c_c, D => \ORATETMO_7[4]\, SET => 
        CLEAR_16, Q => \ORATETMO[4]_net_1\);
    
    un2_bnc_cnt_I_65 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \BNC_CNT[9]_net_1\, C
         => \BNC_CNT[10]_net_1\, Y => N_116);
    
    \CRC32[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_99\, CLR => CLEAR_8, Q
         => \CRC32[6]_net_1\);
    
    un4_bnc_res_NE_6 : OR2
      port map(A => un4_bnc_res_16_i_i, B => un4_bnc_res_19_i_i, 
        Y => un4_bnc_res_NE_6_i);
    
    EVNT_NUM_2_I_69 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2[0]\);
    
    \EVENT_DWORD_17_i_0_a2[21]\ : NOR2
      port map(A => \EVENT_DWORD[21]_net_1\, B => N_1229_i_0, Y
         => N_1718);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m15 : MUX2H
      port map(A => ADD_16x16_slow_I14_un1_CO1_N_18, B => 
        ADD_16x16_slow_I14_un1_CO1_N_17, S => \un2_evread[14]\, Y
         => ADD_16x16_slow_I14_un1_CO1_N_16_i_i);
    
    \EVENT_DWORD_17_i_0_o2[3]\ : NOR2FT
      port map(A => N_1768_i, B => N_1454_0, Y => N_190_i);
    
    \FID_2[8]\ : XOR2
      port map(A => \CRC32[4]_net_1\, B => \FID_2_0[8]_net_1\, Y
         => \FID_2[8]_net_1\);
    
    \STATE1_ns_1_iv_0_0[2]\ : AO21TTF
      port map(A => N_1777, B => \STATE1[2]_net_1\, C => 
        \STATE1_ns_1_iv_0_0_7[2]_net_1\, Y => \STATE1_ns[2]\);
    
    FIFO_END_EVNT_88 : MUX2H
      port map(A => \FIFO_END_EVNT\, B => N_532_3, S => 
        un1_STATE1_5, Y => \FIFO_END_EVNT_88\);
    
    \FID[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_179\, CLR => CLEAR_15, Q
         => \FID[9]_net_1\);
    
    \OR_RREQ\ : DFFC
      port map(CLK => CLK_c_c, D => \OR_RREQ_203\, CLR => 
        CLEAR_17, Q => OR_RREQ_net_1);
    
    \CRC32[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_107\, CLR => CLEAR_6, 
        Q => \CRC32[14]_net_1\);
    
    \EVENT_DWORD_17_i_0_0[22]\ : OAI21TTF
      port map(A => \EVENT_DWORD[30]_net_1\, B => N_105_i_0_0, C
         => N_1711, Y => \EVENT_DWORD_17_i_0_0[22]_net_1\);
    
    \EVENT_DWORD[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_156\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[18]_net_1\);
    
    un2_bnc_cnt_I_136 : XOR2
      port map(A => N_66, B => \BNC_CNT[21]_net_1\, Y => I_136);
    
    un1_ORATETMO_1_I_28 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_4[0]\);
    
    \FID_6_r[28]\ : OA21
      port map(A => N_1536_i, B => \FID_6_iv_0_0_0_i[28]\, C => 
        N_532_3_4, Y => \FID_6[28]\);
    
    \CRC32_2_i_0_a2_s[17]\ : NOR2
      port map(A => \STATE1[0]_net_1\, B => \STATE1[3]_net_1\, Y
         => N_1585);
    
    \CRC32_2_0_a3_i[7]\ : NOR2FT
      port map(A => N_532_3_0, B => N_249_i_i_0, Y => N_1596);
    
    un2_bnc_cnt_I_13 : XOR2
      port map(A => N_154, B => \BNC_CNT[3]_net_1\, Y => I_13_3);
    
    un2_bnc_cnt_I_77 : XOR2
      port map(A => N_108, B => \BNC_CNT[13]_net_1\, Y => I_77_0);
    
    \FID_6_iv_0_0_1[17]\ : OAI21FTT
      port map(A => REG_60, B => N_1574_1, C => 
        \FID_6_iv_0_0_0[17]_net_1\, Y => \FID_6_iv_0_0_1_i[17]\);
    
    EVNT_NUM_2_I_54 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \EVNT_NUM[4]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    \un2_i2c_chain_0_0_0[0]\ : OR3
      port map(A => N_1674, B => N_1764, C => N_1773, Y => N_93);
    
    \CRC32_2_i_0[15]\ : NOR2FT
      port map(A => N_532_3_1, B => N_251_i_i_0, Y => N_1219);
    
    \EVENT_DWORD_17_i_a2[29]\ : NOR2
      port map(A => I2C_RDATA(9), B => N_1768_i, Y => N_1682);
    
    un1_I2C_RREQ_1_sqmuxa_0_0_0_i2_i_o2 : NAND2
      port map(A => \STATE1[1]_net_1\, B => \STATE1[2]_net_1\, Y
         => N_215);
    
    \CRC32_2_i_0[25]\ : NOR2FT
      port map(A => N_532_3_2, B => N_1780_i_0, Y => N_1141);
    
    PDL_RADDR_213 : MUX2H
      port map(A => \CNT[3]_net_1\, B => \PDL_RADDR[3]_net_1\, S
         => STATE1_1_sqmuxa_1, Y => \PDL_RADDR_213\);
    
    un5_evread : OR3
      port map(A => un5_evread_11_i, B => un5_evread_8_i, C => 
        un5_evread_7_0_i, Y => un5_evread_i_0);
    
    \un2_i2c_chain_0_i_0_2[2]\ : OAI21
      port map(A => N_186, B => \CNT[3]_net_1\, C => 
        \un2_i2c_chain_0_i_0_0[2]_net_1\, Y => 
        \un2_i2c_chain_0_i_0_2_i[2]\);
    
    \STATE1_ns_i_0_a2_3[1]\ : NOR2FT
      port map(A => \STATE1[0]_net_1\, B => N_522, Y => N_7189_i);
    
    READ_ADC_FLAG_90_0_0_o2 : NOR2
      port map(A => N_258_i_0, B => N_268_i_0, Y => N_288_i);
    
    BNC_CNT_244 : MUX2H
      port map(A => \BNC_CNT[28]_net_1\, B => 
        \BNC_CNT_3[28]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_244\);
    
    \CRC32[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_105\, CLR => CLEAR_6, 
        Q => \CRC32[12]_net_1\);
    
    \OR_RADDR[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \OR_RADDR_204\, CLR => 
        CLEAR_16, Q => \OR_RADDR[0]_net_1\);
    
    \EVENT_DWORD_17_0_a2[30]\ : AND2
      port map(A => N_1590, B => PDL_RDATA(6), Y => 
        \EVENT_DWORD_17[30]\);
    
    un2_bnc_cnt_I_224 : XOR2
      port map(A => N_4, B => \BNC_CNT[31]_net_1\, Y => I_224);
    
    I2C_RREQ_1_sqmuxa_0_a5_0_a2 : NOR2FT
      port map(A => N_1592, B => N_215, Y => I2C_RREQ_1_sqmuxa);
    
    EVENT_DWORD_150 : MUX2H
      port map(A => \EVENT_DWORD[12]_net_1\, B => 
        \EVENT_DWORD_17[12]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_150\);
    
    BNC_CNT_230 : MUX2H
      port map(A => \BNC_CNT[14]_net_1\, B => 
        \BNC_CNT_3[14]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_230\);
    
    un4_bnc_res_NE_16 : OR3
      port map(A => un4_bnc_res_3_i_i, B => un4_bnc_res_30_i_i, C
         => un4_bnc_res_31_i_i, Y => un4_bnc_res_NE_16_i);
    
    \EVENT_DWORD_17_r[12]\ : AND3FFT
      port map(A => N_1654, B => \EVENT_DWORD_17_i_0_0[12]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[12]\);
    
    un4_bnc_res_NE_13 : OR2
      port map(A => un4_bnc_res_4_i_i, B => un4_bnc_res_6_i_i, Y
         => un4_bnc_res_NE_13_i);
    
    \STATE1[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[3]\, CLR => 
        CLEAR_19, Q => \STATE1[3]_net_1\);
    
    \un2_i2c_chain_0_0_0_o2_0[1]\ : OR2
      port map(A => \CNT_0[0]_net_1\, B => \CNT_0[3]_net_1\, Y
         => N_219);
    
    BNC_LIMIT_r : DFFC
      port map(CLK => ALICLK_c, D => \BNC_LIMIT\, CLR => CLEAR_5, 
        Q => \BNC_LIMIT_r\);
    
    \un2_i2c_chain_0_0_0_o2[1]\ : OR2FT
      port map(A => \CNT_0[2]_net_1\, B => \CNT_0[1]_net_1\, Y
         => N_218);
    
    \FID_6_iv_0_0_0[24]\ : OAI21FTT
      port map(A => \EVNT_NUM[8]_net_1\, B => N_1575_1, C => 
        N_1489, Y => \FID_6_iv_0_0_0_i[24]\);
    
    \EVENT_DWORD_17_i_0_a2_0[4]\ : NOR2
      port map(A => \EVENT_DWORD[14]_net_1\, B => N_190_i, Y => 
        N_327);
    
    \BNC_CNT[17]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_233\, CLR => 
        CLEAR_3, Q => \BNC_CNT[17]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I6_un4_CO1_6_tz_0 : AND2
      port map(A => \REG[37]\, B => \REG[35]\, Y => 
        ADD_16x16_slow_I6_un4_CO1_6_tz_0);
    
    EVENT_DWORD_149 : MUX2H
      port map(A => \EVENT_DWORD[11]_net_1\, B => 
        \EVENT_DWORD_17[11]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_149\);
    
    \STATE1_ns_i_0_5[1]\ : NAND3
      port map(A => \STATE1_ns_i_0_4[1]_net_1\, B => 
        \STATE1_ns_i_0_2[1]_net_1\, C => N_1564, Y => 
        \STATE1_ns_i_0_5_i[1]\);
    
    \PDL_RADDR[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RADDR_212\, CLR => 
        CLEAR_17, Q => \PDL_RADDR[2]_net_1\);
    
    un2_bnc_cnt_I_185 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[30]\, 
        C => \DWACT_FINC_E[21]\, Y => N_31);
    
    \FID_6_iv_0_0_a2_1[14]\ : NOR2FT
      port map(A => \EVENT_DWORD[14]_net_1\, B => N_620_4_1, Y
         => N_1511_i);
    
    FID_200 : MUX2H
      port map(A => \FID[30]_net_1\, B => \FID_6[30]\, S => 
        N_205_0, Y => \FID_200\);
    
    FAULT_STAT_126 : MUX2H
      port map(A => \FAULT_STAT_3\, B => \FAULT_STAT\, S => 
        \FAULT_STAT_1_sqmuxa\, Y => \FAULT_STAT_126\);
    
    \STATE1_ns_1_iv_0_0_5[2]\ : NAND3FTT
      port map(A => \STATE1_ns_1_iv_0_0_2_i[2]\, B => 
        \STATE1_ns_1_iv_0_0_3[2]_net_1\, C => 
        \STATE1_ns_0_0_0_i_0[3]_net_1\, Y => 
        \STATE1_ns_1_iv_0_0_5_i[2]\);
    
    un4_bnc_res_14 : XOR2
      port map(A => \BNC_CNT[14]_net_1\, B => REG_418, Y => 
        un4_bnc_res_14_i_i);
    
    \FID_2_0[9]\ : XOR2
      port map(A => \CRC32[17]_net_1\, B => \CRC32[29]_net_1\, Y
         => \FID_2_0[9]_net_1\);
    
    \DTEST_FIFO\ : DFFC
      port map(CLK => CLK_c_c, D => \DTEST_FIFO_87\, CLR => 
        CLEAR_9, Q => DTEST_FIFO_net_1);
    
    \CRC32_2_i_0_a2_7[17]\ : OR2FT
      port map(A => N_1585_0, B => N_176_0, Y => N_532_3_7);
    
    \un2_i2c_chain_0_0_0_a2_1_0[1]\ : AND2
      port map(A => \CNT[5]_net_1\, B => \CNT_0[2]_net_1\, Y => 
        N_1629_1);
    
    \un2_i2c_chain_0_0_0_o2[3]\ : NOR2FT
      port map(A => N_1766, B => N_197, Y => N_194);
    
    \RDY_CNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \RDY_CNT_8_i_0[1]_net_1\, CLR
         => CLEAR_17, Q => \RDY_CNT[1]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2[22]\ : NOR2
      port map(A => \EVENT_DWORD[22]_net_1\, B => N_1229_i_0, Y
         => N_1710);
    
    \un2_i2c_chain_0_0_0_0_1_tz[5]\ : OA21FTT
      port map(A => \CNT[0]_net_1\, B => N_188, C => 
        \un2_i2c_chain_0_0_0_a2_9_0[5]_net_1\, Y => 
        \un2_i2c_chain_0_0_0_0_1_tz[5]_net_1\);
    
    \OR_RADDR[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \OR_RADDR_209\, CLR => 
        CLEAR_16, Q => \OR_RADDR[5]_net_1\);
    
    EVNT_NUM_2_I_46 : XOR2
      port map(A => \EVNT_NUM[10]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_11_1[0]\, Y => \EVNT_NUM_2[10]\);
    
    \EVENT_DWORD_17_i_0_a2_0[17]\ : NOR2
      port map(A => \EVENT_DWORD[17]_net_1\, B => N_1229_i_1, Y
         => N_292);
    
    \un2_i2c_chain_0_0_0_0_x3[5]\ : XOR2FT
      port map(A => \CNT[0]_net_1\, B => N_197, Y => 
        N_265_i_i_0_i);
    
    \EVENT_DWORD_17_i_0_a2_0[20]\ : NOR2
      port map(A => I2C_RDATA(0), B => N_1768_i, Y => N_1703);
    
    \EVENT_DWORD_17_i_0_0[14]\ : OAI21TTF
      port map(A => \EVENT_DWORD[22]_net_1\, B => N_105_i_0_1, C
         => N_1658, Y => \EVENT_DWORD_17_i_0_0[14]_net_1\);
    
    \BNC_CNT_3[15]\ : AND2
      port map(A => I_91_0, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[15]_net_1\);
    
    \FID_2_0[6]\ : XOR2
      port map(A => \CRC32[14]_net_1\, B => \CRC32[26]_net_1\, Y
         => \FID_2_0[6]_net_1\);
    
    EVENT_DWORD_162 : MUX2H
      port map(A => \EVENT_DWORD[24]_net_1\, B => 
        \EVENT_DWORD_17[24]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_162\);
    
    READ_OR_FLAG_91_i_0_a2_0 : NOR2FT
      port map(A => N_252, B => \READ_OR_FLAG\, Y => N_1540);
    
    \CNT_0[3]\ : DFFC
      port map(CLK => CLK_c_c, D => N_81, CLR => CLEAR_0, Q => 
        \CNT_0[3]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m7_1 : AND2
      port map(A => \REG[42]\, B => \REG[44]\, Y => 
        ADD_16x16_slow_I14_un1_CO1_m7_1);
    
    \RDY_CNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \RDY_CNT_8_i_0[0]_net_1\, CLR
         => CLEAR_17, Q => \RDY_CNT[0]_net_1\);
    
    un2_bnc_cnt_I_182 : AND3
      port map(A => \DWACT_FINC_E[7]\, B => \DWACT_FINC_E[9]\, C
         => \DWACT_FINC_E[12]\, Y => \DWACT_FINC_E[30]\);
    
    \EVENT_DWORD[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_140\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[2]_net_1\);
    
    I2C_RREQ_1_sqmuxa_0_o3_i_a2 : NOR2
      port map(A => N_192, B => N_199, Y => N_1771);
    
    BNC_CNT_229 : MUX2H
      port map(A => \BNC_CNT[13]_net_1\, B => 
        \BNC_CNT_3[13]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_229\);
    
    un2_bnc_cnt_I_9 : XOR2
      port map(A => N_157, B => \BNC_CNT[2]_net_1\, Y => I_9_2);
    
    \EVENT_DWORD_17_i_0_1[25]\ : OAI21FTF
      port map(A => N_1454, B => OR_RDATA(5), C => 
        \EVENT_DWORD_17_i_0_0[25]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[25]_net_1\);
    
    \CNT_8_i_o3_0[0]\ : OA21FTT
      port map(A => N_1758_1, B => N_199, C => N_1757, Y => 
        N_1600);
    
    un2_bnc_cnt_I_143 : XOR2
      port map(A => N_61, B => \BNC_CNT[22]_net_1\, Y => I_143);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m7_3 : NAND3
      port map(A => \REG[40]\, B => \REG[45]\, C => \REG[46]\, Y
         => ADD_16x16_slow_I14_un1_CO1_m7_3_i);
    
    \CRC32[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_104\, CLR => CLEAR_6, 
        Q => \CRC32[11]_net_1\);
    
    \un2_i2c_chain_0_0_0_a2_1[1]\ : OR2FT
      port map(A => N_1764, B => \CNT_0[1]_net_1\, Y => N_1631);
    
    \STATE1_0[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns_i_0[1]_net_1\, CLR
         => CLEAR_0, Q => \STATE1_0[1]_net_1\);
    
    \BNC_CNT[1]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_217\, CLR => 
        CLEAR_3, Q => \BNC_CNT[1]_net_1\);
    
    un1_CNT_1_I_24 : XOR2
      port map(A => \CNT[4]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => I_24_2);
    
    \EVENT_DWORD_17_i_0_1[28]\ : OAI21FTF
      port map(A => N_1454, B => OR_RDATA(8), C => 
        \EVENT_DWORD_17_i_0_0[28]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[28]_net_1\);
    
    un4_bnc_res_24 : XOR2
      port map(A => \BNC_CNT[24]_net_1\, B => REG_428, Y => 
        un4_bnc_res_24_i_i);
    
    \un2_i2c_chain_0_0_0_a2_3_1[4]\ : NOR2FT
      port map(A => \CNT_0[0]_net_1\, B => N_186, Y => N_1691_1);
    
    FID_172 : MUX2H
      port map(A => \FID[2]_net_1\, B => \FID_6[2]\, S => N_205, 
        Y => \FID_172\);
    
    \ORATETMO[0]\ : DFFS
      port map(CLK => CLK_c_c, D => \ORATETMO_7[0]\, SET => 
        CLEAR_16, Q => \ORATETMO_i_i[0]\);
    
    un1_STATE1_1_sqmuxa_0_0_o2 : NOR2FT
      port map(A => \STATE1_0[3]_net_1\, B => \PDL_RACK_sync\, Y
         => N_207);
    
    \STATE1[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[2]\, CLR => 
        CLEAR_19, Q => \STATE1[2]_net_1\);
    
    \FID_6_iv_0_0_x2[13]\ : XOR2FT
      port map(A => \CRC32[9]_net_1\, B => \CRC32[21]_net_1\, Y
         => N_269_i_0_i);
    
    \EVENT_DWORD_17_i_0_a2[1]\ : NOR2
      port map(A => \EVENT_DWORD[11]_net_1\, B => N_190_i, Y => 
        N_329);
    
    \CRC32_2_i_0_a2_0[17]\ : OR2FT
      port map(A => N_1585, B => N_176_0, Y => N_532_3_0);
    
    un4_bnc_res_NE_24 : OR3
      port map(A => un4_bnc_res_NE_16_i, B => un4_bnc_res_0_i_i, 
        C => un4_bnc_res_1_i_i, Y => un4_bnc_res_NE_24_i);
    
    un1_REG_1_ADD_16x16_slow_I11_CO1_0_m5_0 : OR3FFT
      port map(A => ADD_16x16_slow_I11_CO1_0_m5_0_a4_0, B => 
        ADD_16x16_slow_I11_CO1_0_m5_0_a4, C => \un2_evread_1[14]\, 
        Y => ADD_16x16_slow_I11_CO1_0_m5_0);
    
    \FID[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_172\, CLR => CLEAR_14, Q
         => \FID[2]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2_0[10]\ : NOR2
      port map(A => \EVENT_DWORD[20]_net_1\, B => N_190_i_0, Y
         => N_1652);
    
    \FID_6_iv_0_0[19]\ : OAI21FTT
      port map(A => \EVNT_NUM[3]_net_1\, B => N_1575_1, C => 
        N_323, Y => \FID_6_iv_0_0_i[19]\);
    
    \EVENT_DWORD_17_i_0_0[5]\ : OAI21TTF
      port map(A => \EVENT_DWORD[13]_net_1\, B => N_105_i_0, C
         => N_332, Y => \EVENT_DWORD_17_i_0_0[5]_net_1\);
    
    \CNT_8_i[5]\ : AND2
      port map(A => N_185_i, B => I_26, Y => \CNT_8_i[5]_net_1\);
    
    un2_bnc_cnt_I_94 : AND2
      port map(A => \DWACT_FINC_E[7]\, B => \DWACT_FINC_E[9]\, Y
         => \DWACT_FINC_E[10]\);
    
    \FID[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_195\, CLR => CLEAR_14, Q
         => \FID[25]_net_1\);
    
    EVENT_DWORD_164 : MUX2H
      port map(A => \EVENT_DWORD[26]_net_1\, B => 
        \EVENT_DWORD_17[26]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_164\);
    
    un1_CNT_1_I_30 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \CNT[4]_net_1\, Y => I_30);
    
    \CNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => N_81, CLR => CLEAR_6, Q => 
        \CNT[3]_net_1\);
    
    \BNC_CNT_3[6]\ : AND2
      port map(A => I_31_0, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[6]_net_1\);
    
    \FID[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_191\, CLR => CLEAR_14, Q
         => \FID[21]_net_1\);
    
    \ORATETMO[2]\ : DFFS
      port map(CLK => CLK_c_c, D => \ORATETMO_7[2]\, SET => 
        CLEAR_16, Q => \ORATETMO[2]_net_1\);
    
    \BNC_CNT[31]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_247\, CLR => 
        CLEAR_4, Q => \BNC_CNT[31]_net_1\);
    
    \FID_6_r[0]\ : OA21
      port map(A => N_1500_i, B => \FID_6_0_iv_0_0_0_i[0]\, C => 
        N_532_3_6, Y => \FID_6[0]\);
    
    \FID_6_0_iv_0_0_0[3]\ : OAI21FTT
      port map(A => REG_46, B => N_1574_0, C => N_311, Y => 
        \FID_6_0_iv_0_0_0_i[3]\);
    
    \CRC32[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_124\, CLR => CLEAR_8, 
        Q => \CRC32[31]_net_1\);
    
    \FID_6_iv_0_0_a2_1[16]\ : NOR2FT
      port map(A => \EVENT_DWORD[16]_net_1\, B => N_620_4_1, Y
         => N_1534_i);
    
    \EVENT_DWORD_17_i_0_a2_0[3]\ : NOR2
      port map(A => \EVENT_DWORD[3]_net_1\, B => N_1229_i, Y => 
        N_1618);
    
    \BNC_CNT[14]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_230\, CLR => 
        CLEAR_2, Q => \BNC_CNT[14]_net_1\);
    
    L1AS : DFFC
      port map(CLK => ALICLK_c, D => \L1AS_1\, CLR => HWRES_c_12, 
        Q => REG_328);
    
    \ORATETMO[3]\ : DFFS
      port map(CLK => CLK_c_c, D => \ORATETMO_7[3]\, SET => 
        CLEAR_16, Q => \ORATETMO_i_i[3]\);
    
    EVENT_DWORD_166 : MUX2H
      port map(A => \EVENT_DWORD[28]_net_1\, B => 
        \EVENT_DWORD_17[28]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_166\);
    
    EVENT_DWORD_152 : MUX2H
      port map(A => \EVENT_DWORD[14]_net_1\, B => 
        \EVENT_DWORD_17[14]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_152\);
    
    \FID_6_iv_0_0_a2_1[11]\ : NOR2FT
      port map(A => \EVENT_DWORD[11]_net_1\, B => N_620_4_0, Y
         => N_1475_i);
    
    un1_STATE1_11_0_i : AND3FTT
      port map(A => N_1541_i, B => N_253, C => N_1586, Y => N_182);
    
    \un2_i2c_chain_0_0_0_a3_1[3]\ : OR2
      port map(A => N_1763, B => \CNT_0[3]_net_1\, Y => N_1775);
    
    \STATE1_ns_i_0_4[1]\ : OAI21FTF
      port map(A => N_252, B => N_1195_1, C => N_193, Y => 
        \STATE1_ns_i_0_4[1]_net_1\);
    
    \FID_6_iv_0_0_0[10]\ : OAI21
      port map(A => N_1575_0, B => \FID_2_i[10]\, C => N_1471, Y
         => \FID_6_iv_0_0_0_i[10]\);
    
    \un2_i2c_chain_0_0_0_0[4]\ : OA21FTT
      port map(A => N_189, B => N_199, C => N_1692, Y => 
        \un2_i2c_chain_0_0_0_0[4]_net_1\);
    
    \EVENT_DWORD[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_141\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[3]_net_1\);
    
    FID_189 : MUX2H
      port map(A => \FID[19]_net_1\, B => \FID_6[19]\, S => 
        N_205_1, Y => \FID_189\);
    
    \FID[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_190\, CLR => CLEAR_14, Q
         => \FID[20]_net_1\);
    
    \BNC_CNT_3[2]\ : AND2
      port map(A => I_9_2, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[2]_net_1\);
    
    \FID_6_iv_0_0_a2_2[17]\ : NOR2FT
      port map(A => \EVENT_DWORD[17]_net_1\, B => N_620_4_1, Y
         => N_1555_i);
    
    un2_bnc_cnt_I_66 : XOR2
      port map(A => N_116, B => \BNC_CNT[11]_net_1\, Y => I_66_0);
    
    \CRC32_2_i_0_a2_3[17]\ : OR2FT
      port map(A => N_1585_0, B => N_176_0, Y => N_532_3_3);
    
    \CRC32_2_i_0_x2[26]\ : XOR2FT
      port map(A => \CRC32[26]_net_1\, B => 
        \EVENT_DWORD[26]_net_1\, Y => N_287_i_i_0);
    
    BNC_CNT_240 : MUX2H
      port map(A => \BNC_CNT[24]_net_1\, B => 
        \BNC_CNT_3[24]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_240\);
    
    un2_bnc_cnt_I_62 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[5]\, Y => \DWACT_FINC_E[6]\);
    
    \FID_6_r[14]\ : OA21
      port map(A => N_1511_i, B => \FID_6_iv_0_0_0_i[14]\, C => 
        N_532_3_5, Y => \FID_6[14]\);
    
    \CRC32_2_i_0_x2[8]\ : XOR2FT
      port map(A => \CRC32[8]_net_1\, B => \EVENT_DWORD[8]_net_1\, 
        Y => N_282_i_i_0);
    
    \STATE2_ns_i_i_a2_i[1]\ : AND2
      port map(A => \STATE2[2]_net_1\, B => \TRIGGER_sync\, Y => 
        \STATE2_ns_i_i_a2_i[1]_net_1\);
    
    \STATE1_ns_1_iv_0_0_o3[0]\ : OAI21FTT
      port map(A => N_1752_1, B => N_193, C => 
        \STATE1_ns_1_iv_0_0_o3_4[0]_net_1\, Y => N_1778);
    
    \CRC32_2_i_0_x2[23]\ : XOR2FT
      port map(A => \CRC32[23]_net_1\, B => 
        \EVENT_DWORD[23]_net_1\, Y => N_1781_i_0);
    
    STATE1_tr9_i_a4_0_o2 : NOR2
      port map(A => \L2ASS\, B => PULSE(2), Y => N_1470);
    
    \CRC32[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_97\, CLR => CLEAR_8, Q
         => \CRC32[4]_net_1\);
    
    \BNC_CNT[26]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_242\, CLR => 
        CLEAR_3, Q => \BNC_CNT[26]_net_1\);
    
    \FID_6_iv_0_0_a2_0[10]\ : OR2FT
      port map(A => REG_53, B => N_1574_0, Y => N_1471);
    
    \CRC32_2_i_0[3]\ : NOR2FT
      port map(A => N_532_3_0, B => N_272_i_i_0, Y => N_1123);
    
    un1_REG_1_G_6_0 : OR2
      port map(A => \REG[33]\, B => \REG[32]\, Y => G_6_0);
    
    un5_evread_6 : OR3
      port map(A => \REG[37]\, B => \REG[40]\, C => \REG[36]\, Y
         => un5_evread_6_i);
    
    un1_REG_1_G_0_x2 : XOR2
      port map(A => ADD_16x16_slow_I14_S_0, B => G_0_o2, Y => 
        G_0_x2);
    
    un2_bnc_cnt_I_73 : XOR2
      port map(A => N_111, B => \BNC_CNT[12]_net_1\, Y => I_73_0);
    
    \BNC_CNT[2]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_218\, CLR => 
        CLEAR_4, Q => \BNC_CNT[2]_net_1\);
    
    \BNC_CNT_3[7]\ : AND2
      port map(A => I_38_0, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[7]_net_1\);
    
    READ_OR_FLAG_91_i_0 : NOR3FTT
      port map(A => \STATE1_d[7]\, B => N_1539, C => N_1540, Y
         => \READ_OR_FLAG_91_i_0\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \un2_i2c_chain_0_0_0_a2_9_0[5]\ : OR2FT
      port map(A => \CNT_0[3]_net_1\, B => N_1767, Y => 
        \un2_i2c_chain_0_0_0_a2_9_0[5]_net_1\);
    
    un4_bnc_res_11 : XOR2
      port map(A => \BNC_CNT[11]_net_1\, B => REG_415, Y => 
        un4_bnc_res_11_i_i);
    
    un1_EVENT_DWORD_0_sqmuxa_0_o5_0_a2_0_a2_0_a2_0 : NOR2FT
      port map(A => \OR_RACK_sync\, B => N_1762, Y => N_1454_0);
    
    READ_ADC_FLAG_90_0_0_x2 : XOR2
      port map(A => \STATE1[1]_net_1\, B => \STATE1[3]_net_1\, Y
         => N_268_i_0);
    
    EVENT_DWORD_154 : MUX2H
      port map(A => \EVENT_DWORD[16]_net_1\, B => 
        \EVENT_DWORD_17[16]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_154\);
    
    \ORATETMO_7_0_0[3]\ : OR2
      port map(A => N_233, B => I_21, Y => \ORATETMO_7[3]\);
    
    EVRDYi_202 : MUX2H
      port map(A => EVREAD_i_0, B => \EVRDY_c\, S => \un1_reg154\, 
        Y => \EVRDYi_202\);
    
    \EVENT_DWORD_17_i_0_a2[3]\ : NOR2
      port map(A => \EVENT_DWORD[13]_net_1\, B => N_190_i, Y => 
        N_1616);
    
    \STATE1_ns_0_0_0_o3[3]\ : NOR2
      port map(A => \STATE1[0]_net_1\, B => \STATE1[1]_net_1\, Y
         => N_1601);
    
    \CRC32_2_i_0_a2_6[17]\ : OR2FT
      port map(A => N_1585_0, B => N_176_0, Y => N_532_3_6);
    
    un1_ORATETMO_1_I_14 : XOR2
      port map(A => \ORATETMO_i_i[3]\, B => N_701_i_0_0, Y => 
        \DWACT_ADD_CI_0_partial_sum[3]\);
    
    EVNT_NUM_2_I_72 : AND2
      port map(A => \EVNT_NUM[6]_net_1\, B => \EVNT_NUM[7]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_2[0]\);
    
    un1_reg154 : OAI21FTF
      port map(A => un5_evread_i_0, B => \FIFO_END_EVNT\, C => 
        \un2_evread[15]_net_1\, Y => \un1_reg154\);
    
    CRC32_111 : MUX2H
      port map(A => \CRC32[18]_net_1\, B => N_1382, S => N_1469_1, 
        Y => \CRC32_111\);
    
    un1_REG_1_ADD_16x16_slow_I6_un1_CO1_0_a0_2 : NOR2
      port map(A => \REG[32]\, B => \REG[34]\, Y => 
        ADD_16x16_slow_I2_un1_CO1_0_a0_0);
    
    \CRC32_2_i_0[11]\ : NOR2FT
      port map(A => N_532_3_1, B => N_250_i_i_0, Y => N_1218);
    
    \FID[31]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_201\, CLR => CLEAR_15, Q
         => \FID[31]_net_1\);
    
    EVENT_DWORD_156 : MUX2H
      port map(A => \EVENT_DWORD[18]_net_1\, B => 
        \EVENT_DWORD_17[18]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_156\);
    
    \CRC32_2_i_0[21]\ : NOR2FT
      port map(A => N_532_3_2, B => N_275_i_i_0, Y => N_1220);
    
    un4_bnc_res_NE_25 : OR3
      port map(A => un4_bnc_res_NE_18_i, B => un4_bnc_res_NE_5_i, 
        C => un4_bnc_res_NE_6_i, Y => un4_bnc_res_NE_25_i);
    
    \un2_i2c_chain_0_i_0_a3_1[2]\ : NAND2
      port map(A => \CNT[1]_net_1\, B => \CNT[2]_net_1\, Y => 
        N_1766);
    
    \FID_6_r[4]\ : OA21
      port map(A => N_343_i, B => \FID_6_iv_0_0_0_i[4]\, C => 
        N_532_3_6, Y => \FID_6[4]\);
    
    \EVENT_DWORD_17_i_0_1[21]\ : OAI21FTF
      port map(A => N_1454_0, B => OR_RDATA(1), C => 
        \EVENT_DWORD_17_i_0_0[21]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[21]_net_1\);
    
    CRC32_121 : MUX2H
      port map(A => \CRC32[28]_net_1\, B => N_1385, S => N_1469_0, 
        Y => \CRC32_121\);
    
    un2_bnc_cnt_I_149 : AND3
      port map(A => \BNC_CNT[0]_net_1\, B => \BNC_CNT[1]_net_1\, 
        C => \BNC_CNT[2]_net_1\, Y => \DWACT_FINC_E[34]\);
    
    \OR_RADDR[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \OR_RADDR_207\, CLR => 
        CLEAR_16, Q => \OR_RADDR[3]_net_1\);
    
    \un2_i2c_chain_0_0_0_1_0[5]\ : OAI21FTT
      port map(A => N_213, B => N_1775, C => N_1724, Y => 
        \un2_i2c_chain_0_0_0_1_0_i[5]\);
    
    BNC_CNT_228 : MUX2H
      port map(A => \BNC_CNT[12]_net_1\, B => 
        \BNC_CNT_3[12]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_228\);
    
    \PDL_RREQ\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RREQ_136\, CLR => 
        CLEAR_17, Q => PDL_RREQ_net_1);
    
    \FID_6_0_iv_0_0_a2[31]\ : NOR2FT
      port map(A => REG_74, B => N_1574, Y => N_1497_i);
    
    CHANNEL_130 : MUX2H
      port map(A => \CHANNEL[0]_net_1\, B => N_97, S => 
        I2C_RREQ_1_sqmuxa, Y => \CHANNEL_130\);
    
    \EVENT_DWORD_17_r[5]\ : AND3FFT
      port map(A => N_333, B => \EVENT_DWORD_17_i_0_0[5]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[5]\);
    
    un1_REG_1_ADD_16x16_slow_I0_un1_CO1 : OR2FT
      port map(A => \REG[32]\, B => \un2_evread[15]_net_1\, Y => 
        I0_un1_CO1);
    
    CRC32_115 : MUX2H
      port map(A => \CRC32[22]_net_1\, B => N_1292, S => N_1469_0, 
        Y => \CRC32_115\);
    
    \CNT_8_i[1]\ : AND2
      port map(A => N_185_i, B => I_21_0, Y => \CNT_8_i[1]_net_1\);
    
    BNC_CNT_227 : MUX2H
      port map(A => \BNC_CNT[11]_net_1\, B => 
        \BNC_CNT_3[11]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_227\);
    
    \EVENT_DWORD_17_i_0_0[16]\ : OAI21TTF
      port map(A => \EVENT_DWORD[24]_net_1\, B => N_105_i_0_1, C
         => N_1661, Y => \EVENT_DWORD_17_i_0_0[16]_net_1\);
    
    BNC_CNT_226 : MUX2H
      port map(A => \BNC_CNT[10]_net_1\, B => 
        \BNC_CNT_3[10]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_226\);
    
    un1_REG_1_G_13_i_a2 : NAND2
      port map(A => N220, B => \REG[40]\, Y => I8_un4_CO1);
    
    un4_bnc_res_21 : XOR2
      port map(A => \BNC_CNT[21]_net_1\, B => REG_425, Y => 
        un4_bnc_res_21_i_i);
    
    \FID[30]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_200\, CLR => CLEAR_14, Q
         => \FID[30]_net_1\);
    
    \EVENT_DWORD_17_r[21]\ : AND3FFT
      port map(A => N_1718, B => \EVENT_DWORD_17_i_0_1[21]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[21]\);
    
    \CRC32[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_117\, CLR => CLEAR_7, 
        Q => \CRC32[24]_net_1\);
    
    \EVNT_NUM[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[1]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[1]_net_1\);
    
    \OR_RADDR_3_i_0[2]\ : AND2
      port map(A => N_532_3_3, B => \CNT_0[2]_net_1\, Y => N_685);
    
    STATE1_1_sqmuxa_1_0_a5_0_o3 : OR2FT
      port map(A => N_189, B => N_186, Y => N_192);
    
    \CRC32_2_i_0[31]\ : NOR2FT
      port map(A => N_532_3_2, B => N_276_i_i_0, Y => N_1222);
    
    \REG_1[35]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I3_S, CLR => 
        CLEAR_18, Q => \REG[35]\);
    
    un1_STATE1_17_i_0_0_a2_0 : NOR2FT
      port map(A => \STATE1_0[1]_net_1\, B => N_120_i, Y => N_305);
    
    FID_194 : MUX2H
      port map(A => \FID[24]_net_1\, B => \FID_6[24]\, S => 
        N_205_0, Y => \FID_194\);
    
    \FID_2[7]\ : XOR2FT
      port map(A => \CRC32[3]_net_1\, B => \FID_2_0[7]_net_1\, Y
         => \FID_2_i[7]\);
    
    un2_bnc_cnt_I_209 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \DWACT_FINC_E[25]\, Y => N_14);
    
    \BNC_CNT[10]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_226\, CLR => 
        CLEAR_2, Q => \BNC_CNT[10]_net_1\);
    
    BNC_LIMIT_2 : AND2FT
      port map(A => un4_bnc_res_i, B => LBSP_c(2), Y => 
        \BNC_LIMIT_2\);
    
    un1_ORATETMO_1_I_13 : XOR2
      port map(A => \ORATETMO[4]_net_1\, B => N_701_i_0_0, Y => 
        \DWACT_ADD_CI_0_partial_sum[4]\);
    
    un4_bnc_res_NE_5 : OR2
      port map(A => un4_bnc_res_22_i_i, B => un4_bnc_res_25_i_i, 
        Y => un4_bnc_res_NE_5_i);
    
    \STATE1_ns_i_0_a2_5[1]\ : NOR3FFT
      port map(A => N_1470, B => N_166, C => N_120_i, Y => 
        N_1568_i);
    
    FID_187 : MUX2H
      port map(A => \FID[17]_net_1\, B => \FID_6[17]\, S => 
        N_205_1, Y => \FID_187\);
    
    \STATE1_ns_1_iv_0_0[0]\ : OAI21TTF
      port map(A => N_1586, B => 
        \STATE1_ns_1_iv_0_0_a2_0[0]_net_1\, C => N_1614, Y => 
        \STATE1_ns[0]\);
    
    \CRC32[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_115\, CLR => CLEAR_7, 
        Q => \CRC32[22]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I3_S_0 : XOR2FT
      port map(A => \REG[35]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I3_S_0);
    
    STATE1_tr16_1_0_a2_0_a2_0_a2_0_a2_0 : OR2FT
      port map(A => N_1573, B => N_221, Y => N_620_4_0);
    
    \RDY_CNT_8_i_0[0]\ : AND2
      port map(A => N_267, B => \DWACT_ADD_CI_0_partial_sum_0[0]\, 
        Y => \RDY_CNT_8_i_0[0]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2[14]\ : NOR2
      port map(A => \EVENT_DWORD[14]_net_1\, B => N_1229_i_1, Y
         => N_1657);
    
    OR_RADDR_205 : MUX2H
      port map(A => \OR_RADDR[1]_net_1\, B => N_687, S => N_248, 
        Y => \OR_RADDR_205\);
    
    \I2C_CHAIN\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_CHAIN_128\, CLR => 
        CLEAR_15, Q => I2C_CHAIN_net_1);
    
    BNC_CNT_219 : MUX2H
      port map(A => \BNC_CNT[3]_net_1\, B => \BNC_CNT_3[3]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_219\);
    
    \FID_6_r[25]\ : OA21
      port map(A => N_1493_i, B => \FID_6_iv_0_0_0_i[25]\, C => 
        N_532_3_4, Y => \FID_6[25]\);
    
    \FID_6_iv_0_0_0[22]\ : OAI21FTT
      port map(A => \EVNT_NUM[6]_net_1\, B => N_1575_1, C => 
        N_1513, Y => \FID_6_iv_0_0_0_i[22]\);
    
    \CNT_0[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_8_i[0]_net_1\, CLR => 
        CLEAR_0, Q => \CNT_0[0]_net_1\);
    
    un2_bnc_cnt_I_24 : XOR2
      port map(A => N_146, B => \BNC_CNT[5]_net_1\, Y => I_24_1);
    
    un1_CNT_1_I_22 : XOR2
      port map(A => \CNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_22_0);
    
    \STATE1_ns_i_0_a2_0[1]\ : OA21FTT
      port map(A => \READ_PDL_FLAG\, B => \READ_ADC_FLAG\, C => 
        N_1576_1, Y => N_1563_i);
    
    \STATE1_0[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[0]\, CLR => 
        CLEAR_0, Q => \STATE1_0[0]_net_1\);
    
    REG_1_20_127_i_a2 : AO21
      port map(A => N_226_i_0, B => N_701_i_0_0, C => \REG[20]\, 
        Y => \REG_1_20_127_i_a2\);
    
    CRC32_101 : MUX2H
      port map(A => \CRC32[8]_net_1\, B => N_1378, S => N_1469, Y
         => \CRC32_101\);
    
    L1AF2 : DFFC
      port map(CLK => ALICLK_c, D => \L1AF1\, CLR => HWRES_c_12, 
        Q => \L1AF2\);
    
    \un2_i2c_chain_0_0_0_a2_0[0]\ : NOR2
      port map(A => \CNT_0[5]_net_1\, B => \CNT_0[4]_net_1\, Y
         => N_1764);
    
    \FID_6_iv_0_0_a2_1[13]\ : NOR2FT
      port map(A => \EVENT_DWORD[13]_net_1\, B => N_620_4_1, Y
         => N_1531_i);
    
    \BNC_CNT_3[5]\ : AND2
      port map(A => I_24_1, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[5]_net_1\);
    
    EVENT_DWORD_143 : MUX2H
      port map(A => \EVENT_DWORD[5]_net_1\, B => 
        \EVENT_DWORD_17[5]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_143\);
    
    \BNC_CNT[22]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_238\, CLR => 
        CLEAR_3, Q => \BNC_CNT[22]_net_1\);
    
    BNC_CNT_231 : MUX2H
      port map(A => \BNC_CNT[15]_net_1\, B => 
        \BNC_CNT_3[15]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_231\);
    
    \un2_i2c_chain_0_0_0_a2_8[5]\ : AND3
      port map(A => N_1770, B => N_188, C => \CNT[1]_net_1\, Y
         => N_1725_i);
    
    STATE1_1_sqmuxa_1_0_a5_0_o2 : OR2
      port map(A => N_188, B => N_192, Y => N_193);
    
    \CRC32[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_109\, CLR => CLEAR_6, 
        Q => \CRC32[16]_net_1\);
    
    \STATE1_ns_1_iv_0_0_a2_4_1[2]\ : NOR3FFT
      port map(A => PULSE(2), B => REG_i_0(5), C => 
        EVNT_TRG_net_1, Y => \STATE1_ns_1_iv_0_0_a2_4_1[2]_net_1\);
    
    EVNT_NUM_2_I_42 : XOR2
      port map(A => \EVNT_NUM[5]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => \EVNT_NUM_2[5]\);
    
    \EVENT_DWORD_17_i_0_0[24]\ : OAI21TTF
      port map(A => N_105_i_0_0, B => PDL_RDATA(0), C => N_1707, 
        Y => \EVENT_DWORD_17_i_0_0[24]_net_1\);
    
    un2_bnc_cnt_I_69 : AND3
      port map(A => \BNC_CNT[9]_net_1\, B => \BNC_CNT[10]_net_1\, 
        C => \BNC_CNT[11]_net_1\, Y => \DWACT_FINC_E[7]\);
    
    un1_STATE1_1_sqmuxa_1_i_i : OR2
      port map(A => N_1454, B => N_248, Y => N_203);
    
    \EVENT_DWORD_17_i_0_a2[18]\ : NOR2
      port map(A => \EVENT_DWORD[18]_net_1\, B => N_1229_i_1, Y
         => N_1666);
    
    EVENT_DWORD_165 : MUX2H
      port map(A => \EVENT_DWORD[27]_net_1\, B => 
        \EVENT_DWORD_17[27]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_165\);
    
    \CNT_8_i_a3[0]\ : NOR2
      port map(A => N_252, B => N_188, Y => N_1759_i);
    
    N_752_i_i_o2 : OR2FT
      port map(A => \STATE1[1]_net_1\, B => N_221, Y => N_252);
    
    \FID_2_0[7]\ : XOR2
      port map(A => \CRC32[15]_net_1\, B => \CRC32[27]_net_1\, Y
         => \FID_2_0[7]_net_1\);
    
    \CNT_0[2]\ : DFFC
      port map(CLK => CLK_c_c, D => N_78, CLR => CLEAR_0, Q => 
        \CNT_0[2]_net_1\);
    
    \CRC32_2_i_0[8]\ : NOR2FT
      port map(A => N_532_3_1, B => N_282_i_i_0, Y => N_1378);
    
    CRC32_105 : MUX2H
      port map(A => \CRC32[12]_net_1\, B => N_1290, S => N_1469_1, 
        Y => \CRC32_105\);
    
    READ_PDL_FLAG_92_0_0_a2_1 : NOR3FFT
      port map(A => \READ_PDL_FLAG\, B => N_166, C => 
        \STATE1_0[3]_net_1\, Y => N_1671);
    
    FID_186 : MUX2H
      port map(A => \FID[16]_net_1\, B => \FID_6[16]\, S => 
        N_205_1, Y => \FID_186\);
    
    PDL_RADDR_210 : MUX2H
      port map(A => \CNT[0]_net_1\, B => \PDL_RADDR[0]_net_1\, S
         => STATE1_1_sqmuxa_1, Y => \PDL_RADDR_210\);
    
    \FID_6_iv_0_0_a2_1[24]\ : NOR2FT
      port map(A => \EVENT_DWORD[24]_net_1\, B => N_620_4_1, Y
         => N_1490_i);
    
    FID_188 : MUX2H
      port map(A => \FID[18]_net_1\, B => \FID_6[18]\, S => 
        N_205_1, Y => \FID_188\);
    
    BNC_CNT_235 : MUX2H
      port map(A => \BNC_CNT[19]_net_1\, B => 
        \BNC_CNT_3[19]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_235\);
    
    \FID_6_r[13]\ : OA21
      port map(A => N_1531_i, B => \FID_6_iv_0_0_0_i[13]\, C => 
        N_532_3_5, Y => \FID_6[13]\);
    
    \STATE1_ns_1_iv_0_0_o3_4[0]\ : AND3FFT
      port map(A => \STATE1_ns_1_iv_0_0_o3_2_i[0]\, B => 
        \STATE1_ns_1_iv_0_0_o3_1_i[0]\, C => N_1575, Y => 
        \STATE1_ns_1_iv_0_0_o3_4[0]_net_1\);
    
    un2_bnc_cnt_I_146 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \BNC_CNT[21]_net_1\, 
        C => \BNC_CNT[22]_net_1\, Y => \DWACT_FINC_E[33]\);
    
    \REG_1[42]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I10_S, CLR => 
        CLEAR_19, Q => \REG[42]\);
    
    \STATE1_ns_0_0_0_a2_1[3]\ : NOR2FT
      port map(A => N_1733_1, B => N_620_4, Y => N_1733_i);
    
    un1_REG_1_ADD_16x16_slow_I11_S : XOR2
      port map(A => I10_un1_CO1, B => ADD_16x16_slow_I11_S_0, Y
         => ADD_16x16_slow_I11_S);
    
    \REG_1[41]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I9_S, CLR => 
        CLEAR_19, Q => \REG[41]\);
    
    \EVENT_DWORD_17_r[2]\ : AND3FFT
      port map(A => N_1644, B => \EVENT_DWORD_17_i_0_0[2]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[2]\);
    
    \STATE1_ns_1_iv_0_0_o3_0[0]\ : AOI21TTF
      port map(A => N_226_i_0, B => N_1752_1, C => N_1750, Y => 
        \STATE1_ns_1_iv_0_0_o3_0[0]_net_1\);
    
    \CRC32[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_114\, CLR => CLEAR_7, 
        Q => \CRC32[21]_net_1\);
    
    \FID_6_0_iv_0_0_0[0]\ : OAI21FTT
      port map(A => REG_43, B => N_1574_0, C => N_1502, Y => 
        \FID_6_0_iv_0_0_0_i[0]\);
    
    un1_REG_1_G_16_0_o2 : NAND2
      port map(A => ADD_16x16_slow_I8_un1_CO1_0, B => I8_un4_CO1, 
        Y => I8_un1_CO1);
    
    CRC32_97 : MUX2H
      port map(A => \CRC32[4]_net_1\, B => N_1216, S => N_1469, Y
         => \CRC32_97\);
    
    un2_bnc_cnt_I_55 : AND3
      port map(A => \DWACT_FINC_E[4]\, B => \BNC_CNT[8]_net_1\, C
         => \BNC_CNT[9]_net_1\, Y => N_123);
    
    \FID[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_183\, CLR => CLEAR_13, Q
         => \FID[13]_net_1\);
    
    \CNT_8_i_o3[0]\ : OA21FTF
      port map(A => \STATE1_0[2]_net_1\, B => N_1600, C => 
        N_1759_i, Y => N_183);
    
    PDL_RADDR_212 : MUX2H
      port map(A => \CNT[2]_net_1\, B => \PDL_RADDR[2]_net_1\, S
         => STATE1_1_sqmuxa_1, Y => \PDL_RADDR_212\);
    
    un1_EVENT_DWORD_0_sqmuxa_0_0_a2_0_0_a2 : NAND3FTT
      port map(A => N_105_i_0, B => \STATE1[3]_net_1\, C => 
        \PDL_RACK_sync\, Y => N_520);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \un2_i2c_chain_0_0_0_3[4]\ : OAI21FTT
      port map(A => N_1776, B => N_1765, C => 
        \un2_i2c_chain_0_0_0_0[4]_net_1\, Y => 
        \un2_i2c_chain_0_0_0_3_i[4]\);
    
    \STATE2[2]\ : DFFS
      port map(CLK => CLK_c_c, D => \STATE2_ns[0]\, SET => 
        CLEAR_20, Q => \STATE2[2]_net_1\);
    
    FID_201 : MUX2H
      port map(A => \FID[31]_net_1\, B => \FID_6[31]\, S => 
        N_205_0, Y => \FID_201\);
    
    \BNC_CNT_3[3]\ : AND2
      port map(A => I_13_3, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[3]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I1_S_0 : XOR2FT
      port map(A => \REG[33]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I1_S_0);
    
    CYC_STAT_0 : DFFC
      port map(CLK => CLK_c_c, D => \CYC_STAT_0_2\, CLR => 
        HWRES_c_11, Q => \CYC_STAT_0\);
    
    un1_STATE1_11_0_i_a2_0_0_a2 : NAND2
      port map(A => N_1601, B => \STATE1[2]_net_1\, Y => N_1586);
    
    un1_REG_1_ADD_16x16_slow_I10_S : XOR2
      port map(A => N224, B => ADD_16x16_slow_I10_S_0, Y => 
        ADD_16x16_slow_I10_S);
    
    \EVENT_DWORD_17_i_0_0[15]\ : OAI21TTF
      port map(A => \EVENT_DWORD[23]_net_1\, B => N_105_i_0_1, C
         => N_1623, Y => \EVENT_DWORD_17_i_0_0[15]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m14_2 : NOR2
      port map(A => \REG[41]\, B => \REG[42]\, Y => 
        ADD_16x16_slow_I14_un1_CO1_m14_2);
    
    \FID_6_r[19]\ : OA21
      port map(A => N_324_i, B => \FID_6_iv_0_0_i[19]\, C => 
        N_532_3_4, Y => \FID_6[19]\);
    
    \EVENT_DWORD[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_163\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[25]_net_1\);
    
    \STATE1_ns_0_0_0[3]\ : NAND3FFT
      port map(A => N_1733_i, B => \STATE1_ns_0_0_0_2_i[3]\, C
         => STATE1_1_sqmuxa_1, Y => \STATE1_ns[3]\);
    
    \EVENT_DWORD_17_i_0_0[18]\ : OAI21TTF
      port map(A => \EVENT_DWORD[26]_net_1\, B => N_105_i_0_1, C
         => N_1667, Y => \EVENT_DWORD_17_i_0_0[18]_net_1\);
    
    I2C_RREQ_1_sqmuxa_0_a5_0_a2_0 : NOR2
      port map(A => N_1771, B => \STATE1[0]_net_1\, Y => N_1592);
    
    \FID_6_iv_0_0_0[25]\ : OAI21FTT
      port map(A => \EVNT_NUM[9]_net_1\, B => N_1575_1, C => 
        N_1492, Y => \FID_6_iv_0_0_0_i[25]\);
    
    FID_195 : MUX2H
      port map(A => \FID[25]_net_1\, B => \FID_6[25]\, S => 
        N_205_0, Y => \FID_195\);
    
    \un2_i2c_chain_0_0_0_0[6]\ : AO21TTF
      port map(A => N_202_i_i_0, B => N_1638_1, C => N_1640, Y
         => \un2_i2c_chain_0_0_0_0_i[6]\);
    
    L2ASS : DFFC
      port map(CLK => CLK_c_c, D => \REG[334]\, CLR => CLEAR_15, 
        Q => \L2ASS\);
    
    \EVENT_DWORD_17_i_0_a2[24]\ : NOR2
      port map(A => \EVENT_DWORD[24]_net_1\, B => N_1229_i_0, Y
         => N_1706);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m14_3 : OR3FTT
      port map(A => ADD_16x16_slow_I14_un1_CO1_m14_2, B => 
        \REG[44]\, C => \REG[39]\, Y => 
        ADD_16x16_slow_I14_un1_CO1_m14_3_i);
    
    N_1205_i_i_o2 : NOR3
      port map(A => N_1205_i_i_o2_2_i, B => \ORATETMO_i_i[3]\, C
         => \ORATETMO[4]_net_1\, Y => N_226_i_0);
    
    un1_STATE1_18_0_0_a2 : NOR2FT
      port map(A => \STATE1_0[0]_net_1\, B => N_215, Y => 
        N_1673_i);
    
    \BNC_CNT[27]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_243\, CLR => 
        CLEAR_3, Q => \BNC_CNT[27]_net_1\);
    
    un1_REG_1_G_0_o2 : AO21TTF
      port map(A => I12_un1_CO1, B => \REG[45]\, C => 
        ADD_16x16_slow_I13_CO1_0, Y => G_0_o2);
    
    un1_REG_1_ADD_16x16_slow_I5_CO1_1 : AO21
      port map(A => ADD_16x16_slow_I3_CO1_0_a0_1, B => 
        ADD_16x16_slow_I5_CO1_0_a0_3, C => 
        ADD_16x16_slow_I3_CO1_1_0_i_i, Y => 
        ADD_16x16_slow_I5_CO1_0);
    
    \FID_6_0_iv_0_a2_3[0]\ : OR2FT
      port map(A => \EVENT_DWORD[0]_net_1\, B => N_620_4_0, Y => 
        N_1502);
    
    EVENT_DWORD_155 : MUX2H
      port map(A => \EVENT_DWORD[17]_net_1\, B => 
        \EVENT_DWORD_17[17]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_155\);
    
    un1_REG_1_G_5_i_a2 : NAND2
      port map(A => I10_un1_CO1, B => \REG[43]\, Y => I11_un3_CO1);
    
    \CHANNEL[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \CHANNEL_132\, CLR => CLEAR_5, 
        Q => \CHANNEL[2]_net_1\);
    
    STATE1_s6_0_a3_0_a2_0_a2 : OR2
      port map(A => \STATE1_0[0]_net_1\, B => N_215, Y => 
        \STATE1_d[7]\);
    
    \EVENT_DWORD[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_149\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[11]_net_1\);
    
    READ_OR_FLAG_91_i_0_a2 : NOR3
      port map(A => N_258_i_0, B => \STATE1[1]_net_1\, C => 
        \STATE1[3]_net_1\, Y => N_1539);
    
    \PDL_RADDR[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RADDR_210\, CLR => 
        CLEAR_17, Q => \PDL_RADDR[0]_net_1\);
    
    EVNT_NUM_2_I_40 : XOR2
      port map(A => \EVNT_NUM[9]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, Y => \EVNT_NUM_2[9]\);
    
    \FID_6_iv_0_0_0[6]\ : OAI21
      port map(A => N_1575_0, B => \FID_2_i[6]\, C => N_316, Y
         => \FID_6_iv_0_0_0_i[6]\);
    
    \REG_1[46]\ : DFFC
      port map(CLK => CLK_c_c, D => G_0_x2, CLR => CLEAR_19, Q
         => \REG[46]\);
    
    \BNC_CNT[13]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_229\, CLR => 
        CLEAR_2, Q => \BNC_CNT[13]_net_1\);
    
    un4_bnc_res_3 : XOR2
      port map(A => \BNC_CNT[3]_net_1\, B => REG_407, Y => 
        un4_bnc_res_3_i_i);
    
    \RDY_CNT_8_i_0_a2[0]\ : NOR3FTT
      port map(A => \PDL_RACK_sync\, B => N_243, C => N_105_i_0_0, 
        Y => N_1582);
    
    un1_REG_1_G_7_0_o2 : NAND2
      port map(A => ADD_16x16_slow_I11_CO1_0_m5_0, B => 
        I11_un3_CO1, Y => N228);
    
    N_161_i_0_a2 : NOR2FT
      port map(A => \STATE1_0[2]_net_1\, B => N_195, Y => 
        N_161_i_0);
    
    FID_170 : MUX2H
      port map(A => \FID[0]_net_1\, B => \FID_6[0]\, S => N_205, 
        Y => \FID_170\);
    
    un1_CNT_1_I_33 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    \EVENT_DWORD_17_0_a2_0_0_a2[31]\ : NOR2FT
      port map(A => \STATE1_0[3]_net_1\, B => N_105_i_0_0, Y => 
        N_1590);
    
    \EVNT_NUM[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[2]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[2]_net_1\);
    
    \BNC_CNT_3[1]\ : AND2
      port map(A => I_5_2, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[1]_net_1\);
    
    un1_STATE1_17_i_0_i4_0_a2_0_a2_0_i2_0_o2 : OR2
      port map(A => \STATE1_0[2]_net_1\, B => \STATE1_0[1]_net_1\, 
        Y => N_176);
    
    \STATE1_ns_1_iv_0_1_o2_3_o3_0[0]\ : AND2
      port map(A => \PDL_RACK_sync\, B => N_193, Y => N_237);
    
    \CRC32_2_i_0[6]\ : NOR2FT
      port map(A => N_532_3_0, B => N_281_i_i_0, Y => N_1377);
    
    EVENT_DWORD_141 : MUX2H
      port map(A => \EVENT_DWORD[3]_net_1\, B => 
        \EVENT_DWORD_17[3]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_141\);
    
    \EVENT_DWORD_17_i_0_a2[28]\ : NOR2
      port map(A => \EVENT_DWORD[28]_net_1\, B => N_1229_i_0, Y
         => N_1694);
    
    \EVENT_DWORD_17_i_0_0[8]\ : OAI21TTF
      port map(A => \EVENT_DWORD[16]_net_1\, B => N_105_i_0_1, C
         => N_1664, Y => \EVENT_DWORD_17_i_0_0[8]_net_1\);
    
    un2_bnc_cnt_I_34 : AND3
      port map(A => \BNC_CNT[3]_net_1\, B => \BNC_CNT[4]_net_1\, 
        C => \BNC_CNT[5]_net_1\, Y => \DWACT_FINC_E[2]\);
    
    un1_ORATETMO_1_I_17_i_0 : NOR2FT
      port map(A => N_193, B => N_252, Y => N_701_i_0_0);
    
    un4_bnc_res_15 : XOR2
      port map(A => \BNC_CNT[15]_net_1\, B => REG_419, Y => 
        un4_bnc_res_15_i_i);
    
    un1_STATE1_19_i_i : NAND3FTT
      port map(A => N_1587, B => N_522, C => N_253, Y => N_205);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m14_2_0 : OR3
      port map(A => \REG[45]\, B => \REG[46]\, C => \REG[40]\, Y
         => ADD_16x16_slow_I14_un1_CO1_m14_2_0_i);
    
    \FID_6_0_iv_0_a2_0[31]\ : NOR2FT
      port map(A => \EVENT_DWORD[31]_net_1\, B => N_620_4, Y => 
        N_1498_i);
    
    \FID_6_iv_0_0_a2_1[5]\ : NOR2
      port map(A => \EVENT_DWORD[5]_net_1\, B => N_620_4, Y => 
        N_1522);
    
    \FID_6_iv_0_0_a2_1[26]\ : NOR2FT
      port map(A => \EVENT_DWORD[26]_net_1\, B => N_620_4, Y => 
        N_1496_i);
    
    BNC_CNT_218 : MUX2H
      port map(A => \BNC_CNT[2]_net_1\, B => \BNC_CNT_3[2]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_218\);
    
    \FID_6_0_iv_0_0_a2[3]\ : NOR2
      port map(A => GA_c(3), B => N_235, Y => N_309_i);
    
    \un2_i2c_chain_0_i_0_o2_0[2]\ : NAND2
      port map(A => \CNT[2]_net_1\, B => N_1767, Y => N_213);
    
    N_105_i_0_a2_0_a2 : OR2
      port map(A => \STATE1_0[0]_net_1\, B => N_176, Y => 
        N_105_i_0);
    
    \FID_6_iv_0_0_a2_0[24]\ : OR2FT
      port map(A => REG_67, B => N_1574, Y => N_1489);
    
    \un2_i2c_chain_0_i_0_x3[2]\ : XOR2FT
      port map(A => \CNT[0]_net_1\, B => \CNT[1]_net_1\, Y => 
        N_202_i_i_0);
    
    \FID_6_iv_0_0_a2_1[21]\ : NOR2FT
      port map(A => \EVENT_DWORD[21]_net_1\, B => N_620_4_1, Y
         => N_1484_i);
    
    \EVENT_DWORD_17_r[24]\ : AND3FFT
      port map(A => N_1706, B => \EVENT_DWORD_17_i_0_1[24]_net_1\, 
        C => N_532_3_6, Y => \EVENT_DWORD_17[24]\);
    
    \FID_6_iv_0_0_a2_1[9]\ : NOR2
      port map(A => \EVENT_DWORD[9]_net_1\, B => N_620_4, Y => 
        N_1528);
    
    un1_REG_1_ADD_16x16_slow_I2_S : XOR2
      port map(A => N208, B => ADD_16x16_slow_I2_S_0, Y => 
        ADD_16x16_slow_I2_S);
    
    un1_EVENT_DWORD_0_sqmuxa_0_0_o2 : OA21FTF
      port map(A => N_1593, B => N_215, C => N_1454_0, Y => N_234);
    
    \CRC32[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_106\, CLR => CLEAR_6, 
        Q => \CRC32[13]_net_1\);
    
    BNC_CNT_217 : MUX2H
      port map(A => \BNC_CNT[1]_net_1\, B => \BNC_CNT_3[1]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_217\);
    
    FID_181 : MUX2H
      port map(A => \FID[11]_net_1\, B => \FID_6[11]\, S => 
        N_205_1, Y => \FID_181\);
    
    CYC_STAT_89 : MUX2H
      port map(A => CLEAR_PSM_FLAGS_i_0, B => \CYC_STAT\, S => 
        \CYC_STAT_1_sqmuxa\, Y => \CYC_STAT_89\);
    
    BNC_CNT_216 : MUX2H
      port map(A => \BNC_CNT[0]_net_1\, B => \BNC_CNT_3[0]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_216\);
    
    \EVENT_DWORD_17_i_o2_1_o2_1[7]\ : OA21FTF
      port map(A => \STATE1_0[0]_net_1\, B => N_180, C => 
        N_1755_i, Y => N_1229_i_1);
    
    PDL_RADDR_211 : MUX2H
      port map(A => \CNT[1]_net_1\, B => \PDL_RADDR[1]_net_1\, S
         => STATE1_1_sqmuxa_1, Y => \PDL_RADDR_211\);
    
    FID_183 : MUX2H
      port map(A => \FID[13]_net_1\, B => \FID_6[13]\, S => 
        N_205_1, Y => \FID_183\);
    
    BNC_CNT_241 : MUX2H
      port map(A => \BNC_CNT[25]_net_1\, B => 
        \BNC_CNT_3[25]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_241\);
    
    un2_bnc_cnt_I_98 : XOR2
      port map(A => N_93_0, B => \BNC_CNT[16]_net_1\, Y => I_98);
    
    un4_bnc_res_12 : XOR2
      port map(A => \BNC_CNT[12]_net_1\, B => REG_416, Y => 
        un4_bnc_res_12_i_i);
    
    \CRC32_2_i_0[9]\ : NOR2FT
      port map(A => N_532_3_1, B => N_283_i_i_0, Y => N_1379);
    
    \CRC32_2_i_0_x2[5]\ : XOR2FT
      port map(A => \CRC32[5]_net_1\, B => \EVENT_DWORD[5]_net_1\, 
        Y => N_280_i_i_0);
    
    \FID_6_iv_0_0_a2_1[15]\ : NOR2FT
      port map(A => \EVENT_DWORD[15]_net_1\, B => N_620_4_1, Y
         => N_1478_i);
    
    EVNT_TRG_1_f0_i_0 : OA21TTF
      port map(A => EVNT_TRG_net_1, B => \STATE2[1]_net_1\, C => 
        \STATE2[0]_net_1\, Y => N_1147);
    
    \EVNT_NUM[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[6]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[6]_net_1\);
    
    \un2_i2c_chain_0_0_0_a3[1]\ : OR2FT
      port map(A => \CNT[3]_net_1\, B => \CNT_0[2]_net_1\, Y => 
        N_1769);
    
    READ_ADC_FLAG : DFFC
      port map(CLK => CLK_c_c, D => \READ_ADC_FLAG_90_0_0\, CLR
         => CLEAR_17, Q => \READ_ADC_FLAG\);
    
    \FID_6_0_iv_0_a2_1[2]\ : OR2FT
      port map(A => \EVENT_DWORD[2]_net_1\, B => N_620_4_0, Y => 
        N_1519);
    
    \EVENT_DWORD_17_i_0_a2[16]\ : NOR2
      port map(A => \EVENT_DWORD[16]_net_1\, B => N_1229_i_1, Y
         => N_1660);
    
    \EVENT_DWORD_17_i_0_1[20]\ : OAI21FTF
      port map(A => N_1454_0, B => OR_RDATA(0), C => 
        \EVENT_DWORD_17_i_0_0[20]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[20]_net_1\);
    
    \CRC32_2_i[19]\ : NOR2FT
      port map(A => N_532_3_1, B => N_273_i_i_0, Y => N_1468);
    
    \un2_i2c_chain_0_0_0_a2_0_1[6]\ : NOR2
      port map(A => N_1763, B => N_1769, Y => N_1638_1);
    
    un1_STATE1_2_0_i_a3_i : NAND2
      port map(A => N_532_3, B => N_620_4, Y => N_1469);
    
    BNC_CNT_245 : MUX2H
      port map(A => \BNC_CNT[29]_net_1\, B => 
        \BNC_CNT_3[29]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_245\);
    
    un4_bnc_res_25 : XOR2
      port map(A => \BNC_CNT[25]_net_1\, B => REG_429, Y => 
        un4_bnc_res_25_i_i);
    
    \FID_2_0[11]\ : XOR2
      port map(A => \CRC32[19]_net_1\, B => \CRC32[31]_net_1\, Y
         => \FID_2_0[11]_net_1\);
    
    \BNC_CNT_3[24]\ : AND2
      port map(A => I_166, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[24]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I1_un3_CO1_0 : AND2
      port map(A => \REG[32]\, B => \REG[33]\, Y => 
        ADD_16x16_slow_I1_un3_CO1_0);
    
    \STATE1_ns_i_0_a2_6[1]\ : NOR3FFT
      port map(A => EVNT_TRG_net_1, B => REG_i_0(5), C => 
        N_532_3_3, Y => N_1569_i);
    
    EVENT_DWORD_147 : MUX2H
      port map(A => \EVENT_DWORD[9]_net_1\, B => 
        \EVENT_DWORD_17[9]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_147\);
    
    un4_bnc_res_NE_0 : OR3
      port map(A => un4_bnc_res_NE_29_i, B => un4_bnc_res_NE_25_i, 
        C => un4_bnc_res_NE_24_i, Y => un4_bnc_res_i_0);
    
    \un2_i2c_chain_0_0_0_a2_1[6]\ : NOR3FFT
      port map(A => N_199, B => N_1770, C => \CNT_0[1]_net_1\, Y
         => N_1639_i);
    
    un1_STATE1_11_0_i_a2 : NOR2FT
      port map(A => \STATE1_0[0]_net_1\, B => N_176, Y => 
        N_1541_i);
    
    un1_REG_1_ADD_16x16_slow_I11_CO1_0_m5_0_a4_0 : OR3
      port map(A => ADD_16x16_slow_I11_CO1_0tt_m3_0_a2, B => 
        I6_un4_CO1, C => ADD_16x16_slow_I11_CO1_0_m5_0_a4_0_0, Y
         => ADD_16x16_slow_I11_CO1_0_m5_0_a4_0);
    
    \BNC_CNT_3[0]\ : NOR2FT
      port map(A => un4_bnc_res_i_0, B => \BNC_CNT[0]_net_1\, Y
         => \BNC_CNT_3[0]_net_1\);
    
    un1_ORATETMO_1_I_11 : XOR2
      port map(A => \ORATETMO[2]_net_1\, B => N_701_i_0_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_1[0]\);
    
    \CNT_8_i[3]\ : AND2
      port map(A => N_185_i, B => I_23, Y => N_81);
    
    \BNC_CNT[24]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_240\, CLR => 
        CLEAR_3, Q => \BNC_CNT[24]_net_1\);
    
    STATE1_tr16_1_0_a2_0_a2_0_a2_0_a2_1 : OR2FT
      port map(A => N_1573, B => N_221, Y => N_620_4_1);
    
    \EVENT_DWORD_17_i_0_0[26]\ : OAI21TTF
      port map(A => N_105_i_0_0, B => PDL_RDATA(2), C => N_1699, 
        Y => \EVENT_DWORD_17_i_0_0[26]_net_1\);
    
    un4_bnc_res_7 : XOR2
      port map(A => \BNC_CNT[7]_net_1\, B => REG_411, Y => 
        un4_bnc_res_7_i_i);
    
    \EVENT_DWORD_17_i_0_0[17]\ : OAI21TTF
      port map(A => \EVENT_DWORD[25]_net_1\, B => N_105_i_0_1, C
         => N_291, Y => \EVENT_DWORD_17_i_0_0[17]_net_1\);
    
    CRC32_113 : MUX2H
      port map(A => \CRC32[20]_net_1\, B => N_1383, S => N_1469_1, 
        Y => \CRC32_113\);
    
    CRC32_117 : MUX2H
      port map(A => \CRC32[24]_net_1\, B => N_1293, S => N_1469_0, 
        Y => \CRC32_117\);
    
    un1_REG_1_ADD_16x16_slow_I3_CO1 : AO21TTF
      port map(A => I2_un1_CO1, B => \REG[35]\, C => 
        ADD_16x16_slow_I3_CO1_0, Y => N212);
    
    CRC32_93 : MUX2H
      port map(A => \CRC32[0]_net_1\, B => N_1287, S => N_1469, Y
         => \CRC32_93\);
    
    \FID_6_r[21]\ : OA21
      port map(A => N_1484_i, B => \FID_6_iv_0_0_0_i[21]\, C => 
        N_532_3_4, Y => \FID_6[21]\);
    
    \FID_2_0[4]\ : XOR2
      port map(A => \CRC32[12]_net_1\, B => \CRC32[24]_net_1\, Y
         => \FID_2_0[4]_net_1\);
    
    \EVENT_DWORD_17_i_0_0[11]\ : OAI21TTF
      port map(A => \EVENT_DWORD[19]_net_1\, B => N_105_i_0_1, C
         => N_335, Y => \EVENT_DWORD_17_i_0_0[11]_net_1\);
    
    CRC32_123 : MUX2H
      port map(A => \CRC32[30]_net_1\, B => N_1294, S => N_1469_0, 
        Y => \CRC32_123\);
    
    un5_evread_7_0 : OR3FTT
      port map(A => \un5_evread_4\, B => \REG[45]\, C => 
        \REG[38]\, Y => un5_evread_7_0_i);
    
    un4_bnc_res_22 : XOR2
      port map(A => \BNC_CNT[22]_net_1\, B => REG_426, Y => 
        un4_bnc_res_22_i_i);
    
    \EVNT_NUM[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[7]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[7]_net_1\);
    
    \STATE1_ns_1_iv_0_o2_0[0]\ : NOR2
      port map(A => EVNT_TRG_net_1, B => REG_0, Y => N_1183_i);
    
    OR_RADDR_209 : MUX2H
      port map(A => \OR_RADDR[5]_net_1\, B => N_679, S => N_248, 
        Y => \OR_RADDR_209\);
    
    \FID_6_iv_0_0_0[21]\ : OAI21FTT
      port map(A => \EVNT_NUM[5]_net_1\, B => N_1575_1, C => 
        N_1483, Y => \FID_6_iv_0_0_0_i[21]\);
    
    \FID_6_r[27]\ : OA21
      port map(A => N_1544_i, B => \FID_6_iv_0_0_i[27]\, C => 
        N_532_3_4, Y => \FID_6[27]\);
    
    \un2_i2c_chain_0_0_0_a2_1[0]\ : AND2
      port map(A => \CNT[5]_net_1\, B => \CNT_0[3]_net_1\, Y => 
        N_1773);
    
    \FID[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_187\, CLR => CLEAR_13, Q
         => \FID[17]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I12_un1_CO1_0_tz_0 : NOR2FT
      port map(A => ADD_16x16_slow_I11_CO1_0_m5_0, B => \REG[44]\, 
        Y => ADD_16x16_slow_I12_un1_CO1_0_tz_0);
    
    un1_ORATETMO_1_I_25 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_5[0]\);
    
    L2RF3 : DFFC
      port map(CLK => ALICLK_c, D => \L2RF2\, CLR => HWRES_c_12, 
        Q => \L2RF3\);
    
    \STATE1[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns_i_0[1]_net_1\, CLR
         => CLEAR_19, Q => \STATE1[1]_net_1\);
    
    L2RF1 : DFFC
      port map(CLK => ALICLK_c, D => L2R_c_c, CLR => HWRES_c_12, 
        Q => \L2RF1\);
    
    un2_bnc_cnt_I_155 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[33]\, Y => N_52);
    
    \FID_2[9]\ : XOR2
      port map(A => \CRC32[5]_net_1\, B => \FID_2_0[9]_net_1\, Y
         => \FID_2[9]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2_0[23]\ : NOR2
      port map(A => I2C_RDATA(3), B => N_1768_i, Y => N_1715);
    
    un1_CNT_1_I_15 : XOR2
      port map(A => \CNT[0]_net_1\, B => 
        \un1_EVENT_DWORD_0_sqmuxa_0_0\, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \EVENT_DWORD_17_r[18]\ : AND3FFT
      port map(A => N_1666, B => \EVENT_DWORD_17_i_0_0[18]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[18]\);
    
    un1_REG_1_ADD_16x16_slow_I13_CO1_0_a0_2 : OR2
      port map(A => \REG[40]\, B => \REG[41]\, Y => 
        ADD_16x16_slow_I13_CO1_0_a0_2_i);
    
    PDL_RADDR_215 : MUX2H
      port map(A => \CNT[5]_net_1\, B => \PDL_RADDR[5]_net_1\, S
         => STATE1_1_sqmuxa_1, Y => \PDL_RADDR_215\);
    
    \STATE1[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[0]\, CLR => 
        CLEAR_19, Q => \STATE1[0]_net_1\);
    
    \CNT_0[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_8_i[5]_net_1\, CLR => 
        CLEAR_0, Q => \CNT_0[5]_net_1\);
    
    \FID_6_iv_0_0_a2_0[26]\ : OR2FT
      port map(A => REG_69, B => N_1574, Y => N_1495);
    
    \FID_6_r[8]\ : AND3FFT
      port map(A => N_1525, B => \FID_6_iv_0_0_0[8]_net_1\, C => 
        N_532_3_5, Y => \FID_6[8]\);
    
    \FID_6_0_iv_0_0_a2[0]\ : NOR2
      port map(A => GA_c(0), B => N_235, Y => N_1500_i);
    
    un4_bnc_res_10 : XOR2
      port map(A => \BNC_CNT[10]_net_1\, B => REG_414, Y => 
        un4_bnc_res_10_i_i);
    
    \EVENT_DWORD_17_r[4]\ : AND3FFT
      port map(A => N_326, B => \EVENT_DWORD_17_i_0_0[4]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[4]\);
    
    un2_bnc_cnt_I_51 : AND2
      port map(A => \BNC_CNT[8]_net_1\, B => \DWACT_FINC_E[4]\, Y
         => N_126);
    
    FID_192 : MUX2H
      port map(A => \FID[22]_net_1\, B => \FID_6[22]\, S => 
        N_205_0, Y => \FID_192\);
    
    un2_bnc_cnt_I_56 : XOR2
      port map(A => N_123, B => \BNC_CNT[10]_net_1\, Y => I_56_0);
    
    \FID_6_iv_0_0_a2_0[21]\ : OR2FT
      port map(A => REG_64, B => N_1574_1, Y => N_1483);
    
    un1_REG_1_G_15_0_a2 : AND2
      port map(A => I6_un1_CO1_i_0_i, B => \REG[39]\, Y => 
        I7_un3_CO1);
    
    \EVENT_DWORD_17_i_0_o2_i[3]\ : OAI21FTT
      port map(A => N_120_i, B => N_176, C => I2C_RACK, Y => 
        N_1768_i);
    
    BNC_CNT_224 : MUX2H
      port map(A => \BNC_CNT[8]_net_1\, B => \BNC_CNT_3[8]_net_1\, 
        S => LBSP_c_1(2), Y => \BNC_CNT_224\);
    
    \EVENT_DWORD_17_i_o2_1_o2[7]\ : OA21FTF
      port map(A => \STATE1_0[0]_net_1\, B => N_180, C => 
        N_1755_i, Y => N_1229_i);
    
    un2_bnc_cnt_I_52 : XOR2
      port map(A => N_126, B => \BNC_CNT[9]_net_1\, Y => I_52_0);
    
    un1_STATE1_5_0_0_0 : OR2FT
      port map(A => N_532_3_0, B => N_161_i_0, Y => un1_STATE1_5);
    
    \BNC_CNT[5]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_221\, CLR => 
        CLEAR_4, Q => \BNC_CNT[5]_net_1\);
    
    \ORATETMO_7_0_0[0]\ : OR2
      port map(A => N_233, B => \DWACT_ADD_CI_0_partial_sum_1[0]\, 
        Y => \ORATETMO_7[0]\);
    
    \CRC32_2_i[29]\ : NOR2FT
      port map(A => N_532_3_2, B => N_248_i_i_0, Y => N_1594);
    
    un2_bnc_cnt_I_189 : AND3
      port map(A => \BNC_CNT[24]_net_1\, B => \BNC_CNT[25]_net_1\, 
        C => \BNC_CNT[26]_net_1\, Y => \DWACT_FINC_E[22]\);
    
    un1_REG_1_ADD_16x16_slow_I13_CO1_0_a0_3 : OR3FTT
      port map(A => ADD_16x16_slow_I13_CO1_0_a0_0, B => \REG[43]\, 
        C => \REG[42]\, Y => ADD_16x16_slow_I13_CO1_0_a0_3_i);
    
    \EVENT_DWORD_17_r[26]\ : AND3FFT
      port map(A => N_1698, B => \EVENT_DWORD_17_i_0_1[26]_net_1\, 
        C => N_532_3_6, Y => \EVENT_DWORD_17[26]\);
    
    un2_bnc_cnt_I_152 : AND3
      port map(A => \DWACT_FINC_E[34]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[5]\, Y => \DWACT_FINC_E[29]\);
    
    un1_STATE1_17_i_0_i4_0_a2_0_a2_0_i2_0_o2_i : INV
      port map(A => \STATE1[2]_net_1\, Y => \STATE1_i_0[2]\);
    
    N_105_i_0_a2_0_a2_0 : OR2
      port map(A => \STATE1_0[0]_net_1\, B => N_176, Y => 
        N_105_i_0_0);
    
    \CRC32[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_119\, CLR => CLEAR_7, 
        Q => \CRC32[26]_net_1\);
    
    EVNT_NUM_2_I_32 : XOR2
      port map(A => \EVNT_NUM[0]_net_1\, B => N_161_i_0, Y => 
        \DWACT_ADD_CI_0_partial_sum_2[0]\);
    
    \EVENT_DWORD_17_r[27]\ : AND3FFT
      port map(A => N_1679, B => \EVENT_DWORD_17_i_1[27]_net_1\, 
        C => N_532_3_6, Y => \EVENT_DWORD_17[27]\);
    
    \EVENT_DWORD_17_i_0_a2[26]\ : NOR2
      port map(A => \EVENT_DWORD[26]_net_1\, B => N_1229_i_0, Y
         => N_1698);
    
    \FID_6_iv_0_a2_0[19]\ : OR2FT
      port map(A => REG_62, B => N_1574_1, Y => N_323);
    
    \CRC32[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_93\, CLR => CLEAR_6, Q
         => \CRC32[0]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2_0[13]\ : NOR2
      port map(A => \EVENT_DWORD[13]_net_1\, B => N_1229_i_1, Y
         => N_339);
    
    CHIP_ADDR_133 : MUX2H
      port map(A => \CHIP_ADDR[0]_net_1\, B => N_94, S => 
        I2C_RREQ_1_sqmuxa, Y => \CHIP_ADDR_133\);
    
    un1_REG_1_ADD_16x16_slow_I5_CO1_0_a0_2 : NOR2
      port map(A => \REG[32]\, B => \REG[33]\, Y => 
        ADD_16x16_slow_I3_CO1_0_a0_1);
    
    \EVENT_DWORD_17_i_1[29]\ : OAI21FTF
      port map(A => N_1454, B => OR_RDATA(9), C => 
        \EVENT_DWORD_17_i_0[29]_net_1\, Y => 
        \EVENT_DWORD_17_i_1[29]_net_1\);
    
    \EVENT_DWORD_17_r[7]\ : AND3FFT
      port map(A => N_1621, B => \EVENT_DWORD_17_i_0_0[7]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[7]\);
    
    \EVENT_DWORD_17_i_0[29]\ : OAI21TTF
      port map(A => N_105_i_0_0, B => PDL_RDATA(5), C => N_1682, 
        Y => \EVENT_DWORD_17_i_0[29]_net_1\);
    
    CRC32_103 : MUX2H
      port map(A => \CRC32[10]_net_1\, B => N_1289, S => N_1469_1, 
        Y => \CRC32_103\);
    
    CRC32_107 : MUX2H
      port map(A => \CRC32[14]_net_1\, B => N_1291, S => N_1469_1, 
        Y => \CRC32_107\);
    
    un2_bnc_cnt_I_44 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => N_131);
    
    un1_STATE1_18_0_0_1 : NAND3FTT
      port map(A => N_1673_i, B => N_1672, C => N_1762, Y => 
        un1_STATE1_18_1);
    
    \REG_1[33]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I1_S, CLR => 
        CLEAR_18, Q => \REG[33]\);
    
    \STATE2_ns_a3_0_a2_0_a2[0]\ : NOR2
      port map(A => \STATE2[1]_net_1\, B => \TRIGGER_sync\, Y => 
        \STATE2_ns[0]\);
    
    \CRC32_2_i_0[2]\ : NOR2FT
      port map(A => N_532_3_0, B => N_261_i_i_0, Y => N_1375);
    
    OR_RADDR_204 : MUX2H
      port map(A => \OR_RADDR[0]_net_1\, B => N_689, S => N_248, 
        Y => \OR_RADDR_204\);
    
    \EVENT_DWORD_17_i_0_a2_0[5]\ : NOR2
      port map(A => \EVENT_DWORD[5]_net_1\, B => N_1229_i, Y => 
        N_333);
    
    \EVENT_DWORD_17_i_0_a2_0[22]\ : NOR2
      port map(A => I2C_RDATA(2), B => N_1768_i, Y => N_1711);
    
    \FID_6_iv_0_0_a2_1[23]\ : NOR2FT
      port map(A => \EVENT_DWORD[23]_net_1\, B => N_620_4_1, Y
         => N_1487_i);
    
    \EVENT_DWORD_17_i_0_a2[0]\ : NOR2
      port map(A => \EVENT_DWORD[0]_net_1\, B => N_1229_i, Y => 
        N_1641);
    
    un2_bnc_cnt_I_203 : XOR2
      port map(A => N_19_0, B => \BNC_CNT[28]_net_1\, Y => I_203);
    
    \FID_6_iv_0_a2_1[27]\ : NOR2FT
      port map(A => \EVENT_DWORD[27]_net_1\, B => N_620_4, Y => 
        N_1544_i);
    
    un4_bnc_res_NE : OR3
      port map(A => un4_bnc_res_NE_29_i, B => un4_bnc_res_NE_25_i, 
        C => un4_bnc_res_NE_24_i, Y => un4_bnc_res_i);
    
    BNC_CNT_233 : MUX2H
      port map(A => \BNC_CNT[17]_net_1\, B => 
        \BNC_CNT_3[17]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_233\);
    
    un4_bnc_res_20 : XOR2
      port map(A => \BNC_CNT[20]_net_1\, B => REG_424, Y => 
        un4_bnc_res_20_i_i);
    
    un1_REG_1_ADD_16x16_slow_I11_CO1_0_m5_0_a4_0_1 : OR2
      port map(A => ADD_16x16_slow_I6_un1_CO1_0, B => \REG[43]\, 
        Y => ADD_16x16_slow_I11_CO1_0_m5_0_a4_0_0);
    
    \STATE1_ns_1_iv_0_0_a2_3_1[2]\ : NOR3FFT
      port map(A => \OR_RACK_sync\, B => \STATE1_i_0[2]\, C => 
        N_222, Y => \STATE1_ns_1_iv_0_0_a2_3_1[2]_net_1\);
    
    EVENT_DWORD_168 : MUX2H
      port map(A => \EVENT_DWORD[30]_net_1\, B => 
        \EVENT_DWORD_17[30]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_168\);
    
    CRC32_112 : MUX2H
      port map(A => \CRC32[19]_net_1\, B => N_1468, S => N_1469_1, 
        Y => \CRC32_112\);
    
    \CHANNEL[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \CHANNEL_130\, CLR => CLEAR_5, 
        Q => \CHANNEL[0]_net_1\);
    
    un1_ORATETMO_1_I_20 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, Y => I_20_2);
    
    CRC32_122 : MUX2H
      port map(A => \CRC32[29]_net_1\, B => N_1594, S => N_1469_0, 
        Y => \CRC32_122\);
    
    \un2_i2c_chain_0_0_0_a2_1_0[3]\ : NOR2FT
      port map(A => \CNT_0[0]_net_1\, B => N_1775, Y => 
        \un2_i2c_chain_0_0_0_a2_1_0[3]_net_1\);
    
    \BNC_CNT_3[14]\ : AND2
      port map(A => I_84_0, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[14]_net_1\);
    
    un1_STATE1_1_sqmuxa_0_0_a2 : OR2
      port map(A => N_105_i_0, B => N_207, Y => N_1672);
    
    \CRC32[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_112\, CLR => CLEAR_7, 
        Q => \CRC32[19]_net_1\);
    
    \EVENT_DWORD_17_i_a2[9]\ : NOR2
      port map(A => \EVENT_DWORD[19]_net_1\, B => N_190_i, Y => 
        N_294);
    
    un4_bnc_res_NE_27 : OR3
      port map(A => un4_bnc_res_NE_20_i, B => un4_bnc_res_NE_14_i, 
        C => un4_bnc_res_NE_15_i, Y => un4_bnc_res_NE_27_i);
    
    CYC_STAT_1 : DFFC
      port map(CLK => CLK_c_c, D => \CYC_STAT_1_2\, CLR => 
        HWRES_c_11, Q => \CYC_STAT_1\);
    
    \BNC_CNT[20]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_236\, CLR => 
        CLEAR_3, Q => \BNC_CNT[20]_net_1\);
    
    \EVENT_DWORD_17_i_0_0[25]\ : OAI21TTF
      port map(A => N_105_i_0_0, B => PDL_RDATA(1), C => N_1736, 
        Y => \EVENT_DWORD_17_i_0_0[25]_net_1\);
    
    un1_CNT_1_I_34 : AND2
      port map(A => \CNT[2]_net_1\, B => \CNT[3]_net_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    \EVENT_DWORD_17_r[15]\ : AND3FFT
      port map(A => N_1624, B => \EVENT_DWORD_17_i_0_0[15]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[15]\);
    
    \CRC32_2_i_0_x2[6]\ : XOR2FT
      port map(A => \CRC32[6]_net_1\, B => \EVENT_DWORD[6]_net_1\, 
        Y => N_281_i_i_0);
    
    un1_REG_1_G_26_0_o2 : AND2
      port map(A => ADD_16x16_slow_I2_un1_CO1_0_a0_0, B => 
        ADD_16x16_slow_I6_un1_CO1_0_a0_2, Y => N_43);
    
    un1_REG_1_ADD_16x16_slow_I4_S_0 : XOR2FT
      port map(A => \REG[36]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I4_S_0);
    
    \EVENT_DWORD_17_i_0_0[28]\ : OAI21TTF
      port map(A => N_105_i_0_0, B => PDL_RDATA(4), C => N_1695, 
        Y => \EVENT_DWORD_17_i_0_0[28]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I7_S_0 : XOR2FT
      port map(A => \REG[39]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I7_S_0);
    
    \FID_6_iv_0_0_0[8]\ : OAI21TTF
      port map(A => N_1574, B => REG_51, C => N_1523, Y => 
        \FID_6_iv_0_0_0[8]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I11_CO1_0_m5_0_a4 : OR3
      port map(A => ADD_16x16_slow_I11_CO1_0tt_m3_0_a2, B => 
        \REG[39]\, C => \REG[43]\, Y => 
        ADD_16x16_slow_I11_CO1_0_m5_0_a4);
    
    un4_bnc_res_NE_14 : OR3
      port map(A => un4_bnc_res_2_i_i, B => un4_bnc_res_14_i_i, C
         => un4_bnc_res_17_i_i, Y => un4_bnc_res_NE_14_i);
    
    \CRC32_2_0_a3_i_x2[7]\ : XOR2FT
      port map(A => \CRC32[7]_net_1\, B => \EVENT_DWORD[7]_net_1\, 
        Y => N_249_i_i_0);
    
    CRC32_95 : MUX2H
      port map(A => \CRC32[2]_net_1\, B => N_1375, S => N_1469, Y
         => \CRC32_95\);
    
    \EVENT_DWORD_17_i_0_a2_0[12]\ : NOR2
      port map(A => \EVENT_DWORD[22]_net_1\, B => N_190_i_0, Y
         => N_1655);
    
    STATE1_1_sqmuxa_1_0_a5_0_a2 : OR3FFT
      port map(A => N_193, B => N_1195_1, C => \PDL_RACK_sync\, Y
         => STATE1_1_sqmuxa_1);
    
    un1_CNT_1_I_26 : XOR2
      port map(A => \CNT[5]_net_1\, B => I_30, Y => I_26);
    
    \STATE1_ns_0_0_0_2[3]\ : NAND3FTT
      port map(A => \STATE1_ns_0_0_0_0_i[3]\, B => N_1734, C => 
        \STATE1_ns_0_0_0_i_0[3]_net_1\, Y => 
        \STATE1_ns_0_0_0_2_i[3]\);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m14 : NOR3
      port map(A => I6_un1_CO1_i_0_i, B => 
        ADD_16x16_slow_I14_un1_CO1_m14_3_i, C => 
        ADD_16x16_slow_I14_un1_CO1_m14_2_0_i, Y => 
        ADD_16x16_slow_I14_un1_CO1_N_18);
    
    PDL_RACK_sync : DFFC
      port map(CLK => CLK_c_c, D => PDL_RACK, CLR => CLEAR_17, Q
         => \PDL_RACK_sync\);
    
    \EVENT_DWORD_17_r[1]\ : AND3FFT
      port map(A => N_330, B => \EVENT_DWORD_17_i_0_0[1]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[1]\);
    
    CRC32_94 : MUX2H
      port map(A => \CRC32[1]_net_1\, B => N_1288, S => N_1469, Y
         => \CRC32_94\);
    
    \EVENT_DWORD_17_0_a2[31]\ : AND2
      port map(A => N_1590, B => PDL_RDATA(7), Y => 
        \EVENT_DWORD_17[31]\);
    
    \REG_1[34]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I2_S, CLR => 
        CLEAR_18, Q => \REG[34]\);
    
    \BNC_CNT_3[9]\ : AND2
      port map(A => I_52_0, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[9]_net_1\);
    
    un2_bnc_cnt_I_105 : XOR2
      port map(A => N_88, B => \BNC_CNT[17]_net_1\, Y => I_105);
    
    un2_bnc_cnt_I_213 : AND3
      port map(A => \BNC_CNT[27]_net_1\, B => \BNC_CNT[28]_net_1\, 
        C => \BNC_CNT[29]_net_1\, Y => \DWACT_FINC_E[26]\);
    
    \FID_6_r[7]\ : OA21
      port map(A => N_320_i, B => \FID_6_iv_0_0_0_i[7]\, C => 
        N_532_3_5, Y => \FID_6[7]\);
    
    \un2_i2c_chain_0_0_0[4]\ : OR3
      port map(A => \un2_i2c_chain_0_0_0_3_i[4]\, B => 
        \un2_i2c_chain_0_0_0_2_i[4]\, C => 
        \un2_i2c_chain_0_0_0_1_i[4]\, Y => N_97);
    
    EVNT_NUM_2_I_50 : XOR2
      port map(A => \EVNT_NUM[4]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\, Y => \EVNT_NUM_2[4]\);
    
    un1_REG_1_ADD_16x16_slow_I7_CO1_1 : OA21TTF
      port map(A => ADD_16x16_slow_I7_CO1_0_a0_2_i, B => 
        ADD_16x16_slow_I7_CO1_0_a0_3_i, C => 
        ADD_16x16_slow_I3_CO1_1_0_i_i, Y => 
        ADD_16x16_slow_I7_CO1_0);
    
    \STATE1_ns_1_iv_0_0_o3_1[0]\ : OAI21TTF
      port map(A => N_120_i, B => N_1613, C => N_7200_i, Y => 
        \STATE1_ns_1_iv_0_0_o3_1_i[0]\);
    
    \FID_6_iv_0_0_a2_1_0_a2_0[28]\ : OR2FT
      port map(A => \STATE1_0[1]_net_1\, B => N_195, Y => 
        N_1575_0);
    
    \BNC_CNT_3[29]\ : AND2
      port map(A => I_210, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[29]_net_1\);
    
    un2_bnc_cnt_I_223 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \DWACT_FINC_E[27]\, Y => N_4);
    
    \FID_6_r[18]\ : OA21
      port map(A => N_1550_i, B => \FID_6_iv_0_0_1_i[18]\, C => 
        N_532_3_4, Y => \FID_6[18]\);
    
    \FID_6_iv_0_0_0[13]\ : OAI21
      port map(A => N_1575_0, B => N_269_i_0_i, C => N_1530, Y
         => \FID_6_iv_0_0_0_i[13]\);
    
    \EVENT_DWORD[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_161\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[23]_net_1\);
    
    \STATE1_ns_1_iv_0_1_o2_3_a3_1[0]\ : AND2
      port map(A => N_1758_1, B => N_1771, Y => N_1746);
    
    \un2_i2c_chain_0_0_0_a2_2[3]\ : NAND3
      port map(A => N_312_1, B => \CNT[0]_net_1\, C => 
        \CNT[1]_net_1\, Y => N_312);
    
    un1_REG_1_ADD_16x16_slow_I12_un1_CO1_0 : AO21
      port map(A => ADD_16x16_slow_I12_un1_CO1_0_tz_0, B => 
        I11_un3_CO1, C => \un2_evread_1[14]\, Y => 
        ADD_16x16_slow_I12_un1_CO1_0);
    
    \FID[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_185\, CLR => CLEAR_13, Q
         => \FID[15]_net_1\);
    
    \CRC32[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_94\, CLR => CLEAR_7, Q
         => \CRC32[1]_net_1\);
    
    EVENT_DWORD_158 : MUX2H
      port map(A => \EVENT_DWORD[20]_net_1\, B => 
        \EVENT_DWORD_17[20]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_158\);
    
    READ_ADC_FLAG_90_0_0 : AO21FTF
      port map(A => N_288_i, B => \READ_ADC_FLAG\, C => 
        \STATE1_d[7]\, Y => \READ_ADC_FLAG_90_0_0\);
    
    \EVENT_DWORD_17_i_0_0[0]\ : OAI21TTF
      port map(A => \EVENT_DWORD[8]_net_1\, B => N_105_i_0, C => 
        N_1642, Y => \EVENT_DWORD_17_i_0_0[0]_net_1\);
    
    un2_bnc_cnt_I_210 : XOR2
      port map(A => N_14, B => \BNC_CNT[29]_net_1\, Y => I_210);
    
    un2_bnc_cnt_I_186 : XOR2
      port map(A => N_31, B => \BNC_CNT[26]_net_1\, Y => I_186);
    
    \BNC_CNT_3[26]\ : AND2
      port map(A => I_186, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[26]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I4_un1_CO1 : AO21TTF
      port map(A => N212, B => \REG[36]\, C => 
        ADD_16x16_slow_I4_un1_CO1_0, Y => I4_un1_CO1);
    
    un1_ORATETMO_1_I_27 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_1_4[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\);
    
    \FID_6_iv_0_0_a2_0[6]\ : OR2FT
      port map(A => REG_49, B => N_1574_0, Y => N_316);
    
    \FID[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_181\, CLR => CLEAR_13, Q
         => \FID[11]_net_1\);
    
    un1_ORATETMO_1_I_16 : XOR2
      port map(A => \ORATETMO_i_i[1]\, B => N_701_i_0, Y => 
        \DWACT_ADD_CI_0_partial_sum[1]\);
    
    L1AF3 : DFFC
      port map(CLK => ALICLK_c, D => \L1AF2\, CLR => HWRES_c_12, 
        Q => \L1AF3\);
    
    CRC32_102 : MUX2H
      port map(A => \CRC32[9]_net_1\, B => N_1379, S => N_1469, Y
         => \CRC32_102\);
    
    \EVENT_DWORD[29]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_167\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[29]_net_1\);
    
    \un2_evread[15]\ : OA21FTT
      port map(A => \FIFO_END_EVNT\, B => EVREAD, C => 
        \un2_evread_0[14]\, Y => \un2_evread[15]_net_1\);
    
    \CRC32_2_i_0_a2_4[17]\ : OR2FT
      port map(A => N_1585_0, B => N_176_0, Y => N_532_3_4);
    
    un2_bnc_cnt_I_220 : AND2
      port map(A => \DWACT_FINC_E[26]\, B => \BNC_CNT[30]_net_1\, 
        Y => \DWACT_FINC_E[27]\);
    
    \FID_6_iv_0_0_0[7]\ : OAI21
      port map(A => N_1575_0, B => \FID_2_i[7]\, C => N_319, Y
         => \FID_6_iv_0_0_0_i[7]\);
    
    \OR_RADDR_3_i_0[0]\ : AND2
      port map(A => N_532_3_3, B => \CNT_0[0]_net_1\, Y => N_689);
    
    un1_REG_1_G_10_0_a2 : NOR3
      port map(A => ADD_16x16_slow_I2_un1_CO1_0_a0_0, B => 
        \FIFO_END_EVNT\, C => I_16, Y => N_55);
    
    \FID_6_r[3]\ : OA21
      port map(A => N_309_i, B => \FID_6_0_iv_0_0_0_i[3]\, C => 
        N_532_3_6, Y => \FID_6[3]\);
    
    \CRC32_2_i_0[12]\ : NOR2FT
      port map(A => N_532_3_1, B => N_256_i_i_0, Y => N_1290);
    
    \EVENT_DWORD_17_i_0_a2[13]\ : NOR2
      port map(A => \EVENT_DWORD[23]_net_1\, B => N_190_i_0, Y
         => N_338);
    
    \FID_6_iv_0_0_a2_0[23]\ : OR2FT
      port map(A => REG_66, B => N_1574_1, Y => N_1486);
    
    un1_STATE1_17_i_0_0_a2 : NOR2FT
      port map(A => \STATE1_0[3]_net_1\, B => N_176, Y => N_304);
    
    EVNT_NUM_2_I_47 : XOR2
      port map(A => \EVNT_NUM[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, Y => \EVNT_NUM_2[2]\);
    
    \CRC32_2_i_0[22]\ : NOR2FT
      port map(A => N_532_3_2, B => N_1782_i_0, Y => N_1292);
    
    CHANNEL_132 : MUX2H
      port map(A => \CHANNEL[2]_net_1\, B => N_99, S => 
        I2C_RREQ_1_sqmuxa, Y => \CHANNEL_132\);
    
    \un2_i2c_chain_0_0_0_o2[4]\ : NOR2
      port map(A => \CNT[1]_net_1\, B => \CNT[2]_net_1\, Y => 
        N_197);
    
    un1_I2C_RREQ_1_sqmuxa_0_0_0 : OAI21FTT
      port map(A => N_293, B => N_215, C => N_532_3_0, Y => 
        un1_I2C_RREQ_1_sqmuxa);
    
    \FID_6_r[26]\ : OA21
      port map(A => N_1496_i, B => \FID_6_iv_0_0_0_i[26]\, C => 
        N_532_3_4, Y => \FID_6[26]\);
    
    un2_bnc_cnt_I_59 : AND3
      port map(A => \BNC_CNT[6]_net_1\, B => \BNC_CNT[7]_net_1\, 
        C => \BNC_CNT[8]_net_1\, Y => \DWACT_FINC_E[5]\);
    
    un1_REG_1_ADD_16x16_slow_I7_CO1_0_a0_3 : OR3
      port map(A => un5_evread_7, B => \REG[32]\, C => \REG[33]\, 
        Y => ADD_16x16_slow_I7_CO1_0_a0_3_i);
    
    \un2_i2c_chain_0_0_0_o2_0[6]\ : NAND2
      port map(A => N_1765, B => N_1775, Y => N_1612);
    
    un1_RDY_CNT_I_10 : XOR2
      port map(A => \RDY_CNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP_1[0]\, Y => I_10);
    
    BNC_CNT_220 : MUX2H
      port map(A => \BNC_CNT[4]_net_1\, B => \BNC_CNT_3[4]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_220\);
    
    \CRC32[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_116\, CLR => CLEAR_7, 
        Q => \CRC32[23]_net_1\);
    
    \CRC32[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_108\, CLR => CLEAR_6, 
        Q => \CRC32[15]_net_1\);
    
    \STATE2_ns_0_0[2]\ : AO21FTT
      port map(A => \STATE2[2]_net_1\, B => \TRIGGER_sync\, C => 
        \STATE2[1]_net_1\, Y => \STATE2_ns[2]\);
    
    \FID[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_176\, CLR => CLEAR_15, Q
         => \FID[6]_net_1\);
    
    \FID[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_180\, CLR => CLEAR_13, Q
         => \FID[10]_net_1\);
    
    \EVNT_NUM[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[9]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[9]_net_1\);
    
    \un2_i2c_chain_0_0_0_a2_2_1[3]\ : NOR2
      port map(A => \CNT[2]_net_1\, B => N_1765, Y => N_312_1);
    
    un2_bnc_cnt_I_115 : XOR2
      port map(A => N_81_0, B => \BNC_CNT[18]_net_1\, Y => I_115);
    
    un2_bnc_cnt_I_165 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[18]\, Y => N_45);
    
    L1AS_1 : OR3
      port map(A => \L1AF1\, B => \L1AF2\, C => \L1AF3\, Y => 
        \L1AS_1\);
    
    un1_REG_1_ADD_16x16_slow_I5_CO1 : AO21TTF
      port map(A => I4_un1_CO1, B => \REG[37]\, C => 
        ADD_16x16_slow_I5_CO1_0, Y => N216);
    
    un1_EVENT_DWORD_0_sqmuxa_0_o5_0_a2_0_a2_0_a2 : NOR2FT
      port map(A => \OR_RACK_sync\, B => N_1762, Y => N_1454);
    
    EVNT_NUM_2_I_60 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_0[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_0[0]\);
    
    \FID_6_iv_0_0_a2_1[12]\ : NOR2FT
      port map(A => \EVENT_DWORD[12]_net_1\, B => N_620_4_0, Y
         => N_1508_i);
    
    un2_bnc_cnt_I_125 : AND2
      port map(A => \BNC_CNT[18]_net_1\, B => \BNC_CNT[19]_net_1\, 
        Y => \DWACT_FINC_E[14]\);
    
    \FID_6_iv_0_0_0[20]\ : OAI21FTT
      port map(A => \EVNT_NUM[4]_net_1\, B => N_1575_1, C => 
        N_1480, Y => \FID_6_iv_0_0_0_i[20]\);
    
    DTEST_FIFO_87 : MUX2H
      port map(A => DTEST_FIFO_net_1, B => N_532_3, S => N_795, Y
         => \DTEST_FIFO_87\);
    
    FID_179 : MUX2H
      port map(A => \FID[9]_net_1\, B => \FID_6[9]\, S => N_205, 
        Y => \FID_179\);
    
    un1_REG_1_ADD_16x16_slow_I1_CO1_0 : OAI21FTF
      port map(A => \un5_evread_1\, B => \REG[33]\, C => 
        \un2_evread[14]\, Y => ADD_16x16_slow_I1_CO1_0);
    
    \un2_i2c_chain_0_0_0_o2_0[3]\ : OR2FT
      port map(A => N_219, B => \CNT[5]_net_1\, Y => N_1603);
    
    \CRC32_2_i_0_x2[31]\ : XOR2FT
      port map(A => \CRC32[31]_net_1\, B => 
        \EVENT_DWORD[31]_net_1\, Y => N_276_i_i_0);
    
    L2AF2 : DFFC
      port map(CLK => ALICLK_c, D => \L2AF1\, CLR => HWRES_c_12, 
        Q => \L2AF2\);
    
    BNC_CNT_243 : MUX2H
      port map(A => \BNC_CNT[27]_net_1\, B => 
        \BNC_CNT_3[27]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_243\);
    
    \FID[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_173\, CLR => CLEAR_15, Q
         => \FID[3]_net_1\);
    
    \BNC_CNT[15]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_231\, CLR => 
        CLEAR_2, Q => \BNC_CNT[15]_net_1\);
    
    un1_REG_1_G_10_0_o2 : OR3
      port map(A => I6_un4_CO1, B => N_55, C => N_54, Y => 
        I6_un1_CO1_i_0_i);
    
    un1_REG_1_ADD_16x16_slow_I8_un1_CO1_0_tz_0 : OR2
      port map(A => ADD_16x16_slow_I7_CO1_0, B => \REG[40]\, Y
         => ADD_16x16_slow_I8_un1_CO1_0_tz_0);
    
    \FID[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_196\, CLR => CLEAR_14, Q
         => \FID[26]_net_1\);
    
    un4_bnc_res_NE_15 : OR3
      port map(A => un4_bnc_res_NE_1_i, B => un4_bnc_res_20_i_i, 
        C => un4_bnc_res_23_i_i, Y => un4_bnc_res_NE_15_i);
    
    \FID_2_0[10]\ : XOR2
      port map(A => \CRC32[18]_net_1\, B => \CRC32[30]_net_1\, Y
         => \FID_2_0[10]_net_1\);
    
    un1_REG_1_G_8_0_x2 : XOR2
      port map(A => I_16, B => \FIFO_END_EVNT\, Y => G_8_0_x2);
    
    \STATE1_ns_1_iv_0_0_a3_2[0]\ : OR3FTT
      port map(A => N_1601, B => \STATE1[3]_net_1\, C => N_1183_i, 
        Y => N_1750);
    
    un2_bnc_cnt_I_162 : AND2
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        Y => \DWACT_FINC_E[18]\);
    
    \FID_6_iv_0_0_a2_1[25]\ : NOR2FT
      port map(A => \EVENT_DWORD[25]_net_1\, B => N_620_4, Y => 
        N_1493_i);
    
    \FID_6_iv_0_0_0[9]\ : OAI21TTF
      port map(A => N_1574, B => REG_52, C => N_1526, Y => 
        \FID_6_iv_0_0_0[9]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2[6]\ : NOR2
      port map(A => \EVENT_DWORD[6]_net_1\, B => N_1229_i, Y => 
        N_1648);
    
    \EVENT_DWORD[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_143\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[5]_net_1\);
    
    \un2_i2c_chain_0_0_0_1[1]\ : AOI21TTF
      port map(A => N_219, B => N_1629_1, C => N_1631, Y => 
        \un2_i2c_chain_0_0_0_1[1]_net_1\);
    
    \EVENT_DWORD_17_i_0_0[10]\ : OAI21TTF
      port map(A => \EVENT_DWORD[18]_net_1\, B => N_105_i_0_1, C
         => N_1652, Y => \EVENT_DWORD_17_i_0_0[10]_net_1\);
    
    \EVENT_DWORD_17_i_0_0[21]\ : OAI21TTF
      port map(A => \EVENT_DWORD[29]_net_1\, B => N_105_i_0_0, C
         => N_1719, Y => \EVENT_DWORD_17_i_0_0[21]_net_1\);
    
    un2_bnc_cnt_I_38 : XOR2
      port map(A => N_136, B => \BNC_CNT[7]_net_1\, Y => I_38_0);
    
    un2_bnc_cnt_I_122 : XOR2
      port map(A => N_76, B => \BNC_CNT[19]_net_1\, Y => I_122);
    
    \BNC_CNT[23]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_239\, CLR => 
        CLEAR_3, Q => \BNC_CNT[23]_net_1\);
    
    \FID_6_iv_0_0_0[16]\ : OAI21FTT
      port map(A => \EVNT_NUM[0]_net_1\, B => N_1575_1, C => 
        N_1533, Y => \FID_6_iv_0_0_0_i[16]\);
    
    \EVENT_DWORD[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_165\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[27]_net_1\);
    
    \CHIP_ADDR[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \CHIP_ADDR_135\, CLR => 
        CLEAR_5, Q => \CHIP_ADDR[2]_net_1\);
    
    un1_EVENT_DWORD_0_sqmuxa_0_0 : NAND2
      port map(A => N_234, B => N_520, Y => 
        \un1_EVENT_DWORD_0_sqmuxa_0_0\);
    
    \FID_6_iv_0_0_a2_2[18]\ : NOR2FT
      port map(A => \EVENT_DWORD[18]_net_1\, B => N_620_4_1, Y
         => N_1550_i);
    
    \EVENT_DWORD_17_r[9]\ : AND3FFT
      port map(A => N_295, B => \EVENT_DWORD_17_i_0[9]_net_1\, C
         => N_532_3_8, Y => \EVENT_DWORD_17[9]\);
    
    EVNT_NUM_2_I_48 : XOR2
      port map(A => \EVNT_NUM[11]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_4[0]\, Y => \EVNT_NUM_2[11]\);
    
    \FID_6_r[20]\ : OA21
      port map(A => N_1481_i, B => \FID_6_iv_0_0_0_i[20]\, C => 
        N_532_3_4, Y => \FID_6[20]\);
    
    OR_RADDR_207 : MUX2H
      port map(A => \OR_RADDR[3]_net_1\, B => N_683, S => N_248, 
        Y => \OR_RADDR_207\);
    
    BNC_CNT_232 : MUX2H
      port map(A => \BNC_CNT[16]_net_1\, B => 
        \BNC_CNT_3[16]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_232\);
    
    N_1470_i : INV
      port map(A => N_1470, Y => N_1470_i_0);
    
    \BNC_CNT[7]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_223\, CLR => 
        CLEAR_4, Q => \BNC_CNT[7]_net_1\);
    
    FAULT_STROBE_0_2_i : OR2FT
      port map(A => REG_c(23), B => \CLEAR_PSM_FLAGS\, Y => 
        \FAULT_STROBE_0_2_i\);
    
    \STATE1_ns_1_iv_0_1_o2_2_0_o2[0]\ : NAND2
      port map(A => \RDY_CNT[0]_net_1\, B => \RDY_CNT[1]_net_1\, 
        Y => N_243);
    
    \FID_2[11]\ : XOR2FT
      port map(A => \CRC32[7]_net_1\, B => \FID_2_0[11]_net_1\, Y
         => \FID_2_i[11]\);
    
    \BNC_CNT_3[19]\ : AND2
      port map(A => I_122, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[19]_net_1\);
    
    EVENT_DWORD_140 : MUX2H
      port map(A => \EVENT_DWORD[2]_net_1\, B => 
        \EVENT_DWORD_17[2]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_140\);
    
    un2_bnc_cnt_I_80 : AND2
      port map(A => \BNC_CNT[12]_net_1\, B => \BNC_CNT[13]_net_1\, 
        Y => \DWACT_FINC_E[8]\);
    
    \EVENT_DWORD_17_i_0_a2[23]\ : NOR2
      port map(A => \EVENT_DWORD[23]_net_1\, B => N_1229_i_0, Y
         => N_1714);
    
    \FID_6_r[22]\ : OA21
      port map(A => N_1514_i, B => \FID_6_iv_0_0_0_i[22]\, C => 
        N_532_3_4, Y => \FID_6[22]\);
    
    STATE1_tr10_0_a3_0_a2 : AND2
      port map(A => N_1573, B => N_1585, Y => \STATE1_d[9]\);
    
    \FID_6_iv_0_0_a2[17]\ : OR2FT
      port map(A => \EVNT_NUM[1]_net_1\, B => N_1575_1, Y => 
        N_1552);
    
    un4_bnc_res_4 : XOR2
      port map(A => \BNC_CNT[4]_net_1\, B => REG_408, Y => 
        un4_bnc_res_4_i_i);
    
    \REG_1[39]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I7_S, CLR => 
        CLEAR_18, Q => \REG[39]\);
    
    \BNC_CNT_3[16]\ : AND2
      port map(A => I_98, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[16]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I3_S : XOR2
      port map(A => I2_un1_CO1, B => ADD_16x16_slow_I3_S_0, Y => 
        ADD_16x16_slow_I3_S);
    
    \STATE1_ns_1_iv_0_0_a3_0_1[0]\ : NOR3FFT
      port map(A => \PDL_RACK_sync\, B => N_243, C => 
        \STATE1_0[1]_net_1\, Y => 
        \STATE1_ns_1_iv_0_0_a3_0_1[0]_net_1\);
    
    un1_REG_1_G_14_0_o2 : OR2
      port map(A => ADD_16x16_slow_I7_CO1_0, B => I7_un3_CO1, Y
         => N220);
    
    un1_REG_1_ADD_16x16_slow_I8_S_0 : XOR2FT
      port map(A => \REG[40]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I8_S_0);
    
    un1_REG_1_ADD_16x16_slow_I6_S_0 : XOR2FT
      port map(A => \REG[38]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I6_S_0);
    
    \REG_1[45]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I13_S, CLR => 
        CLEAR_19, Q => \REG[45]\);
    
    \FID_6_r[2]\ : OA21
      port map(A => N_1517_i, B => \FID_6_0_iv_0_0_0_i[2]\, C => 
        N_532_3_6, Y => \FID_6[2]\);
    
    \CNT[4]\ : DFFC
      port map(CLK => CLK_c_c, D => N_84, CLR => CLEAR_6, Q => 
        \CNT[4]_net_1\);
    
    \un2_i2c_chain_0_0_0_a2_4[1]\ : NOR2
      port map(A => \CNT[3]_net_1\, B => N_1767, Y => N_1776);
    
    \PDL_RADDR[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RADDR_215\, CLR => 
        CLEAR_17, Q => \PDL_RADDR[5]_net_1\);
    
    \EVENT_DWORD_17_i_0[19]\ : OAI21TTF
      port map(A => \EVENT_DWORD[27]_net_1\, B => N_105_i_0_1, C
         => N_1675, Y => \EVENT_DWORD_17_i_0[19]_net_1\);
    
    un4_bnc_res_31 : XOR2
      port map(A => \BNC_CNT[31]_net_1\, B => REG_435, Y => 
        un4_bnc_res_31_i_i);
    
    un1_STATE1_11_0_i_m2 : MUX2H
      port map(A => N_1575, B => N_221, S => \STATE1[2]_net_1\, Y
         => N_253);
    
    \FID_6_iv_0_0_a2_1[7]\ : NOR2FT
      port map(A => \EVENT_DWORD[7]_net_1\, B => N_620_4_0, Y => 
        N_320_i);
    
    \CRC32[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_103\, CLR => CLEAR_6, 
        Q => \CRC32[10]_net_1\);
    
    \OR_RADDR[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \OR_RADDR_208\, CLR => 
        CLEAR_16, Q => \OR_RADDR[4]_net_1\);
    
    \CRC32_2_i_0_a2_2[17]\ : OR2FT
      port map(A => N_1585_0, B => N_176_0, Y => N_532_3_2);
    
    un2_bnc_cnt_I_104 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[10]\, C
         => \DWACT_FINC_E[11]\, Y => N_88);
    
    \CRC32_2_i_0_x2[11]\ : XOR2FT
      port map(A => \CRC32[11]_net_1\, B => 
        \EVENT_DWORD[11]_net_1\, Y => N_250_i_i_0);
    
    \un2_i2c_chain_0_0_0_a2[6]\ : NOR3FFT
      port map(A => \CNT_0[0]_net_1\, B => N_1612, C => N_1766, Y
         => N_1637_i);
    
    \STATE1_ns_i_0_o2_0[1]\ : OR3FTT
      port map(A => I2C_RACK, B => N_222, C => N_120_i, Y => 
        N_289);
    
    \CNT[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_8_i[5]_net_1\, CLR => 
        CLEAR_6, Q => \CNT[5]_net_1\);
    
    \CRC32_2_i_0[13]\ : NOR2FT
      port map(A => N_532_3_1, B => N_284_i_i_0, Y => N_1380);
    
    un4_bnc_res_13 : XOR2
      port map(A => \BNC_CNT[13]_net_1\, B => REG_417, Y => 
        un4_bnc_res_13_i_i);
    
    \PDL_RADDR[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RADDR_213\, CLR => 
        CLEAR_17, Q => \PDL_RADDR[3]_net_1\);
    
    \CRC32_2_i_0[23]\ : NOR2FT
      port map(A => N_532_3_2, B => N_1781_i_0, Y => N_1221);
    
    TRIGGER_sync : DFFC
      port map(CLK => CLK_c_c, D => \BNC_LIMIT_stretched\, CLR
         => CLEAR_20, Q => \TRIGGER_sync\);
    
    un1_REG_1_ADD_16x16_slow_I4_un1_CO1_0_a0_1 : OR2FT
      port map(A => ADD_16x16_slow_I4_un1_CO1_0_a0_0, B => 
        \REG[33]\, Y => ADD_16x16_slow_I4_un1_CO1_0_a0_1_i);
    
    un1_REG_1_ADD_16x16_slow_I13_S_0 : XOR2FT
      port map(A => \REG[45]\, B => \un2_evread_1[14]\, Y => 
        ADD_16x16_slow_I13_S_0);
    
    FID_177 : MUX2H
      port map(A => \FID[7]_net_1\, B => \FID_6[7]\, S => N_205, 
        Y => \FID_177\);
    
    \EVENT_DWORD_17_i_a2_0[29]\ : NOR2
      port map(A => \EVENT_DWORD[29]_net_1\, B => N_1229_i_0, Y
         => N_1683);
    
    \CHANNEL[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \CHANNEL_131\, CLR => CLEAR_5, 
        Q => \CHANNEL[1]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I15_Y : XOR2
      port map(A => ADD_16x16_slow_I15_Y_0, B => 
        I14_un1_CO1_i_0_i, Y => ADD_16x16_slow_I15_Y);
    
    CHIP_ADDR_134 : MUX2H
      port map(A => \CHIP_ADDR[1]_net_1\, B => N_721_i_0, S => 
        I2C_RREQ_1_sqmuxa, Y => \CHIP_ADDR_134\);
    
    un1_CNT_1_I_28 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \CNT_0[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \un2_i2c_chain_0_i_0_a2[2]\ : NOR2FT
      port map(A => N_213, B => N_1763, Y => N_298_i);
    
    \CRC32_2_i_0_x2[4]\ : XOR2FT
      port map(A => \CRC32[4]_net_1\, B => \EVENT_DWORD[4]_net_1\, 
        Y => N_274_i_i_0);
    
    FID_190 : MUX2H
      port map(A => \FID[20]_net_1\, B => \FID_6[20]\, S => 
        N_205_1, Y => \FID_190\);
    
    un1_ORATETMO_1_I_12 : XOR2
      port map(A => \ORATETMO_i_i[3]\, B => N_701_i_0_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\);
    
    \CRC32[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_98\, CLR => CLEAR_8, Q
         => \CRC32[5]_net_1\);
    
    un1_STATE1_19_i_i_0 : NAND3FTT
      port map(A => N_1587, B => N_522, C => N_253, Y => N_205_0);
    
    \STATE1_ns_1_iv_0_1_o2_3_a3[0]\ : NOR3FTT
      port map(A => \STATE1[0]_net_1\, B => \STATE1[1]_net_1\, C
         => N_237, Y => N_1744);
    
    \FID_6_iv_0_0_a2_0[25]\ : OR2FT
      port map(A => REG_68, B => N_1574, Y => N_1492);
    
    \un2_i2c_chain_0_i_0_a3_0[2]\ : OR2FT
      port map(A => \CNT_0[5]_net_1\, B => \CNT_0[4]_net_1\, Y
         => N_1765);
    
    un4_bnc_res_NE_9 : OR2
      port map(A => un4_bnc_res_24_i_i, B => un4_bnc_res_27_i_i, 
        Y => un4_bnc_res_NE_9_i);
    
    un2_bnc_cnt_I_195 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[30]\, 
        C => \DWACT_FINC_E[23]\, Y => N_24);
    
    EVNT_NUM_2_I_45 : XOR2
      port map(A => \EVNT_NUM[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP_0[0]\, Y => \EVNT_NUM_2[1]\);
    
    \CRC32[30]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_123\, CLR => CLEAR_8, 
        Q => \CRC32[30]_net_1\);
    
    READ_PDL_FLAG : DFFC
      port map(CLK => CLK_c_c, D => \READ_PDL_FLAG_92_0_0\, CLR
         => CLEAR_18, Q => \READ_PDL_FLAG\);
    
    \CRC32[29]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_122\, CLR => CLEAR_8, 
        Q => \CRC32[29]_net_1\);
    
    \EVENT_DWORD[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_146\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[8]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2[2]\ : NOR2
      port map(A => \EVENT_DWORD[2]_net_1\, B => N_1229_i, Y => 
        N_1644);
    
    \CRC32_2_i_0[17]\ : NOR2FT
      port map(A => N_532_3_1, B => N_1779_i_0, Y => N_1140);
    
    \CRC32_2_i_0[27]\ : NOR2FT
      port map(A => N_532_3_2, B => N_242_i_i_0, Y => N_1142);
    
    \EVENT_DWORD[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_153\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[15]_net_1\);
    
    \CRC32_2_i_0_a2_5[17]\ : OR2FT
      port map(A => N_1585_0, B => N_176_0, Y => N_532_3_5);
    
    \EVENT_DWORD_17_i_a2_0[19]\ : NOR2
      port map(A => \EVENT_DWORD[19]_net_1\, B => N_1229_i_1, Y
         => N_1676);
    
    \CRC32_2_i_0_a2[17]\ : OR2FT
      port map(A => N_1585, B => N_176, Y => N_532_3);
    
    un4_bnc_res_23 : XOR2
      port map(A => \BNC_CNT[23]_net_1\, B => REG_427, Y => 
        un4_bnc_res_23_i_i);
    
    EVENT_DWORD_169 : MUX2H
      port map(A => \EVENT_DWORD[31]_net_1\, B => 
        \EVENT_DWORD_17[31]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_169\);
    
    un2_bnc_cnt_I_114 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[10]\, 
        C => \DWACT_FINC_E[12]\, Y => N_81_0);
    
    \CRC32[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_110\, CLR => CLEAR_7, 
        Q => \CRC32[17]_net_1\);
    
    FID_176 : MUX2H
      port map(A => \FID[6]_net_1\, B => \FID_6[6]\, S => N_205, 
        Y => \FID_176\);
    
    CRC32_98 : MUX2H
      port map(A => \CRC32[5]_net_1\, B => N_1376, S => N_1469, Y
         => \CRC32_98\);
    
    FID_178 : MUX2H
      port map(A => \FID[8]_net_1\, B => \FID_6[8]\, S => N_205, 
        Y => \FID_178\);
    
    un2_bnc_cnt_I_192 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        C => \DWACT_FINC_E[22]\, Y => \DWACT_FINC_E[23]\);
    
    un2_bnc_cnt_I_172 : AND3
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[19]\, Y => N_40);
    
    un1_CNT_1_I_1 : AND2
      port map(A => \CNT[0]_net_1\, B => 
        \un1_EVENT_DWORD_0_sqmuxa_0_0\, Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    \EVENT_DWORD_17_r[23]\ : AND3FFT
      port map(A => N_1714, B => \EVENT_DWORD_17_i_0_1[23]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[23]\);
    
    un4_bnc_res_NE_21 : OR3
      port map(A => un4_bnc_res_NE_11_i, B => un4_bnc_res_8_i_i, 
        C => un4_bnc_res_9_i_i, Y => un4_bnc_res_NE_21_i);
    
    \STATE1_ns_0_0_a2_1_a2_0_a2[3]\ : NOR2FT
      port map(A => N_1573, B => N_120_i, Y => N_1195_1);
    
    \ORATETMO_7_0_0[2]\ : OR2
      port map(A => N_233, B => I_20_2, Y => \ORATETMO_7[2]\);
    
    \EVENT_DWORD_17_i_0_a2[7]\ : NOR2
      port map(A => \EVENT_DWORD[17]_net_1\, B => N_190_i, Y => 
        N_1620);
    
    un1_ORATETMO_1_I_24 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0_2[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_1_0[0]\);
    
    \un2_i2c_chain_0_0_0_a2_1[4]\ : OR3
      port map(A => N_219, B => N_1763, C => N_197, Y => 
        \un2_i2c_chain_0_0_0_a2_1[4]_net_1\);
    
    \STATE1_ns_1_iv_0_0_o2[2]\ : NAND2FT
      port map(A => \RDY_CNT[0]_net_1\, B => \RDY_CNT[1]_net_1\, 
        Y => N_222);
    
    READ_PDL_FLAG_92_0_0_a2 : OR3FFT
      port map(A => \READ_PDL_FLAG\, B => N_266, C => 
        \STATE1_0[1]_net_1\, Y => N_1669_i);
    
    event_meb : event_fifo
      port map(FID(31) => \FID[31]_net_1\, FID(30) => 
        \FID[30]_net_1\, FID(29) => \FID[29]_net_1\, FID(28) => 
        \FID[28]_net_1\, FID(27) => \FID[27]_net_1\, FID(26) => 
        \FID[26]_net_1\, FID(25) => \FID[25]_net_1\, FID(24) => 
        \FID[24]_net_1\, FID(23) => \FID[23]_net_1\, FID(22) => 
        \FID[22]_net_1\, FID(21) => \FID[21]_net_1\, FID(20) => 
        \FID[20]_net_1\, FID(19) => \FID[19]_net_1\, FID(18) => 
        \FID[18]_net_1\, FID(17) => \FID[17]_net_1\, FID(16) => 
        \FID[16]_net_1\, FID(15) => \FID[15]_net_1\, FID(14) => 
        \FID[14]_net_1\, FID(13) => \FID[13]_net_1\, FID(12) => 
        \FID[12]_net_1\, FID(11) => \FID[11]_net_1\, FID(10) => 
        \FID[10]_net_1\, FID(9) => \FID[9]_net_1\, FID(8) => 
        \FID[8]_net_1\, FID(7) => \FID[7]_net_1\, FID(6) => 
        \FID[6]_net_1\, FID(5) => \FID[5]_net_1\, FID(4) => 
        \FID[4]_net_1\, FID(3) => \FID[3]_net_1\, FID(2) => 
        \FID[2]_net_1\, FID(1) => \FID[1]_net_1\, FID(0) => 
        \FID[0]_net_1\, DPR(31) => DPR(31), DPR(30) => DPR(30), 
        DPR(29) => DPR(29), DPR(28) => DPR(28), DPR(27) => 
        DPR(27), DPR(26) => DPR(26), DPR(25) => DPR(25), DPR(24)
         => DPR(24), DPR(23) => DPR(23), DPR(22) => DPR(22), 
        DPR(21) => DPR(21), DPR(20) => DPR(20), DPR(19) => 
        DPR(19), DPR(18) => DPR(18), DPR(17) => DPR(17), DPR(16)
         => DPR(16), DPR(15) => DPR(15), DPR(14) => DPR(14), 
        DPR(13) => DPR(13), DPR(12) => DPR(12), DPR(11) => 
        DPR(11), DPR(10) => DPR(10), DPR(9) => DPR(9), DPR(8) => 
        DPR(8), DPR(7) => DPR(7), DPR(6) => DPR(6), DPR(5) => 
        DPR(5), DPR(4) => DPR(4), DPR(3) => DPR(3), DPR(2) => 
        DPR(2), DPR(1) => DPR(1), DPR(0) => DPR(0), WRB => \WRB\, 
        CLEAR_i_0 => CLEAR_i_0, NRDMEB => NRDMEB, CLK_c_c => 
        CLK_c_c, FF_c => FF_c, EF => EF);
    
    \CRC32_2_i_0_x2[15]\ : XOR2FT
      port map(A => \CRC32[15]_net_1\, B => 
        \EVENT_DWORD[15]_net_1\, Y => N_251_i_i_0);
    
    un1_REG_1_ADD_16x16_slow_I6_un4_CO1_4 : AOI21TTF
      port map(A => \REG[34]\, B => \REG[33]\, C => 
        \FIFO_END_EVNT\, Y => N_7210_i);
    
    un2_bnc_cnt_I_48 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[3]\, Y => \DWACT_FINC_E[4]\);
    
    PDL_RREQ_136 : MUX2H
      port map(A => PDL_RREQ_net_1, B => N_1195_1, S => 
        un1_STATE1_1_sqmuxa, Y => \PDL_RREQ_136\);
    
    \CRC32_2_i_0_a2_1[17]\ : OR2FT
      port map(A => N_1585, B => N_176_0, Y => N_532_3_1);
    
    EVENT_DWORD_142 : MUX2H
      port map(A => \EVENT_DWORD[4]_net_1\, B => 
        \EVENT_DWORD_17[4]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_142\);
    
    \EVENT_DWORD[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_160\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[22]_net_1\);
    
    BNC_CNT_242 : MUX2H
      port map(A => \BNC_CNT[26]_net_1\, B => 
        \BNC_CNT_3[26]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_242\);
    
    \REG_1[37]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I5_S, CLR => 
        CLEAR_18, Q => \REG[37]\);
    
    OR_RREQ_203 : MUX2H
      port map(A => OR_RREQ_net_1, B => N_252_i_0, S => N_203, Y
         => \OR_RREQ_203\);
    
    un1_CNT_1_I_21 : XOR2
      port map(A => \CNT[1]_net_1\, B => \DWACT_ADD_CI_0_TMP[0]\, 
        Y => I_21_0);
    
    \FID_6_iv_0_0_x2[14]\ : XOR2FT
      port map(A => \CRC32[10]_net_1\, B => \CRC32[22]_net_1\, Y
         => N_270_i_0_i);
    
    CRC32_119 : MUX2H
      port map(A => \CRC32[26]_net_1\, B => N_1384, S => N_1469_0, 
        Y => \CRC32_119\);
    
    \un2_i2c_chain_0_0_0[1]\ : OR3
      port map(A => \un2_i2c_chain_0_0_0_3_i[1]\, B => 
        \un2_i2c_chain_0_0_0_0_i[1]\, C => N_1776, Y => N_94);
    
    N_105_i_0_a2_0_a2_1 : OR2
      port map(A => \STATE1_0[0]_net_1\, B => N_176, Y => 
        N_105_i_0_1);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_0 : MUX2L
      port map(A => \REG[43]\, B => \un2_evread_i_0[14]\, S => 
        ADD_16x16_slow_I14_un1_CO1_N_16_i_i, Y => 
        I14_un1_CO1_i_0_i);
    
    OR_RADDR_206 : MUX2H
      port map(A => \OR_RADDR[2]_net_1\, B => N_685, S => N_248, 
        Y => \OR_RADDR_206\);
    
    \EVENT_DWORD_17_r[29]\ : AND3FFT
      port map(A => N_1683, B => \EVENT_DWORD_17_i_1[29]_net_1\, 
        C => N_532_3_6, Y => \EVENT_DWORD_17[29]\);
    
    \EVENT_DWORD_17_r[20]\ : AND3FFT
      port map(A => N_1702, B => \EVENT_DWORD_17_i_0_1[20]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[20]\);
    
    \FID_6_0_iv_0_a2_3[1]\ : OR2FT
      port map(A => \EVENT_DWORD[1]_net_1\, B => N_620_4_0, Y => 
        N_1505);
    
    \un2_i2c_chain_0_0_0_a2_4[4]\ : OR3
      port map(A => N_1766, B => \CNT_0[0]_net_1\, C => 
        \CNT[5]_net_1\, Y => N_1692);
    
    \FID_6_iv_0_0_a2_1[10]\ : NOR2FT
      port map(A => \EVENT_DWORD[10]_net_1\, B => N_620_4_0, Y
         => N_1472_i);
    
    EVRDYi_202_i : INV
      port map(A => EVREAD, Y => EVREAD_i_0);
    
    un1_REG_1_ADD_16x16_slow_I6_un4_CO1_6_tz : NAND3
      port map(A => ADD_16x16_slow_I6_un4_CO1_6_tz_0, B => 
        \REG[32]\, C => \REG[36]\, Y => 
        ADD_16x16_slow_I6_un4_CO1_5_tz);
    
    \FID_6_iv_0_0_0[18]\ : AOI21TTF
      port map(A => \FAULT_STAT\, B => N_1587, C => N_1547, Y => 
        \FID_6_iv_0_0_0[18]_net_1\);
    
    \CRC32_2_i_0[16]\ : NOR2FT
      port map(A => N_532_3_1, B => N_1783_i_0, Y => N_1381);
    
    \EVENT_DWORD_17_i_0_a2_0[2]\ : NOR2
      port map(A => \EVENT_DWORD[12]_net_1\, B => N_190_i, Y => 
        N_1645);
    
    \EVENT_DWORD_17_i_0_a2_0[26]\ : NOR2
      port map(A => I2C_RDATA(6), B => N_1768_i, Y => N_1699);
    
    FID_184 : MUX2H
      port map(A => \FID[14]_net_1\, B => \FID_6[14]\, S => 
        N_205_1, Y => \FID_184\);
    
    \CRC32_2_i_0[26]\ : NOR2FT
      port map(A => N_532_3_2, B => N_287_i_i_0, Y => N_1384);
    
    un1_REG_1_ADD_16x16_slow_I13_CO1_0_a0_5 : NOR3
      port map(A => ADD_16x16_slow_I7_CO1_0, B => 
        ADD_16x16_slow_I13_CO1_0_a0_2_i, C => 
        ADD_16x16_slow_I13_CO1_0_a0_3_i, Y => 
        ADD_16x16_slow_I13_CO1_0_a0_5);
    
    \REG_1[40]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I8_S, CLR => 
        CLEAR_18, Q => \REG[40]\);
    
    \EVENT_DWORD_17_i_0_a2[10]\ : NOR2
      port map(A => \EVENT_DWORD[10]_net_1\, B => N_1229_i_1, Y
         => N_1651);
    
    CRC32_99 : MUX2H
      port map(A => \CRC32[6]_net_1\, B => N_1377, S => N_1469, Y
         => \CRC32_99\);
    
    \EVENT_DWORD_17_r[11]\ : AND3FFT
      port map(A => N_336, B => \EVENT_DWORD_17_i_0_0[11]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[11]\);
    
    \FID_6_iv_0_0_a2_1[8]\ : NOR2
      port map(A => \EVENT_DWORD[8]_net_1\, B => N_620_4, Y => 
        N_1525);
    
    CYC_STAT : DFFC
      port map(CLK => CLK_c_c, D => \CYC_STAT_89\, CLR => CLEAR_9, 
        Q => \CYC_STAT\);
    
    \STATE1_ns_0_0_0_o2[3]\ : NAND2
      port map(A => N_243, B => N_1601, Y => N_230);
    
    \un2_i2c_chain_0_i_0[2]\ : NOR3
      port map(A => \un2_i2c_chain_0_i_0_3_i[2]\, B => N_298_i, C
         => \un2_i2c_chain_0_i_0_2_i[2]\, Y => N_721_i_0);
    
    BNC_LIMIT_stretched_1 : OR2
      port map(A => \BNC_LIMIT\, B => \BNC_LIMIT_r\, Y => 
        \BNC_LIMIT_stretched_1\);
    
    \FID_6_iv_0_0_a2[5]\ : NOR2
      port map(A => \FID_2[5]_net_1\, B => N_1575, Y => N_1520);
    
    \CNT_8_i_a3_2_1[0]\ : NOR2FT
      port map(A => \STATE1_0[1]_net_1\, B => \STATE1_0[0]_net_1\, 
        Y => N_1758_1);
    
    \FID_2[5]\ : XOR2
      port map(A => \CRC32[1]_net_1\, B => \FID_2_0[5]_net_1\, Y
         => \FID_2[5]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I9_CO1_0_tz_0 : NOR2FT
      port map(A => ADD_16x16_slow_I8_un1_CO1_0, B => \REG[41]\, 
        Y => ADD_16x16_slow_I9_CO1_0_tz_0);
    
    \FID_6_r[15]\ : OA21
      port map(A => N_1478_i, B => \FID_6_iv_0_0_0_i[15]\, C => 
        N_532_3_5, Y => \FID_6[15]\);
    
    \CRC32_2_i_x2[19]\ : XOR2FT
      port map(A => \CRC32[19]_net_1\, B => 
        \EVENT_DWORD[19]_net_1\, Y => N_273_i_i_0);
    
    \CRC32_2_i_0_x2[14]\ : XOR2FT
      port map(A => \CRC32[14]_net_1\, B => 
        \EVENT_DWORD[14]_net_1\, Y => N_257_i_i_0);
    
    un1_REG_1_ADD_16x16_slow_I5_S : XOR2
      port map(A => I4_un1_CO1, B => ADD_16x16_slow_I5_S_0, Y => 
        ADD_16x16_slow_I5_S);
    
    \FID_6_0_iv_0_a2_2_0_a2_0[3]\ : OR2
      port map(A => \STATE1_0[3]_net_1\, B => N_176_0, Y => 
        N_1574_0);
    
    un1_REG_1_ADD_16x16_slow_I15_Y_0 : XOR2FT
      port map(A => \REG[47]\, B => \un2_evread[14]\, Y => 
        ADD_16x16_slow_I15_Y_0);
    
    \EVENT_DWORD[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_162\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[24]_net_1\);
    
    EVENT_DWORD_159 : MUX2H
      port map(A => \EVENT_DWORD[21]_net_1\, B => 
        \EVENT_DWORD_17[21]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_159\);
    
    \CRC32[25]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_118\, CLR => CLEAR_7, 
        Q => \CRC32[25]_net_1\);
    
    un4_bnc_res_19 : XOR2
      port map(A => \BNC_CNT[19]_net_1\, B => REG_423, Y => 
        un4_bnc_res_19_i_i);
    
    un1_REG_1_ADD_16x16_slow_I14_S_0 : XOR2FT
      port map(A => \REG[46]\, B => \un2_evread[14]\, Y => 
        ADD_16x16_slow_I14_S_0);
    
    \FID_6_iv_0_0[27]\ : OAI21FTT
      port map(A => \EVNT_NUM[11]_net_1\, B => N_1575, C => 
        N_1543, Y => \FID_6_iv_0_0_i[27]\);
    
    \STATE1_0[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[3]\, CLR => 
        CLEAR_0, Q => \STATE1_0[3]_net_1\);
    
    CRC32_96 : MUX2H
      port map(A => \CRC32[3]_net_1\, B => N_1123, S => N_1469, Y
         => \CRC32_96\);
    
    EVENT_DWORD_144 : MUX2H
      port map(A => \EVENT_DWORD[6]_net_1\, B => 
        \EVENT_DWORD_17[6]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_144\);
    
    READ_PDL_FLAG_92_0_0 : OR3
      port map(A => N_1195_1, B => N_1671, C => 
        \READ_PDL_FLAG_92_0_0_0\, Y => \READ_PDL_FLAG_92_0_0\);
    
    un2_bnc_cnt_I_108 : AND3
      port map(A => \BNC_CNT[15]_net_1\, B => \BNC_CNT[16]_net_1\, 
        C => \BNC_CNT[17]_net_1\, Y => \DWACT_FINC_E[12]\);
    
    un1_RDY_CNT_I_1 : AND2
      port map(A => \RDY_CNT[0]_net_1\, B => 
        \un1_EVENT_DWORD_0_sqmuxa_0_0\, Y => 
        \DWACT_ADD_CI_0_TMP_1[0]\);
    
    \ORATETMO[1]\ : DFFS
      port map(CLK => CLK_c_c, D => \ORATETMO_7[1]\, SET => 
        CLEAR_16, Q => \ORATETMO_i_i[1]\);
    
    \CNT_0[4]\ : DFFC
      port map(CLK => CLK_c_c, D => N_84, CLR => CLEAR_0, Q => 
        \CNT_0[4]_net_1\);
    
    \STATE1_ns_1_iv_0_0_a3_4_1[0]\ : AND2
      port map(A => \STATE1_0[1]_net_1\, B => \STATE1_0[3]_net_1\, 
        Y => N_1752_1);
    
    \RDY_CNT_8_i_0_o2[0]\ : NOR3FTT
      port map(A => N_532_3_3, B => N_1583, C => N_1582, Y => 
        N_267);
    
    \FID_6_iv_0_0_a2_0[14]\ : OR2FT
      port map(A => REG_57, B => N_1574_1, Y => N_1510);
    
    \FID[24]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_194\, CLR => CLEAR_14, Q
         => \FID[24]_net_1\);
    
    FAULT_STROBE_0 : DFFS
      port map(CLK => CLK_c_c, D => \FAULT_STROBE_0_2_i\, SET => 
        HWRES_c_11, Q => FAULT_STROBE_0_i);
    
    \EVENT_DWORD_17_i_0_a2_0[16]\ : NOR2
      port map(A => \EVENT_DWORD[26]_net_1\, B => N_190_i_0, Y
         => N_1661);
    
    BNC_CNT_221 : MUX2H
      port map(A => \BNC_CNT[5]_net_1\, B => \BNC_CNT_3[5]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_221\);
    
    \EVENT_DWORD_17_i_0_a2[8]\ : NOR2
      port map(A => \EVENT_DWORD[8]_net_1\, B => N_1229_i, Y => 
        N_1663);
    
    \STATE1_ns_1_iv_0_0_a3[0]\ : NOR3FTT
      port map(A => \STATE1[3]_net_1\, B => \OR_RACK_sync\, C => 
        N_1601, Y => N_7200_i);
    
    STATE1_tr10_0_a3_0_a2_0_0_a2 : NOR2FT
      port map(A => \STATE1_0[2]_net_1\, B => \STATE1[1]_net_1\, 
        Y => N_1573);
    
    un1_STATE1_17_i_0_i4_1_a2_0_i2_0_a2_i_0 : INV
      port map(A => \STATE1[3]_net_1\, Y => \STATE1_i_0[3]\);
    
    \ORATETMO_7_0_0_a2[0]\ : NOR3FFT
      port map(A => \ORATETMO_7_0_0_a2_0[0]_net_1\, B => N_1576_1, 
        C => \READ_PDL_FLAG\, Y => N_1576_i);
    
    EVENT_DWORD_146 : MUX2H
      port map(A => \EVENT_DWORD[8]_net_1\, B => 
        \EVENT_DWORD_17[8]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_146\);
    
    \EVENT_DWORD[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_139\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[1]_net_1\);
    
    un4_bnc_res_8 : XOR2
      port map(A => \BNC_CNT[8]_net_1\, B => REG_412, Y => 
        un4_bnc_res_8_i_i);
    
    un1_STATE1_19_i_i_1 : NAND3FTT
      port map(A => N_1587, B => N_522, C => N_253, Y => N_205_1);
    
    \CNT_8_i_a3_1[0]\ : OR3
      port map(A => N_120_i, B => N_188, C => \STATE1_0[1]_net_1\, 
        Y => N_1757);
    
    \EVNT_NUM[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[11]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[11]_net_1\);
    
    un1_REG_1_G_10_0_a2_0 : NOR3
      port map(A => ADD_16x16_slow_I6_un1_CO1_0_a0_2, B => 
        \FIFO_END_EVNT\, C => I_16, Y => N_54);
    
    BNC_LIMIT_stretched : DFFC
      port map(CLK => ALICLK_c, D => \BNC_LIMIT_stretched_1\, CLR
         => CLEAR_5, Q => \BNC_LIMIT_stretched\);
    
    \un2_i2c_chain_0_0_0_o2[6]\ : NAND2
      port map(A => \CNT[2]_net_1\, B => \CNT[3]_net_1\, Y => 
        N_199);
    
    un1_STATE1_17_i_0_0_a2_1 : NOR3
      port map(A => N_120_i, B => \STATE1[2]_net_1\, C => 
        PULSE(3), Y => N_306);
    
    \EVENT_DWORD_17_i_0_0[20]\ : OAI21TTF
      port map(A => \EVENT_DWORD[28]_net_1\, B => N_105_i_0_0, C
         => N_1703, Y => \EVENT_DWORD_17_i_0_0[20]_net_1\);
    
    \BNC_CNT[30]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_246\, CLR => 
        CLEAR_4, Q => \BNC_CNT[30]_net_1\);
    
    CRC32_109 : MUX2H
      port map(A => \CRC32[16]_net_1\, B => N_1381, S => N_1469_1, 
        Y => \CRC32_109\);
    
    \EVENT_DWORD_17_i_o2_1_a2[7]\ : NOR2FT
      port map(A => N_176, B => I2C_RACK, Y => N_1755_i);
    
    \FID_6_iv_0_0_a2_1[22]\ : NOR2FT
      port map(A => \EVENT_DWORD[22]_net_1\, B => N_620_4_1, Y
         => N_1514_i);
    
    un1_REG_1_G_26_0_a2 : NOR3
      port map(A => N_43, B => \FIFO_END_EVNT\, C => I_16, Y => 
        ADD_16x16_slow_I6_un1_CO1_0);
    
    N_1205_i_i_o2_2 : OR3
      port map(A => \ORATETMO_i_i[0]\, B => \ORATETMO_i_i[1]\, C
         => \ORATETMO[2]_net_1\, Y => N_1205_i_i_o2_2_i);
    
    BNC_CNT_225 : MUX2H
      port map(A => \BNC_CNT[9]_net_1\, B => \BNC_CNT_3[9]_net_1\, 
        S => LBSP_c_1(2), Y => \BNC_CNT_225\);
    
    FID_171 : MUX2H
      port map(A => \FID[1]_net_1\, B => \FID_6[1]\, S => N_205, 
        Y => \FID_171\);
    
    EVNT_NUM_2_I_67 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_3[0]\);
    
    un2_bnc_cnt_I_87 : AND3
      port map(A => \BNC_CNT[12]_net_1\, B => \BNC_CNT[13]_net_1\, 
        C => \BNC_CNT[14]_net_1\, Y => \DWACT_FINC_E[9]\);
    
    un1_REG_1_ADD_16x16_slow_I6_S : XOR2
      port map(A => N216, B => ADD_16x16_slow_I6_S_0, Y => 
        ADD_16x16_slow_I6_S);
    
    EVNT_NUM_2_I_73 : AND2
      port map(A => \EVNT_NUM[4]_net_1\, B => \EVNT_NUM[5]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    \EVENT_DWORD_17_i_0_0[1]\ : OAI21TTF
      port map(A => \EVENT_DWORD[9]_net_1\, B => N_105_i_0, C => 
        N_329, Y => \EVENT_DWORD_17_i_0_0[1]_net_1\);
    
    \FID_6_iv_0_0_a2_1[6]\ : NOR2FT
      port map(A => \EVENT_DWORD[6]_net_1\, B => N_620_4_0, Y => 
        N_317_i);
    
    un1_REG_1_ADD_16x16_slow_I9_CO1_0 : AO21
      port map(A => ADD_16x16_slow_I9_CO1_0_tz_0, B => I8_un4_CO1, 
        C => \un2_evread_1[14]\, Y => ADD_16x16_slow_I9_CO1_0);
    
    un4_bnc_res_29 : XOR2
      port map(A => \BNC_CNT[29]_net_1\, B => REG_433, Y => 
        un4_bnc_res_29_i_i);
    
    \STATE1_ns_1_iv_0_0_a2_2[2]\ : NOR3FFT
      port map(A => \STATE1_i_0[3]\, B => N_1573, C => N_193, Y
         => N_1559_i);
    
    FID_173 : MUX2H
      port map(A => \FID[3]_net_1\, B => \FID_6[3]\, S => N_205, 
        Y => \FID_173\);
    
    \FID_6_iv_0_0_0[5]\ : OAI21TTF
      port map(A => N_1574, B => REG_48, C => N_1520, Y => 
        \FID_6_iv_0_0_0[5]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2_0[24]\ : NOR2
      port map(A => I2C_RDATA(4), B => N_1768_i, Y => N_1707);
    
    L2AS_1 : OR3
      port map(A => \L2AF1\, B => \L2AF2\, C => \L2AF3\, Y => 
        \L2AS_1\);
    
    \FID_6_iv_0_0_a2_0[7]\ : OR2FT
      port map(A => REG_50, B => N_1574_0, Y => N_319);
    
    EVNT_NUM_2_I_58 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_3[0]\, B => 
        \EVNT_NUM[8]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\);
    
    \EVENT_DWORD_17_i_0_a2_0[8]\ : NOR2
      port map(A => \EVENT_DWORD[18]_net_1\, B => N_190_i, Y => 
        N_1664);
    
    \EVENT_DWORD_17_i_0_1[23]\ : OAI21FTF
      port map(A => N_1454_0, B => OR_RDATA(3), C => 
        \EVENT_DWORD_17_i_0_0[23]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[23]_net_1\);
    
    \EVENT_DWORD_17_r[22]\ : AND3FFT
      port map(A => N_1710, B => \EVENT_DWORD_17_i_0_1[22]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[22]\);
    
    \un2_i2c_chain_0_0_0_a2_0[4]\ : NOR3FFT
      port map(A => N_216, B => N_1764, C => \CNT_0[2]_net_1\, Y
         => N_1688_i);
    
    un5_evread_4 : NOR2
      port map(A => \REG[42]\, B => \REG[41]\, Y => 
        \un5_evread_4\);
    
    \BNC_CNT[0]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_216\, CLR => 
        CLEAR_2, Q => \BNC_CNT[0]_net_1\);
    
    \EVENT_DWORD[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_144\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[6]_net_1\);
    
    \EVENT_DWORD_17_r[3]\ : AND3FFT
      port map(A => N_1618, B => \EVENT_DWORD_17_i_0_0[3]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[3]\);
    
    un2_bnc_cnt_I_118 : AND3
      port map(A => \DWACT_FINC_E[7]\, B => \DWACT_FINC_E[9]\, C
         => \DWACT_FINC_E[12]\, Y => \DWACT_FINC_E[13]\);
    
    \FID_6_iv_0_0_x2[12]\ : XOR2FT
      port map(A => \CRC32[8]_net_1\, B => \CRC32[20]_net_1\, Y
         => N_271_i_0_i);
    
    \CRC32_2_i_0_x2[21]\ : XOR2FT
      port map(A => \CRC32[21]_net_1\, B => 
        \EVENT_DWORD[21]_net_1\, Y => N_275_i_i_0);
    
    \BNC_CNT[19]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_235\, CLR => 
        CLEAR_3, Q => \BNC_CNT[19]_net_1\);
    
    un1_REG_1_G_6 : NOR3
      port map(A => un5_evread_7, B => G_6_0, C => 
        ADD_16x16_slow_I5_CO1_0_a0_0, Y => G_6);
    
    \CRC32_2_i_0[0]\ : NOR2FT
      port map(A => N_532_3_0, B => N_254_i_i_0, Y => N_1287);
    
    EVNT_NUM_2_I_71 : AND2
      port map(A => \EVNT_NUM[2]_net_1\, B => \EVNT_NUM[3]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_0[0]\);
    
    \BNC_CNT_3[28]\ : AND2
      port map(A => I_203, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[28]_net_1\);
    
    \OR_RADDR[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \OR_RADDR_205\, CLR => 
        CLEAR_16, Q => \OR_RADDR[1]_net_1\);
    
    \FID[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_177\, CLR => CLEAR_15, Q
         => \FID[7]_net_1\);
    
    un2_bnc_cnt_I_159 : AND3
      port map(A => \BNC_CNT[21]_net_1\, B => \BNC_CNT[22]_net_1\, 
        C => \BNC_CNT[23]_net_1\, Y => \DWACT_FINC_E[17]\);
    
    \EVENT_DWORD_17_i_0_a2[20]\ : NOR2
      port map(A => \EVENT_DWORD[20]_net_1\, B => N_1229_i_0, Y
         => N_1702);
    
    un2_bnc_cnt_I_128 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[14]\, Y => N_71);
    
    FIFO_END_EVNT : DFFC
      port map(CLK => CLK_c_c, D => \FIFO_END_EVNT_88\, CLR => 
        CLEAR_15, Q => \FIFO_END_EVNT\);
    
    un1_STATE1_2_0_i_a3_i_0 : NAND2
      port map(A => N_532_3_0, B => N_620_4_0, Y => N_1469_0);
    
    \FID_6_iv_0_0_0[17]\ : AOI21TTF
      port map(A => \CYC_STAT\, B => N_1587, C => N_1552, Y => 
        \FID_6_iv_0_0_0[17]_net_1\);
    
    un1_ORATETMO_1_I_6 : AND2
      port map(A => \ORATETMO[2]_net_1\, B => N_701_i_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\);
    
    un1_REG_1_ADD_16x16_slow_I11_CO1_0tt_m3_0_a2 : OR3FTT
      port map(A => ADD_16x16_slow_I14_un1_CO1_m14_2, B => 
        \REG[40]\, C => ADD_16x16_slow_I7_CO1_0, Y => 
        ADD_16x16_slow_I11_CO1_0tt_m3_0_a2);
    
    un1_REG_1_ADD_16x16_slow_I6_un1_CO1_0_a0_1 : NOR2
      port map(A => \REG[35]\, B => \REG[36]\, Y => 
        ADD_16x16_slow_I4_un1_CO1_0_a0_0);
    
    un2_bnc_cnt_I_135 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[15]\, Y => N_66);
    
    \EVENT_DWORD[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_142\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[4]_net_1\);
    
    CLEAR_PSM_FLAGS : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_d[9]\, CLR => CLEAR_5, 
        Q => \CLEAR_PSM_FLAGS\);
    
    \BNC_CNT[3]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_219\, CLR => 
        CLEAR_4, Q => \BNC_CNT[3]_net_1\);
    
    un2_bnc_cnt_I_90 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[7]\, C
         => \DWACT_FINC_E[9]\, Y => N_98_0);
    
    \FID[28]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_198\, CLR => CLEAR_14, Q
         => \FID[28]_net_1\);
    
    \EVENT_DWORD_17_r[6]\ : AND3FFT
      port map(A => N_1648, B => \EVENT_DWORD_17_i_0_0[6]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[6]\);
    
    \OR_RADDR_3_i_0[4]\ : AND2
      port map(A => N_532_3_3, B => \CNT_0[4]_net_1\, Y => N_681);
    
    \FID_6_iv_0_0_a2[8]\ : NOR2
      port map(A => \FID_2[8]_net_1\, B => N_1575, Y => N_1523);
    
    \FID[22]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_192\, CLR => CLEAR_14, Q
         => \FID[22]_net_1\);
    
    \EVENT_DWORD[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_158\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[20]_net_1\);
    
    \FID_6_r[31]\ : OA21
      port map(A => N_1497_i, B => N_1498_i, C => N_532_3_3, Y
         => \FID_6[31]\);
    
    FID_185 : MUX2H
      port map(A => \FID[15]_net_1\, B => \FID_6[15]\, S => 
        N_205_1, Y => \FID_185\);
    
    \EVENT_DWORD_17_i_0_a2_0[14]\ : NOR2
      port map(A => \EVENT_DWORD[24]_net_1\, B => N_190_i_0, Y
         => N_1658);
    
    READ_OR_FLAG : DFFC
      port map(CLK => CLK_c_c, D => \READ_OR_FLAG_91_i_0\, CLR
         => CLEAR_18, Q => \READ_OR_FLAG\);
    
    un1_REG_1_ADD_16x16_slow_I7_CO1_0_a0_1 : OR2
      port map(A => \REG[37]\, B => \REG[36]\, Y => 
        ADD_16x16_slow_I5_CO1_0_a0_0);
    
    \EVENT_DWORD_17_i_0_a2[4]\ : NOR2
      port map(A => \EVENT_DWORD[4]_net_1\, B => N_1229_i, Y => 
        N_326);
    
    \FID_6_iv_0_0_a2_0[16]\ : OR2FT
      port map(A => REG_59, B => N_1574_1, Y => N_1533);
    
    CRC32_114 : MUX2H
      port map(A => \CRC32[21]_net_1\, B => N_1220, S => N_1469_0, 
        Y => \CRC32_114\);
    
    \un2_i2c_chain_0_i_0_a3[2]\ : OR2FT
      port map(A => \CNT_0[4]_net_1\, B => \CNT_0[5]_net_1\, Y
         => N_1763);
    
    \EVENT_DWORD[26]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_164\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[26]_net_1\);
    
    \CRC32[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_113\, CLR => CLEAR_7, 
        Q => \CRC32[20]_net_1\);
    
    un1_REG_1_G_8_0_a2 : NOR3
      port map(A => G_8_0_a2_2, B => G_8_0_x2, C => N_19, Y => 
        I6_un4_CO1);
    
    EVNT_NUM_2_I_68 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_2_0[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    \EVENT_DWORD_17_i_0_a2_0[0]\ : NOR2
      port map(A => \EVENT_DWORD[10]_net_1\, B => N_190_i, Y => 
        N_1642);
    
    un2_bnc_cnt_I_206 : AND2
      port map(A => \BNC_CNT[27]_net_1\, B => \BNC_CNT[28]_net_1\, 
        Y => \DWACT_FINC_E[25]\);
    
    \STATE1_ns_1_iv_0_0_0[2]\ : OA21FTT
      port map(A => \STATE1_ns_1_iv_0_0_a2_3_1[2]_net_1\, B => 
        N_195, C => N_1557, Y => \STATE1_ns_1_iv_0_0_0[2]_net_1\);
    
    \FID_6_iv_0_0_a2_0[11]\ : OR2FT
      port map(A => REG_54, B => N_1574_0, Y => N_1474);
    
    \FID[29]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_199\, CLR => CLEAR_14, Q
         => \FID[29]_net_1\);
    
    CRC32_124 : MUX2H
      port map(A => \CRC32[31]_net_1\, B => N_1222, S => N_1469_0, 
        Y => \CRC32_124\);
    
    \BNC_CNT[11]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_227\, CLR => 
        CLEAR_2, Q => \BNC_CNT[11]_net_1\);
    
    \EVENT_DWORD_17_i_0[9]\ : OAI21TTF
      port map(A => \EVENT_DWORD[17]_net_1\, B => N_105_i_0_1, C
         => N_294, Y => \EVENT_DWORD_17_i_0[9]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I9_S_0 : XOR2FT
      port map(A => \REG[41]\, B => \un2_evread_1[14]\, Y => 
        ADD_16x16_slow_I9_S_0);
    
    \BNC_CNT[25]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_241\, CLR => 
        CLEAR_3, Q => \BNC_CNT[25]_net_1\);
    
    un2_bnc_cnt_I_132 : AND3
      port map(A => \BNC_CNT[18]_net_1\, B => \BNC_CNT[19]_net_1\, 
        C => \BNC_CNT[20]_net_1\, Y => \DWACT_FINC_E[15]\);
    
    un1_REG_1_ADD_16x16_slow_I13_S : XOR2
      port map(A => I12_un1_CO1, B => ADD_16x16_slow_I13_S_0, Y
         => ADD_16x16_slow_I13_S);
    
    un4_bnc_res_9 : XOR2
      port map(A => \BNC_CNT[9]_net_1\, B => REG_413, Y => 
        un4_bnc_res_9_i_i);
    
    \OR_RADDR_3_i_0[1]\ : AND2
      port map(A => N_532_3_3, B => \CNT_0[1]_net_1\, Y => N_687);
    
    un1_REG_1_G : NOR2
      port map(A => ADD_16x16_slow_I5_CO1_0_a0_0, B => 
        un5_evread_7, Y => ADD_16x16_slow_I5_CO1_0_a0_3);
    
    \STATE1_ns_1_iv_0_0_o3_2[0]\ : OAI21FTT
      port map(A => \STATE1_ns_1_iv_0_0_a3_0_1[0]_net_1\, B => 
        N_221, C => \STATE1_ns_1_iv_0_0_o3_0[0]_net_1\, Y => 
        \STATE1_ns_1_iv_0_0_o3_2_i[0]\);
    
    BNC_CNT_239 : MUX2H
      port map(A => \BNC_CNT[23]_net_1\, B => 
        \BNC_CNT_3[23]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_239\);
    
    un4_bnc_res_NE_20 : OR3
      port map(A => un4_bnc_res_NE_13_i, B => un4_bnc_res_28_i_i, 
        C => un4_bnc_res_11_i_i, Y => un4_bnc_res_NE_20_i);
    
    \PDL_RADDR[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RADDR_214\, CLR => 
        CLEAR_17, Q => \PDL_RADDR[4]_net_1\);
    
    N_161_i_0_a2_0_i_o2 : NAND2
      port map(A => \STATE1[0]_net_1\, B => \STATE1[3]_net_1\, Y
         => N_195);
    
    un1_REG_1_ADD_16x16_slow_I8_S : XOR2
      port map(A => N220, B => ADD_16x16_slow_I8_S_0, Y => 
        ADD_16x16_slow_I8_S);
    
    \EVENT_DWORD_17_i_0_a2_0[28]\ : NOR2
      port map(A => I2C_RDATA(8), B => N_1768_i, Y => N_1695);
    
    STATE1_tr16_1_0_a2_0_a2_0_a2_0_a2 : OR2FT
      port map(A => N_1573, B => N_221, Y => N_620_4);
    
    \CRC32_2_i_0[18]\ : NOR2FT
      port map(A => N_532_3_1, B => N_285_i_i_0, Y => N_1382);
    
    \FID_6_iv_0_0_a2_0[22]\ : OR2FT
      port map(A => REG_65, B => N_1574_1, Y => N_1513);
    
    L2AF3 : DFFC
      port map(CLK => ALICLK_c, D => \L2AF2\, CLR => HWRES_c_12, 
        Q => \L2AF3\);
    
    \EVENT_DWORD_17_i_0_a2_0[7]\ : NOR2
      port map(A => \EVENT_DWORD[7]_net_1\, B => N_1229_i, Y => 
        N_1621);
    
    \CRC32_2_i_0_x2[1]\ : XOR2FT
      port map(A => \CRC32[1]_net_1\, B => \EVENT_DWORD[1]_net_1\, 
        Y => N_277_i_i_0);
    
    \FID_2_0[8]\ : XOR2
      port map(A => \CRC32[16]_net_1\, B => \CRC32[28]_net_1\, Y
         => \FID_2_0[8]_net_1\);
    
    \CRC32_2_i_0[28]\ : NOR2FT
      port map(A => N_532_3_2, B => N_264_i_i_0, Y => N_1385);
    
    un1_evread_1 : OR2FT
      port map(A => EVREAD, B => \FIFO_END_EVNT\, Y => 
        \un2_evread_1[14]\);
    
    un2_bnc_cnt_I_91 : XOR2
      port map(A => N_98_0, B => \BNC_CNT[15]_net_1\, Y => I_91_0);
    
    \un2_i2c_chain_0_i_0_a2_5[2]\ : OR2
      port map(A => \CNT_0[3]_net_1\, B => \CNT[5]_net_1\, Y => 
        N_1774);
    
    EVNT_NUM_2_I_43 : XOR2
      port map(A => \EVNT_NUM[8]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_3[0]\, Y => \EVNT_NUM_2[8]\);
    
    \CRC32_2_i_0_x2[25]\ : XOR2FT
      port map(A => \CRC32[25]_net_1\, B => 
        \EVENT_DWORD[25]_net_1\, Y => N_1780_i_0);
    
    CHANNEL_131 : MUX2H
      port map(A => \CHANNEL[1]_net_1\, B => N_98, S => 
        I2C_RREQ_1_sqmuxa, Y => \CHANNEL_131\);
    
    EVNT_NUM_2_I_55 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11[0]\, B => 
        \EVNT_NUM[6]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    \EVENT_DWORD[30]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_168\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[30]_net_1\);
    
    \un2_i2c_chain_0_i_0_o2[2]\ : OR2FT
      port map(A => \CNT[4]_net_1\, B => \CNT_0[1]_net_1\, Y => 
        N_186);
    
    L2RS_1 : OR3
      port map(A => \L2RF1\, B => \L2RF2\, C => \L2RF3\, Y => 
        \L2RS_1\);
    
    \CHIP_ADDR[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \CHIP_ADDR_134\, CLR => 
        CLEAR_5, Q => \CHIP_ADDR[1]_net_1\);
    
    CYC_STAT_1_2 : NOR2FT
      port map(A => \CYC_STAT_0\, B => \CLEAR_PSM_FLAGS\, Y => 
        \CYC_STAT_1_2\);
    
    \RDY_CNT_8_i_0_a2_0[0]\ : NOR2
      port map(A => N_222, B => N_234, Y => N_1583);
    
    \BNC_CNT[4]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_220\, CLR => 
        CLEAR_4, Q => \BNC_CNT[4]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I11_S_0 : XOR2FT
      port map(A => \REG[43]\, B => \un2_evread_1[14]\, Y => 
        ADD_16x16_slow_I11_S_0);
    
    \EVENT_DWORD_17_r[14]\ : AND3FFT
      port map(A => N_1657, B => \EVENT_DWORD_17_i_0_0[14]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[14]\);
    
    \EVENT_DWORD_17_i_a2_0[9]\ : NOR2
      port map(A => \EVENT_DWORD[9]_net_1\, B => N_1229_i, Y => 
        N_295);
    
    \STATE2[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE2_ns_i_i_a2_i[1]_net_1\, 
        CLR => CLEAR_20, Q => \STATE2[1]_net_1\);
    
    \un2_i2c_chain_0_i_0_1[2]\ : OA21FTT
      port map(A => N_189, B => N_1766, C => N_300, Y => 
        \un2_i2c_chain_0_i_0_1[2]_net_1\);
    
    \STATE1_ns_i_0_2[1]\ : OA21FTT
      port map(A => N_242, B => N_252, C => 
        \STATE1_ns_i_0_1[1]_net_1\, Y => 
        \STATE1_ns_i_0_2[1]_net_1\);
    
    \REG_1[43]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I11_S, CLR => 
        CLEAR_19, Q => \REG[43]\);
    
    un2_bnc_cnt_I_216 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \DWACT_FINC_E[26]\, Y => N_9);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m7 : AND3FFT
      port map(A => ADD_16x16_slow_I14_un1_CO1_m7_4_i, B => 
        ADD_16x16_slow_I14_un1_CO1_m7_3_i, C => I6_un1_CO1_i_0_i, 
        Y => ADD_16x16_slow_I14_un1_CO1_N_17);
    
    OR_RADDR_208 : MUX2H
      port map(A => \OR_RADDR[4]_net_1\, B => N_681, S => N_248, 
        Y => \OR_RADDR_208\);
    
    EVNT_NUM_2_I_41 : XOR2
      port map(A => \EVNT_NUM[7]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => \EVNT_NUM_2[7]\);
    
    \EVENT_DWORD_17_i_0_1[22]\ : OAI21FTF
      port map(A => N_1454_0, B => OR_RDATA(2), C => 
        \EVENT_DWORD_17_i_0_0[22]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[22]_net_1\);
    
    EVENT_DWORD_163 : MUX2H
      port map(A => \EVENT_DWORD[25]_net_1\, B => 
        \EVENT_DWORD_17[25]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_163\);
    
    un1_REG_1_ADD_16x16_slow_I13_CO1_1 : OAI21FTF
      port map(A => ADD_16x16_slow_I13_CO1_0_a0_5, B => 
        I7_un3_CO1, C => \un2_evread[14]\, Y => 
        ADD_16x16_slow_I13_CO1_0);
    
    \CRC32_2_i_0_x2[18]\ : XOR2FT
      port map(A => \CRC32[18]_net_1\, B => 
        \EVENT_DWORD[18]_net_1\, Y => N_285_i_i_0);
    
    \CRC32[27]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_120\, CLR => CLEAR_7, 
        Q => \CRC32[27]_net_1\);
    
    \FID_6_iv_0_0_0[14]\ : OAI21
      port map(A => N_1575_0, B => N_270_i_0_i, C => N_1510, Y
         => \FID_6_iv_0_0_0_i[14]\);
    
    \EVENT_DWORD_17_i_0_0[6]\ : OAI21TTF
      port map(A => \EVENT_DWORD[14]_net_1\, B => N_105_i_0, C
         => N_1649, Y => \EVENT_DWORD_17_i_0_0[6]_net_1\);
    
    un2_bnc_cnt_I_156 : XOR2
      port map(A => N_52, B => \BNC_CNT[23]_net_1\, Y => I_156);
    
    \FID_6_iv_0_x2[15]\ : XOR2FT
      port map(A => \CRC32[11]_net_1\, B => \CRC32[23]_net_1\, Y
         => N_57_i_0_i);
    
    un1_STATE1_19_i_i_a2 : NOR2FT
      port map(A => N_1585, B => \STATE1_0[1]_net_1\, Y => N_1587);
    
    \EVNT_TRG\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_TRG_125\, CLR => 
        CLEAR_12, Q => EVNT_TRG_net_1);
    
    \EVENT_DWORD_17_i_0_a2_0[18]\ : NOR2
      port map(A => \EVENT_DWORD[28]_net_1\, B => N_190_i_0, Y
         => N_1667);
    
    \EVENT_DWORD_17_i_0_a2[17]\ : NOR2
      port map(A => \EVENT_DWORD[27]_net_1\, B => N_190_i_0, Y
         => N_291);
    
    un4_bnc_res_30 : XOR2
      port map(A => \BNC_CNT[30]_net_1\, B => REG_434, Y => 
        un4_bnc_res_30_i_i);
    
    un1_REG_1_ADD_16x16_slow_I4_un1_CO1_1 : OAI21TTF
      port map(A => ADD_16x16_slow_I4_un1_CO1_0_a0_0_0_i, B => 
        ADD_16x16_slow_I4_un1_CO1_0_a0_1_i, C => 
        ADD_16x16_slow_I3_CO1_1_0_i_i, Y => 
        ADD_16x16_slow_I4_un1_CO1_0);
    
    \un2_i2c_chain_0_i_0_0[2]\ : AOI21TTF
      port map(A => \CNT[4]_net_1\, B => N_1629_1, C => N_1774, Y
         => \un2_i2c_chain_0_i_0_0[2]_net_1\);
    
    CRC32_104 : MUX2H
      port map(A => \CRC32[11]_net_1\, B => N_1218, S => N_1469_1, 
        Y => \CRC32_104\);
    
    WRB_129 : MUX2H
      port map(A => N_182, B => \WRB\, S => N_697, Y => \WRB_129\);
    
    \STATE1_d_i[7]\ : INV
      port map(A => \STATE1_d[7]\, Y => \STATE1_d_i[7]_net_1\);
    
    \CRC32_2_i_0_x2[24]\ : XOR2FT
      port map(A => \CRC32[24]_net_1\, B => 
        \EVENT_DWORD[24]_net_1\, Y => N_279_i_i_0);
    
    BNC_LIMIT : DFFC
      port map(CLK => ALICLK_c, D => \BNC_LIMIT_2\, CLR => 
        CLEAR_5, Q => \BNC_LIMIT\);
    
    \EVENT_DWORD_17_i_0_0[2]\ : OAI21TTF
      port map(A => \EVENT_DWORD[10]_net_1\, B => N_105_i_0, C
         => N_1645, Y => \EVENT_DWORD_17_i_0_0[2]_net_1\);
    
    EVENT_DWORD_145 : MUX2H
      port map(A => \EVENT_DWORD[7]_net_1\, B => 
        \EVENT_DWORD_17[7]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_145\);
    
    FID_199 : MUX2H
      port map(A => \FID[29]_net_1\, B => \FID_6[29]\, S => 
        N_205_0, Y => \FID_199\);
    
    \EVENT_DWORD[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_151\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[13]_net_1\);
    
    \STATE1_ns_1_iv_0_0_a2_0[0]\ : AO21FTT
      port map(A => \READ_PDL_FLAG\, B => \READ_OR_FLAG\, C => 
        \READ_ADC_FLAG\, Y => \STATE1_ns_1_iv_0_0_a2_0[0]_net_1\);
    
    \CRC32[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_96\, CLR => CLEAR_8, Q
         => \CRC32[3]_net_1\);
    
    \BNC_CNT_3[18]\ : AND2
      port map(A => I_115, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[18]_net_1\);
    
    \un2_i2c_chain_0_i_0_a2_1[2]\ : NAND2
      port map(A => N_186, B => N_1773, Y => N_300);
    
    \un2_i2c_chain_0_0_0_a2_0[1]\ : AND3
      port map(A => N_218, B => \CNT[0]_net_1\, C => 
        \CNT[4]_net_1\, Y => N_1630_i);
    
    un2_bnc_cnt_I_101 : AND2
      port map(A => \BNC_CNT[15]_net_1\, B => \BNC_CNT[16]_net_1\, 
        Y => \DWACT_FINC_E[11]\);
    
    \FID_6_r[11]\ : OA21
      port map(A => N_1475_i, B => \FID_6_iv_0_0_0_i[11]\, C => 
        N_532_3_5, Y => \FID_6[11]\);
    
    \CRC32_2_i_0[4]\ : NOR2FT
      port map(A => N_532_3_0, B => N_274_i_i_0, Y => N_1216);
    
    \EVENT_DWORD_17_i_a2[27]\ : NOR2
      port map(A => I2C_RDATA(7), B => N_1768_i, Y => N_1678);
    
    \CRC32[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_102\, CLR => CLEAR_8, 
        Q => \CRC32[9]_net_1\);
    
    \CNT_8_i[2]\ : AND2
      port map(A => N_185_i, B => I_22_0, Y => N_78);
    
    \REG_1[20]\ : DFFC
      port map(CLK => CLK_c_c, D => \REG_1_20_127_i_a2\, CLR => 
        CLEAR_18, Q => \REG[20]\);
    
    G : OR2
      port map(A => \REG[34]\, B => \REG[35]\, Y => un5_evread_7);
    
    FAULT_STROBE : DFFC
      port map(CLK => CLK_c_c, D => \FAULT_STROBE_2\, CLR => 
        HWRES_c_11, Q => \FAULT_STROBE\);
    
    un1_STATE1_2_0_i_a3_i_1 : NAND2
      port map(A => N_532_3_0, B => N_620_4_0, Y => N_1469_1);
    
    \STATE1_ns_0_0_0_a2_1_1[3]\ : NOR2
      port map(A => \READ_ADC_FLAG\, B => \READ_PDL_FLAG\, Y => 
        N_1733_1);
    
    \EVENT_DWORD[28]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_166\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[28]_net_1\);
    
    un4_bnc_res_NE_22 : OR3
      port map(A => un4_bnc_res_NE_9_i, B => un4_bnc_res_18_i_i, 
        C => un4_bnc_res_21_i_i, Y => un4_bnc_res_NE_22_i);
    
    \FID_6_r[17]\ : OA21
      port map(A => N_1555_i, B => \FID_6_iv_0_0_1_i[17]\, C => 
        N_532_3_5, Y => \FID_6[17]\);
    
    \EVENT_DWORD_17_i_o2_1_o3[7]\ : OA21
      port map(A => I2C_RACK, B => \STATE1[3]_net_1\, C => N_1753, 
        Y => N_180);
    
    \EVENT_DWORD[19]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_157\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[19]_net_1\);
    
    \CRC32_2_i_0_x2[2]\ : XOR2FT
      port map(A => \CRC32[2]_net_1\, B => \EVENT_DWORD[2]_net_1\, 
        Y => N_261_i_i_0);
    
    un1_REG_1_ADD_16x16_slow_I0_S : XOR2FT
      port map(A => \REG[32]\, B => \un2_evread[15]_net_1\, Y => 
        ADD_16x16_slow_I0_S);
    
    I2C_RREQ_1_sqmuxa_0_a5_0_a2_i : INV
      port map(A => N_215, Y => N_215_i_0);
    
    FAULT_STAT_1_sqmuxa : OA21TTF
      port map(A => \FAULT_STROBE\, B => FAULT_STROBE_0_i, C => 
        \CLEAR_PSM_FLAGS\, Y => \FAULT_STAT_1_sqmuxa\);
    
    EVNT_NUM_2_I_65 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_0[0]\, B => 
        \EVNT_NUM[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    un1_REG_1_ADD_16x16_slow_I7_S : XOR2
      port map(A => I6_un1_CO1_i_0_i, B => ADD_16x16_slow_I7_S_0, 
        Y => ADD_16x16_slow_I7_S);
    
    un1_REG_1_ADD_16x16_slow_I4_un1_CO1_0_a0_0 : OR2
      port map(A => \REG[32]\, B => \REG[34]\, Y => 
        ADD_16x16_slow_I4_un1_CO1_0_a0_0_0_i);
    
    \FID_6_r[9]\ : AND3FFT
      port map(A => N_1528, B => \FID_6_iv_0_0_0[9]_net_1\, C => 
        N_532_3_5, Y => \FID_6[9]\);
    
    \FID[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_178\, CLR => CLEAR_15, Q
         => \FID[8]_net_1\);
    
    \FID_6_r[24]\ : OA21
      port map(A => N_1490_i, B => \FID_6_iv_0_0_0_i[24]\, C => 
        N_532_3_4, Y => \FID_6[24]\);
    
    un2_bnc_cnt_I_5 : XOR2
      port map(A => \BNC_CNT[0]_net_1\, B => \BNC_CNT[1]_net_1\, 
        Y => I_5_2);
    
    un1_ORATETMO_1_I_21 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12_5[0]\, Y => I_21);
    
    un2_bnc_cnt_I_83 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[7]\, C
         => \DWACT_FINC_E[8]\, Y => N_103);
    
    \REG_1[44]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I12_S, CLR => 
        CLEAR_19, Q => \REG[44]\);
    
    \un2_i2c_chain_0_0_0_0_0[5]\ : AO21FTF
      port map(A => N_265_i_i_0_i, B => N_1764, C => 
        \un2_i2c_chain_0_0_0_a2_11[5]_net_1\, Y => 
        \un2_i2c_chain_0_0_0_0_0_i[5]\);
    
    \CRC32_2_i_0_a2_s_0[17]\ : NOR2
      port map(A => \STATE1[0]_net_1\, B => \STATE1[3]_net_1\, Y
         => N_1585_0);
    
    \CNT_0[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_8_i[1]_net_1\, CLR => 
        CLEAR_0, Q => \CNT_0[1]_net_1\);
    
    \STATE1_ns_i_0_a2_1[1]\ : NAND2
      port map(A => N_222, B => N_1454, Y => N_1564);
    
    \EVENT_DWORD_17_i_0_a2_0[1]\ : NOR2
      port map(A => \EVENT_DWORD[1]_net_1\, B => N_1229_i, Y => 
        N_330);
    
    STATE1_s10_i_o3_i_o4_i_a2_0_i2_i_o2 : OR2FT
      port map(A => \STATE1_0[3]_net_1\, B => \STATE1_0[0]_net_1\, 
        Y => N_221);
    
    un1_REG_1_ADD_16x16_slow_I3_CO1_1 : OAI21FTF
      port map(A => ADD_16x16_slow_I3_CO1_0_a0_1, B => 
        un5_evread_7, C => ADD_16x16_slow_I3_CO1_1_0_i_i, Y => 
        ADD_16x16_slow_I3_CO1_0);
    
    \STATE1_ns_1_iv_0_0_7[2]\ : AND3FFT
      port map(A => N_1559_i, B => \STATE1_ns_1_iv_0_0_5_i[2]\, C
         => N_520, Y => \STATE1_ns_1_iv_0_0_7[2]_net_1\);
    
    \CRC32_2_i_0[1]\ : NOR2FT
      port map(A => N_532_3_0, B => N_277_i_i_0, Y => N_1288);
    
    \FID_2[6]\ : XOR2FT
      port map(A => \CRC32[2]_net_1\, B => \FID_2_0[6]_net_1\, Y
         => \FID_2_i[6]\);
    
    \RDY_CNT_8_i_0[1]\ : AND2
      port map(A => N_267, B => I_10, Y => 
        \RDY_CNT_8_i_0[1]_net_1\);
    
    L1AF1 : DFFC
      port map(CLK => ALICLK_c, D => L1A_c_c, CLR => HWRES_c_11, 
        Q => \L1AF1\);
    
    un1_ORATETMO_1_I_7 : AND2
      port map(A => \ORATETMO_i_i[3]\, B => N_701_i_0, Y => 
        \DWACT_ADD_CI_0_g_array_0_3[0]\);
    
    \STATE1_ns_1_iv_0_0_m2[0]\ : MUX2H
      port map(A => N_1778, B => N_1777, S => \STATE1[2]_net_1\, 
        Y => N_1614);
    
    \FID_6_iv_0_a2_0[27]\ : OR2FT
      port map(A => REG_70, B => N_1574, Y => N_1543);
    
    \FID_6_iv_0_0_a2_1[20]\ : NOR2FT
      port map(A => \EVENT_DWORD[20]_net_1\, B => N_620_4_1, Y
         => N_1481_i);
    
    \FID_6_0_iv_0_a2[29]\ : NOR2FT
      port map(A => REG_72, B => N_1574, Y => N_1545_i);
    
    FID_182 : MUX2H
      port map(A => \FID[12]_net_1\, B => \FID_6[12]\, S => 
        N_205_1, Y => \FID_182\);
    
    EVENT_DWORD_153 : MUX2H
      port map(A => \EVENT_DWORD[15]_net_1\, B => 
        \EVENT_DWORD_17[15]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_153\);
    
    \FID_6_0_iv_0_0_0[2]\ : OAI21FTT
      port map(A => REG_45, B => N_1574_0, C => N_1519, Y => 
        \FID_6_0_iv_0_0_0_i[2]\);
    
    un2_bnc_cnt_I_20 : XOR2
      port map(A => N_149, B => \BNC_CNT[4]_net_1\, Y => I_20_1);
    
    \FID_6_0_iv_0_0_0[1]\ : OAI21FTT
      port map(A => REG_44, B => N_1574_0, C => N_1505, Y => 
        \FID_6_0_iv_0_0_0_i[1]\);
    
    \STATE1_ns_1_iv_0_1_o2_3_o3[0]\ : NOR3
      port map(A => N_1744, B => N_1746, C => 
        \STATE1_ns_1_iv_0_1_o2_3_o3_0[0]_net_1\, Y => N_1777);
    
    \FID_6_iv_0_0_a2_1_0_a2[28]\ : OR2FT
      port map(A => \STATE1[1]_net_1\, B => N_195, Y => N_1575);
    
    un2_bnc_cnt_I_169 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        C => \BNC_CNT[24]_net_1\, Y => \DWACT_FINC_E[19]\);
    
    un2_bnc_cnt_I_111 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \DWACT_FINC_E[5]\, Y => \DWACT_FINC_E[28]\);
    
    un1_REG_1_ADD_16x16_slow_I9_S : XOR2
      port map(A => I8_un1_CO1, B => ADD_16x16_slow_I9_S_0, Y => 
        ADD_16x16_slow_I9_S);
    
    \BNC_CNT_3[23]\ : AND2
      port map(A => I_156, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[23]_net_1\);
    
    \FID_6_iv_0_0_0[23]\ : OAI21FTT
      port map(A => \EVNT_NUM[7]_net_1\, B => N_1575_1, C => 
        N_1486, Y => \FID_6_iv_0_0_0_i[23]\);
    
    EVNT_NUM_2_I_1 : AND2
      port map(A => \EVNT_NUM[0]_net_1\, B => N_161_i_0, Y => 
        \DWACT_ADD_CI_0_TMP_0[0]\);
    
    un2_bnc_cnt_I_129 : XOR2
      port map(A => N_71, B => \BNC_CNT[20]_net_1\, Y => I_129);
    
    \FID_6_iv_0_0_a2_0[13]\ : OR2FT
      port map(A => REG_56, B => N_1574_1, Y => N_1530);
    
    \EVENT_DWORD[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_147\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[9]_net_1\);
    
    un2_bnc_cnt_I_121 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \BNC_CNT[18]_net_1\, Y => N_76);
    
    \STATE1_ns_1_iv_0_0_2[2]\ : OAI21TTF
      port map(A => N_1586, B => N_1733_1, C => N_1558_i, Y => 
        \STATE1_ns_1_iv_0_0_2_i[2]\);
    
    un2_bnc_cnt_I_173 : XOR2
      port map(A => N_40, B => \BNC_CNT[25]_net_1\, Y => I_173);
    
    BNC_CNT_238 : MUX2H
      port map(A => \BNC_CNT[22]_net_1\, B => 
        \BNC_CNT_3[22]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_238\);
    
    \EVENT_DWORD_17_i_0_a2_0[25]\ : NOR2
      port map(A => \EVENT_DWORD[25]_net_1\, B => N_1229_i_0, Y
         => N_1737);
    
    \EVENT_DWORD_17_r[16]\ : AND3FFT
      port map(A => N_1660, B => \EVENT_DWORD_17_i_0_0[16]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[16]\);
    
    \un2_i2c_chain_0_0_0_a2_11[5]\ : OR3FTT
      port map(A => \CNT_0[3]_net_1\, B => N_1763, C => N_216, Y
         => \un2_i2c_chain_0_0_0_a2_11[5]_net_1\);
    
    \STATE1_ns_1_iv_0_0_a2_1[2]\ : NOR3FFT
      port map(A => N_222, B => N_215_i_0, C => N_120_i, Y => 
        N_1558_i);
    
    \EVENT_DWORD_17_i_o2_1_o2_0[7]\ : OA21FTF
      port map(A => \STATE1_0[0]_net_1\, B => N_180, C => 
        N_1755_i, Y => N_1229_i_0);
    
    BNC_CNT_237 : MUX2H
      port map(A => \BNC_CNT[21]_net_1\, B => 
        \BNC_CNT_3[21]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_237\);
    
    BNC_CNT_236 : MUX2H
      port map(A => \BNC_CNT[20]_net_1\, B => 
        \BNC_CNT_3[20]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_236\);
    
    un1_STATE1_19_i_i_a2_0 : OR2FT
      port map(A => PULSE(3), B => N_1574_0, Y => N_522);
    
    un1_REG_1_ADD_16x16_slow_I5_S_0 : XOR2FT
      port map(A => \REG[37]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I5_S_0);
    
    \EVENT_DWORD_17_i_0_a2[15]\ : NOR2
      port map(A => \EVENT_DWORD[25]_net_1\, B => N_190_i_0, Y
         => N_1623);
    
    \FID_6_0_iv_0_a2_2_0_a2_1[3]\ : OR2
      port map(A => \STATE1_0[3]_net_1\, B => N_176_0, Y => 
        N_1574_1);
    
    \EVENT_DWORD[17]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_155\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[17]_net_1\);
    
    \EVENT_DWORD_17_r[17]\ : AND3FFT
      port map(A => N_292, B => \EVENT_DWORD_17_i_0_0[17]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[17]\);
    
    EVENT_DWORD_161 : MUX2H
      port map(A => \EVENT_DWORD[23]_net_1\, B => 
        \EVENT_DWORD_17[23]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_161\);
    
    \CRC32[18]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_111\, CLR => CLEAR_7, 
        Q => \CRC32[18]_net_1\);
    
    BNC_CNT_223 : MUX2H
      port map(A => \BNC_CNT[7]_net_1\, B => \BNC_CNT_3[7]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_223\);
    
    un4_bnc_res_5 : XOR2
      port map(A => \BNC_CNT[5]_net_1\, B => REG_409, Y => 
        un4_bnc_res_5_i_i);
    
    ORATETMO_1_sqmuxa_i_0_o2_i : INV
      port map(A => N_252, Y => N_252_i_0);
    
    \BNC_CNT[18]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_234\, CLR => 
        CLEAR_3, Q => \BNC_CNT[18]_net_1\);
    
    un1_STATE1_18_0_0_0 : NAND3FTT
      port map(A => N_1673_i, B => N_1672, C => N_1762, Y => 
        un1_STATE1_18_0);
    
    un2_bnc_cnt_I_97 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[10]\, C
         => \BNC_CNT[15]_net_1\, Y => N_93_0);
    
    WRB : DFFS
      port map(CLK => CLK_c_c, D => \WRB_129\, SET => CLEAR_20, Q
         => \WRB\);
    
    un1_REG_1_ADD_16x16_slow_I8_un1_CO1_0 : OAI21TTF
      port map(A => ADD_16x16_slow_I8_un1_CO1_0_tz_0, B => 
        I7_un3_CO1, C => \un2_evread_1[14]\, Y => 
        ADD_16x16_slow_I8_un1_CO1_0);
    
    un1_REG_1_ADD_16x16_slow_I12_S_0 : XOR2FT
      port map(A => \REG[44]\, B => \un2_evread_1[14]\, Y => 
        ADD_16x16_slow_I12_S_0);
    
    \CRC32_2_i_0[14]\ : NOR2FT
      port map(A => N_532_3_1, B => N_257_i_i_0, Y => N_1291);
    
    un1_REG_1_ADD_16x16_slow_I2_un1_CO1_1 : OAI21FTF
      port map(A => ADD_16x16_slow_I2_un1_CO1_0_a0_0, B => 
        \REG[33]\, C => ADD_16x16_slow_I3_CO1_1_0_i_i, Y => 
        ADD_16x16_slow_I2_un1_CO1_0);
    
    FID_197 : MUX2H
      port map(A => \FID[27]_net_1\, B => \FID_6[27]\, S => 
        N_205_0, Y => \FID_197\);
    
    \CRC32_2_i_0[24]\ : NOR2FT
      port map(A => N_532_3_2, B => N_279_i_i_0, Y => N_1293);
    
    \CRC32_2_i_0_a2_8[17]\ : OR2FT
      port map(A => N_1585_0, B => N_176_0, Y => N_532_3_8);
    
    \STATE1_ns_1_iv_0_0_1[2]\ : OA21FTT
      port map(A => N_166, B => N_195, C => 
        \STATE1_ns_1_iv_0_0_0[2]_net_1\, Y => 
        \STATE1_ns_1_iv_0_0_1[2]_net_1\);
    
    \FID[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_186\, CLR => CLEAR_13, Q
         => \FID[16]_net_1\);
    
    un4_bnc_res_17 : XOR2
      port map(A => \BNC_CNT[17]_net_1\, B => REG_421, Y => 
        un4_bnc_res_17_i_i);
    
    \BNC_CNT[6]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_222\, CLR => 
        CLEAR_4, Q => \BNC_CNT[6]_net_1\);
    
    \BNC_CNT_3[8]\ : AND2
      port map(A => I_45_0, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[8]_net_1\);
    
    \CRC32_2_i_0_x2[3]\ : XOR2FT
      port map(A => \CRC32[3]_net_1\, B => \EVENT_DWORD[3]_net_1\, 
        Y => N_272_i_i_0);
    
    un1_RDY_CNT_I_8 : XOR2
      port map(A => \RDY_CNT[0]_net_1\, B => 
        \un1_EVENT_DWORD_0_sqmuxa_0_0\, Y => 
        \DWACT_ADD_CI_0_partial_sum_0[0]\);
    
    \FID_6_0_iv_0_a2_0[29]\ : NOR2FT
      port map(A => \EVENT_DWORD[29]_net_1\, B => N_620_4, Y => 
        N_1546_i);
    
    \STATE1_ns_i_0[1]\ : OR3
      port map(A => N_1569_i, B => \STATE1_ns_i_0_5_i[1]\, C => 
        N_7189_i, Y => \STATE1_ns_i_0[1]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2_0[15]\ : NOR2
      port map(A => \EVENT_DWORD[15]_net_1\, B => N_1229_i_1, Y
         => N_1624);
    
    \EVENT_DWORD_17_i_0_0[3]\ : OAI21TTF
      port map(A => \EVENT_DWORD[11]_net_1\, B => N_105_i_0, C
         => N_1616, Y => \EVENT_DWORD_17_i_0_0[3]_net_1\);
    
    \FID_2[10]\ : XOR2FT
      port map(A => \CRC32[6]_net_1\, B => \FID_2_0[10]_net_1\, Y
         => \FID_2_i[10]\);
    
    \un2_i2c_chain_0_i_0_3[2]\ : AO21TTF
      port map(A => N_202_i_i_0, B => N_312_1, C => 
        \un2_i2c_chain_0_i_0_1[2]_net_1\, Y => 
        \un2_i2c_chain_0_i_0_3_i[2]\);
    
    \EVENT_DWORD_17_i_0_0[13]\ : OAI21TTF
      port map(A => \EVENT_DWORD[21]_net_1\, B => N_105_i_0_1, C
         => N_338, Y => \EVENT_DWORD_17_i_0_0[13]_net_1\);
    
    un2_bnc_cnt_I_202 : AND3
      port map(A => \DWACT_FINC_E[24]\, B => \DWACT_FINC_E[23]\, 
        C => \BNC_CNT[27]_net_1\, Y => N_19_0);
    
    \STATE1_ns_i_0_a2[1]\ : NOR2FT
      port map(A => N_289, B => N_215, Y => N_1562_i);
    
    \FID_6_r[6]\ : OA21
      port map(A => N_317_i, B => \FID_6_iv_0_0_0_i[6]\, C => 
        N_532_3_5, Y => \FID_6[6]\);
    
    \FID_6_iv_0_0_a2_1_0_a2_1[28]\ : OR2FT
      port map(A => \STATE1_0[1]_net_1\, B => N_195, Y => 
        N_1575_1);
    
    \STATE1_ns_1_iv_0_0_a2_0[2]\ : OR3FFT
      port map(A => \STATE1[0]_net_1\, B => N_166, C => N_1470, Y
         => N_1557);
    
    \PDL_RADDR[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \PDL_RADDR_211\, CLR => 
        CLEAR_17, Q => \PDL_RADDR[1]_net_1\);
    
    \un2_i2c_chain_0_0_0[6]\ : OR3
      port map(A => \un2_i2c_chain_0_0_0_0_i[6]\, B => N_1637_i, 
        C => N_1639_i, Y => N_99);
    
    \CRC32_2_i_0_x2[30]\ : XOR2FT
      port map(A => \CRC32[30]_net_1\, B => 
        \EVENT_DWORD[30]_net_1\, Y => N_260_i_i_0);
    
    \un2_i2c_chain_0_0_0_2[3]\ : NAND3
      port map(A => N_1633, B => 
        \un2_i2c_chain_0_0_0_a2_4[3]_net_1\, C => N_300, Y => 
        \un2_i2c_chain_0_0_0_2_i[3]\);
    
    \un2_evread_i[14]\ : INV
      port map(A => \un2_evread[14]\, Y => \un2_evread_i_0[14]\);
    
    \FID_6_iv_0_0_a2_0[20]\ : OR2FT
      port map(A => REG_63, B => N_1574_1, Y => N_1480);
    
    \STATE1_ns_0_0_0_i_0[3]\ : OR2
      port map(A => N_215, B => N_289, Y => 
        \STATE1_ns_0_0_0_i_0[3]_net_1\);
    
    \FID_6_r[30]\ : AND3FFT
      port map(A => N_1515, B => N_1516, C => N_532_3_3, Y => 
        \FID_6[30]\);
    
    \BNC_CNT_3[22]\ : AND2
      port map(A => I_143, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[22]_net_1\);
    
    \FID_6_iv_0_0_0[26]\ : OAI21FTT
      port map(A => \EVNT_NUM[10]_net_1\, B => N_1575, C => 
        N_1495, Y => \FID_6_iv_0_0_0_i[26]\);
    
    \FID_6_0_iv_0_0_a2[2]\ : NOR2
      port map(A => GA_c(2), B => N_235, Y => N_1517_i);
    
    EVNT_NUM_2_I_74 : AND2
      port map(A => \EVNT_NUM[8]_net_1\, B => \EVNT_NUM[9]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1_3[0]\);
    
    EVENT_DWORD_167 : MUX2H
      port map(A => \EVENT_DWORD[29]_net_1\, B => 
        \EVENT_DWORD_17[29]\, S => un1_STATE1_18_0, Y => 
        \EVENT_DWORD_167\);
    
    \STATE1_ns_0_0_0_0[3]\ : OAI21FTT
      port map(A => N_207, B => \STATE1_0[2]_net_1\, C => N_1731, 
        Y => \STATE1_ns_0_0_0_0_i[3]\);
    
    un1_STATE1_17_i_0_0 : OR3
      port map(A => N_305, B => N_306, C => N_304, Y => N_697);
    
    \FID[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_171\, CLR => CLEAR_13, Q
         => \FID[1]_net_1\);
    
    CYC_STAT_1_sqmuxa : NOR2
      port map(A => \CLEAR_PSM_FLAGS\, B => \CYC_STAT_1\, Y => 
        \CYC_STAT_1_sqmuxa\);
    
    FID_196 : MUX2H
      port map(A => \FID[26]_net_1\, B => \FID_6[26]\, S => 
        N_205_0, Y => \FID_196\);
    
    \EVNT_NUM[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[5]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[5]_net_1\);
    
    \CRC32_2_i_0[5]\ : NOR2FT
      port map(A => N_532_3_0, B => N_280_i_i_0, Y => N_1376);
    
    \CRC32_2_i_0_x2[12]\ : XOR2FT
      port map(A => \CRC32[12]_net_1\, B => 
        \EVENT_DWORD[12]_net_1\, Y => N_256_i_i_0);
    
    un4_bnc_res_27 : XOR2
      port map(A => \BNC_CNT[27]_net_1\, B => REG_431, Y => 
        un4_bnc_res_27_i_i);
    
    EVENT_DWORD_151 : MUX2H
      port map(A => \EVENT_DWORD[13]_net_1\, B => 
        \EVENT_DWORD_17[13]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_151\);
    
    FID_198 : MUX2H
      port map(A => \FID[28]_net_1\, B => \FID_6[28]\, S => 
        N_205_0, Y => \FID_198\);
    
    un2_bnc_cnt_I_166 : XOR2
      port map(A => N_45, B => \BNC_CNT[24]_net_1\, Y => I_166);
    
    EVENT_DWORD_138 : MUX2H
      port map(A => \EVENT_DWORD[0]_net_1\, B => 
        \EVENT_DWORD_17[0]\, S => un1_STATE1_18, Y => 
        \EVENT_DWORD_138\);
    
    CRC32_118 : MUX2H
      port map(A => \CRC32[25]_net_1\, B => N_1141, S => N_1469_0, 
        Y => \CRC32_118\);
    
    un1_STATE1_18_0_0_a2_0 : OR2
      port map(A => N_195, B => N_176, Y => N_1762);
    
    un2_bnc_cnt_I_16 : AND3
      port map(A => \BNC_CNT[0]_net_1\, B => \BNC_CNT[1]_net_1\, 
        C => \BNC_CNT[2]_net_1\, Y => \DWACT_FINC_E[0]\);
    
    EVNT_NUM_2_I_49 : XOR2
      port map(A => \EVNT_NUM[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => \EVNT_NUM_2[3]\);
    
    un1_REG_1_ADD_16x16_slow_I4_S : XOR2
      port map(A => N212, B => ADD_16x16_slow_I4_S_0, Y => 
        ADD_16x16_slow_I4_S);
    
    \un2_i2c_chain_0_i_0_a3_2[2]\ : OR2FT
      port map(A => \CNT_0[0]_net_1\, B => \CNT_0[1]_net_1\, Y
         => N_1767);
    
    \un2_i2c_chain_0_i_0_o3[2]\ : NOR2FT
      port map(A => \CNT_0[5]_net_1\, B => \CNT_0[0]_net_1\, Y
         => N_189);
    
    un2_bnc_cnt_I_12 : AND3
      port map(A => \BNC_CNT[0]_net_1\, B => \BNC_CNT[1]_net_1\, 
        C => \BNC_CNT[2]_net_1\, Y => N_154);
    
    un1_REG_1_ADD_16x16_slow_I2_un1_CO1 : AO21TTF
      port map(A => N208, B => \REG[34]\, C => 
        ADD_16x16_slow_I2_un1_CO1_0, Y => I2_un1_CO1);
    
    \EVENT_DWORD_17_i_0_0[4]\ : OAI21TTF
      port map(A => \EVENT_DWORD[12]_net_1\, B => N_105_i_0, C
         => N_327, Y => \EVENT_DWORD_17_i_0_0[4]_net_1\);
    
    CRC32_116 : MUX2H
      port map(A => \CRC32[23]_net_1\, B => N_1221, S => N_1469_0, 
        Y => \CRC32_116\);
    
    \BNC_CNT_3[13]\ : AND2
      port map(A => I_77_0, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[13]_net_1\);
    
    \FID_6_r[16]\ : OA21
      port map(A => N_1534_i, B => \FID_6_iv_0_0_0_i[16]\, C => 
        N_532_3_5, Y => \FID_6[16]\);
    
    \FID_2_0[5]\ : XOR2
      port map(A => \CRC32[13]_net_1\, B => \CRC32[25]_net_1\, Y
         => \FID_2_0[5]_net_1\);
    
    \CRC32_2_i_0_x2[28]\ : XOR2FT
      port map(A => \CRC32[28]_net_1\, B => 
        \EVENT_DWORD[28]_net_1\, Y => N_264_i_i_0);
    
    un2_bnc_cnt_I_30 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[1]\, C
         => \BNC_CNT[5]_net_1\, Y => N_141);
    
    \FID_6_0_iv_0_a2_1[3]\ : OR2FT
      port map(A => \EVENT_DWORD[3]_net_1\, B => N_620_4_0, Y => 
        N_311);
    
    \EVENT_DWORD_17_i_a2_0[27]\ : NOR2
      port map(A => \EVENT_DWORD[27]_net_1\, B => N_1229_i_0, Y
         => N_1679);
    
    un1_REG_1_ADD_16x16_slow_I2_S_0 : XOR2FT
      port map(A => \REG[34]\, B => \un2_evread_0[14]\, Y => 
        ADD_16x16_slow_I2_S_0);
    
    \FID_6_r[23]\ : OA21
      port map(A => N_1487_i, B => \FID_6_iv_0_0_0_i[23]\, C => 
        N_532_3_4, Y => \FID_6[23]\);
    
    \EVENT_DWORD_17_i_0_a2[25]\ : NOR2
      port map(A => I2C_RDATA(5), B => N_1768_i, Y => N_1736);
    
    \CRC32_2_i_0_x2[9]\ : XOR2FT
      port map(A => \CRC32[9]_net_1\, B => \EVENT_DWORD[9]_net_1\, 
        Y => N_283_i_i_0);
    
    un1_STATE1_1_sqmuxa_0_0 : NAND2
      port map(A => N_1672, B => STATE1_1_sqmuxa_1, Y => 
        un1_STATE1_1_sqmuxa);
    
    \FID_2[4]\ : XOR2FT
      port map(A => \CRC32[0]_net_1\, B => \FID_2_0[4]_net_1\, Y
         => \FID_2_i[4]\);
    
    un1_evread : OR2FT
      port map(A => EVREAD, B => \FIFO_END_EVNT\, Y => 
        \un2_evread[14]\);
    
    \FID_6_iv_0_0_a2_1[4]\ : NOR2FT
      port map(A => \EVENT_DWORD[4]_net_1\, B => N_620_4_0, Y => 
        N_343_i);
    
    un1_ORATETMO_1_I_26 : AO21
      port map(A => \DWACT_ADD_CI_0_pog_array_0[0]\, B => 
        \DWACT_ADD_CI_0_TMP_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\);
    
    un2_bnc_cnt_I_199 : AND2
      port map(A => \DWACT_FINC_E[29]\, B => \DWACT_FINC_E[30]\, 
        Y => \DWACT_FINC_E[24]\);
    
    un2_bnc_cnt_I_179 : AND3
      port map(A => \DWACT_FINC_E[15]\, B => \DWACT_FINC_E[17]\, 
        C => \DWACT_FINC_E[20]\, Y => \DWACT_FINC_E[21]\);
    
    \CRC32[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_100\, CLR => CLEAR_8, 
        Q => \CRC32[7]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2_0[6]\ : NOR2
      port map(A => \EVENT_DWORD[16]_net_1\, B => N_190_i, Y => 
        N_1649);
    
    \CNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \CNT_8_i[1]_net_1\, CLR => 
        CLEAR_5, Q => \CNT[1]_net_1\);
    
    \BNC_CNT[29]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_245\, CLR => 
        CLEAR_4, Q => \BNC_CNT[29]_net_1\);
    
    \un2_i2c_chain_0_0_0_a2_7[5]\ : OR3FFT
      port map(A => \CNT[4]_net_1\, B => N_1767, C => N_199, Y
         => N_1724);
    
    \FID[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_174\, CLR => CLEAR_15, Q
         => \FID[4]_net_1\);
    
    CYC_STAT_89_i : INV
      port map(A => \CLEAR_PSM_FLAGS\, Y => CLEAR_PSM_FLAGS_i_0);
    
    \un2_i2c_chain_0_0_0_2[4]\ : OAI21TTF
      port map(A => N_1615_i, B => 
        \un2_i2c_chain_0_0_0_a2_0_i[4]\, C => N_1688_i, Y => 
        \un2_i2c_chain_0_0_0_2_i[4]\);
    
    un2_bnc_cnt_I_45 : XOR2
      port map(A => N_131, B => \BNC_CNT[8]_net_1\, Y => I_45_0);
    
    \BNC_CNT_3[20]\ : AND2
      port map(A => I_129, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[20]_net_1\);
    
    \FID_6_iv_0_0_a2_0[15]\ : OR2FT
      port map(A => REG_58, B => N_1574_1, Y => N_1477);
    
    \FID_6_r[29]\ : OA21
      port map(A => N_1545_i, B => N_1546_i, C => N_532_3_4, Y
         => \FID_6[29]\);
    
    BNC_CNT_247 : MUX2H
      port map(A => \BNC_CNT[31]_net_1\, B => 
        \BNC_CNT_3[31]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_247\);
    
    un1_REG_1_G_8_0_a2_2 : NAND3FFT
      port map(A => G_6, B => N_7210_i, C => \REG[38]\, Y => 
        G_8_0_a2_2);
    
    EVNT_NUM_2_I_51 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_0[0]\, B => 
        \EVNT_NUM[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1_0[0]\);
    
    un1_STATE1_17_i_0_i4_0_a2_0_a2_0_i2_0_o2_0 : OR2
      port map(A => \STATE1_0[2]_net_1\, B => \STATE1_0[1]_net_1\, 
        Y => N_176_0);
    
    \EVNT_NUM[0]\ : DFFC
      port map(CLK => CLK_c_c, D => 
        \DWACT_ADD_CI_0_partial_sum_2[0]\, CLR => CLEAR_11, Q => 
        \EVNT_NUM[0]_net_1\);
    
    \BNC_CNT_3[30]\ : AND2
      port map(A => I_217, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[30]_net_1\);
    
    BNC_CNT_246 : MUX2H
      port map(A => \BNC_CNT[30]_net_1\, B => 
        \BNC_CNT_3[30]_net_1\, S => LBSP_c_0(2), Y => 
        \BNC_CNT_246\);
    
    un5_evread_5 : NOR3
      port map(A => \REG[47]\, B => \REG[46]\, C => \REG[39]\, Y
         => \un5_evread_5\);
    
    un1_REG_1_ADD_16x16_slow_I6_un1_CO1_0_a0_0 : NOR2
      port map(A => \REG[38]\, B => \REG[37]\, Y => 
        ADD_16x16_slow_I6_un1_CO1_0_a0_0);
    
    EVENT_DWORD_157 : MUX2H
      port map(A => \EVENT_DWORD[19]_net_1\, B => 
        \EVENT_DWORD_17[19]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_157\);
    
    un1_REG_1_G_6_0_o2 : AO21TTF
      port map(A => N228, B => \REG[44]\, C => 
        ADD_16x16_slow_I12_un1_CO1_0, Y => I12_un1_CO1);
    
    \FID_6_iv_0_0_0[12]\ : OAI21
      port map(A => N_1575_0, B => N_271_i_0_i, C => N_1507, Y
         => \FID_6_iv_0_0_0_i[12]\);
    
    \EVENT_DWORD_17_i_0_a2[5]\ : NOR2
      port map(A => \EVENT_DWORD[15]_net_1\, B => N_190_i, Y => 
        N_332);
    
    un5_evread_1 : OR2FT
      port map(A => \REG[32]\, B => \REG[33]\, Y => 
        \un5_evread_1\);
    
    EVNT_TRG_125 : MUX2H
      port map(A => N_1147, B => EVNT_TRG_net_1, S => 
        \STATE2[2]_net_1\, Y => \EVNT_TRG_125\);
    
    \un2_i2c_chain_0_0_0_0_3[5]\ : OAI21TTF
      port map(A => N_1765, B => 
        \un2_i2c_chain_0_0_0_0_1_tz[5]_net_1\, C => 
        \un2_i2c_chain_0_0_0_1_0_i[5]\, Y => 
        \un2_i2c_chain_0_0_0_0_3_i[5]\);
    
    \CRC32_2_i_0_x2[17]\ : XOR2FT
      port map(A => \CRC32[17]_net_1\, B => 
        \EVENT_DWORD[17]_net_1\, Y => N_1779_i_0);
    
    \CHIP_ADDR[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \CHIP_ADDR_133\, CLR => 
        CLEAR_5, Q => \CHIP_ADDR[0]_net_1\);
    
    un1_REG_1_ADD_16x16_slow_I13_CO1_0_a0_0 : NOR2
      port map(A => \REG[45]\, B => \REG[44]\, Y => 
        ADD_16x16_slow_I13_CO1_0_a0_0);
    
    \un2_i2c_chain_0_0_0_a3[3]\ : NOR2FT
      port map(A => N_189, B => \CNT_0[4]_net_1\, Y => N_1770);
    
    \CRC32_2_i_0_x2[10]\ : XOR2FT
      port map(A => \CRC32[10]_net_1\, B => 
        \EVENT_DWORD[10]_net_1\, Y => N_278_i_i_0);
    
    un5_evread_8 : OR3FTT
      port map(A => \un5_evread_5\, B => \REG[43]\, C => 
        \REG[44]\, Y => un5_evread_8_i);
    
    \EVENT_DWORD[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_150\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[12]_net_1\);
    
    un4_bnc_res_6 : XOR2
      port map(A => \BNC_CNT[6]_net_1\, B => REG_410, Y => 
        un4_bnc_res_6_i_i);
    
    FAULT_STAT_3 : NOR2FT
      port map(A => REG_c(22), B => \CLEAR_PSM_FLAGS\, Y => 
        \FAULT_STAT_3\);
    
    \EVENT_DWORD[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_138\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[0]_net_1\);
    
    un4_bnc_res_NE_1_0 : OR3
      port map(A => un4_bnc_res_NE_29_i, B => un4_bnc_res_NE_25_i, 
        C => un4_bnc_res_NE_24_i, Y => un4_bnc_res_i_1);
    
    un2_bnc_cnt_I_31 : XOR2
      port map(A => N_141, B => \BNC_CNT[6]_net_1\, Y => I_31_0);
    
    \I2C_RREQ\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RREQ_137\, CLR => 
        CLEAR_15, Q => I2C_RREQ_net_1);
    
    CRC32_110 : MUX2H
      port map(A => \CRC32[17]_net_1\, B => N_1140, S => N_1469_1, 
        Y => \CRC32_110\);
    
    \BNC_CNT_3[27]\ : AND2
      port map(A => I_196, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[27]_net_1\);
    
    OR_RACK_sync : DFFC
      port map(CLK => CLK_c_c, D => OR_RACK, CLR => CLEAR_16, Q
         => \OR_RACK_sync\);
    
    un4_bnc_res_NE_11 : OR2
      port map(A => un4_bnc_res_12_i_i, B => un4_bnc_res_15_i_i, 
        Y => un4_bnc_res_NE_11_i);
    
    \EVENT_DWORD_17_i_0_a2_0[21]\ : NOR2
      port map(A => I2C_RDATA(1), B => N_1768_i, Y => N_1719);
    
    \EVENT_DWORD_17_i_0_0[12]\ : OAI21TTF
      port map(A => \EVENT_DWORD[20]_net_1\, B => N_105_i_0_1, C
         => N_1655, Y => \EVENT_DWORD_17_i_0_0[12]_net_1\);
    
    CRC32_108 : MUX2H
      port map(A => \CRC32[15]_net_1\, B => N_1219, S => N_1469_1, 
        Y => \CRC32_108\);
    
    un1_STATE1_24_i_i_o2 : OAI21FTT
      port map(A => N_193, B => \un1_STATE1_24_i_i_a2_1\, C => 
        N_532_3_3, Y => N_248);
    
    \FID_6_r[10]\ : OA21
      port map(A => N_1472_i, B => \FID_6_iv_0_0_0_i[10]\, C => 
        N_532_3_5, Y => \FID_6[10]\);
    
    un4_bnc_res_0 : XOR2
      port map(A => \BNC_CNT[0]_net_1\, B => REG_404, Y => 
        un4_bnc_res_0_i_i);
    
    un4_bnc_res_16 : XOR2
      port map(A => \BNC_CNT[16]_net_1\, B => REG_420, Y => 
        un4_bnc_res_16_i_i);
    
    CRC32_120 : MUX2H
      port map(A => \CRC32[27]_net_1\, B => N_1142, S => N_1469_0, 
        Y => \CRC32_120\);
    
    un2_bnc_cnt_I_142 : AND3
      port map(A => \DWACT_FINC_E[28]\, B => \DWACT_FINC_E[13]\, 
        C => \DWACT_FINC_E[16]\, Y => N_61);
    
    EVNT_NUM_2_I_63 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_3[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_1[0]\);
    
    READ_OR_FLAG_91_i_0_x2 : XOR2
      port map(A => \STATE1[0]_net_1\, B => \STATE1[2]_net_1\, Y
         => N_258_i_0);
    
    EVNT_NUM_2_I_44 : XOR2
      port map(A => \EVNT_NUM[6]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => \EVNT_NUM_2[6]\);
    
    \BNC_CNT[21]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_237\, CLR => 
        CLEAR_3, Q => \BNC_CNT[21]_net_1\);
    
    EVENT_DWORD_148 : MUX2H
      port map(A => \EVENT_DWORD[10]_net_1\, B => 
        \EVENT_DWORD_17[10]\, S => un1_STATE1_18_1, Y => 
        \EVENT_DWORD_148\);
    
    \FID_6_r[5]\ : AND3FFT
      port map(A => N_1522, B => \FID_6_iv_0_0_0[5]_net_1\, C => 
        N_532_3_6, Y => \FID_6[5]\);
    
    un4_bnc_res_18 : XOR2
      port map(A => \BNC_CNT[18]_net_1\, B => REG_422, Y => 
        un4_bnc_res_18_i_i);
    
    un1_CNT_1_I_31 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \CNT_0[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12_0[0]\);
    
    CRC32_106 : MUX2H
      port map(A => \CRC32[13]_net_1\, B => N_1380, S => N_1469_1, 
        Y => \CRC32_106\);
    
    un2_bnc_cnt_I_27 : AND2
      port map(A => \BNC_CNT[3]_net_1\, B => \BNC_CNT[4]_net_1\, 
        Y => \DWACT_FINC_E[1]\);
    
    \un2_i2c_chain_0_0_0_1[4]\ : OAI21FTT
      port map(A => N_1691_1, B => \CNT_0[5]_net_1\, C => 
        \un2_i2c_chain_0_0_0_a2_1[4]_net_1\, Y => 
        \un2_i2c_chain_0_0_0_1_i[4]\);
    
    \BNC_CNT_3[21]\ : AND2
      port map(A => I_136, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[21]_net_1\);
    
    \ORATETMO_7_0_0_a2_1[0]\ : NOR2FT
      port map(A => \STATE1_0[2]_net_1\, B => N_221, Y => 
        N_1576_1);
    
    un1_REG_1_G_11_0_o2 : AO21TTF
      port map(A => I_8, B => \REG[42]\, C => G_11_0_a2_0, Y => 
        I10_un1_CO1);
    
    un1_ORATETMO_1_I_9 : XOR2
      port map(A => \ORATETMO_i_i[1]\, B => N_701_i_0, Y => 
        \DWACT_ADD_CI_0_pog_array_0[0]\);
    
    BNC_CNT_222 : MUX2H
      port map(A => \BNC_CNT[6]_net_1\, B => \BNC_CNT_3[6]_net_1\, 
        S => LBSP_c(2), Y => \BNC_CNT_222\);
    
    FID_191 : MUX2H
      port map(A => \FID[21]_net_1\, B => \FID_6[21]\, S => 
        N_205_0, Y => \FID_191\);
    
    \BNC_CNT_3[31]\ : AND2
      port map(A => I_224, B => un4_bnc_res_i_0, Y => 
        \BNC_CNT_3[31]_net_1\);
    
    FAULT_STAT : DFFC
      port map(CLK => CLK_c_c, D => \FAULT_STAT_126\, CLR => 
        HWRES_c_11, Q => \FAULT_STAT\);
    
    \EVENT_DWORD_17_r[8]\ : AND3FFT
      port map(A => N_1663, B => \EVENT_DWORD_17_i_0_0[8]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[8]\);
    
    \BNC_CNT_3[12]\ : AND2
      port map(A => I_73_0, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[12]_net_1\);
    
    FID_193 : MUX2H
      port map(A => \FID[23]_net_1\, B => \FID_6[23]\, S => 
        N_205_0, Y => \FID_193\);
    
    \EVNT_NUM[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[4]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[4]_net_1\);
    
    un1_ORATETMO_1_I_19 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[1]\, B => 
        \DWACT_ADD_CI_0_TMP_2[0]\, Y => I_19);
    
    \EVENT_DWORD[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_152\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[14]_net_1\);
    
    \CNT_8_i_o2[0]\ : OA21
      port map(A => N_183, B => N_192, C => N_532_3_3, Y => 
        N_185_i);
    
    \FID_6_r[12]\ : OA21
      port map(A => N_1508_i, B => \FID_6_iv_0_0_0_i[12]\, C => 
        N_532_3_5, Y => \FID_6[12]\);
    
    \FID_6_0_iv_0_0_a2[1]\ : NOR2
      port map(A => GA_c(1), B => N_235, Y => N_1503_i);
    
    un4_bnc_res_NE_18 : OR3
      port map(A => un4_bnc_res_NE_7_i, B => un4_bnc_res_5_i_i, C
         => un4_bnc_res_7_i_i, Y => un4_bnc_res_NE_18_i);
    
    \un2_i2c_chain_0_0_0_o2_1[4]\ : AND2
      port map(A => \CNT[0]_net_1\, B => N_1769, Y => N_1615_i);
    
    L2AS : DFFC
      port map(CLK => ALICLK_c, D => \L2AS_1\, CLR => HWRES_c_12, 
        Q => \REG[334]\);
    
    \CRC32_2_i_0[10]\ : NOR2FT
      port map(A => N_532_3_1, B => N_278_i_i_0, Y => N_1289);
    
    un1_REG_1_G_27_i_a2 : OR2
      port map(A => I_16, B => \FIFO_END_EVNT\, Y => 
        ADD_16x16_slow_I3_CO1_1_0_i_i);
    
    un4_bnc_res_NE_1 : OR2
      port map(A => un4_bnc_res_26_i_i, B => un4_bnc_res_29_i_i, 
        Y => un4_bnc_res_NE_1_i);
    
    \CRC32_2_i_0[20]\ : NOR2FT
      port map(A => N_532_3_2, B => N_286_i_i_0, Y => N_1383);
    
    un1_STATE1_24_i_i_a2_1 : OR3
      port map(A => N_252, B => N_242, C => \STATE1[2]_net_1\, Y
         => \un1_STATE1_24_i_i_a2_1\);
    
    \FID_6_iv_0_0_a2[18]\ : OR2FT
      port map(A => \EVNT_NUM[2]_net_1\, B => N_1575_1, Y => 
        N_1547);
    
    \EVENT_DWORD_17_i_0_1[24]\ : OAI21FTF
      port map(A => N_1454_0, B => OR_RDATA(4), C => 
        \EVENT_DWORD_17_i_0_0[24]_net_1\, Y => 
        \EVENT_DWORD_17_i_0_1[24]_net_1\);
    
    READ_PDL_FLAG_92_0_0_o2 : OR2
      port map(A => \STATE1_0[3]_net_1\, B => \STATE1_0[2]_net_1\, 
        Y => N_266);
    
    \FID_6_iv_0_0_a2_0[28]\ : NOR2FT
      port map(A => \EVENT_DWORD[28]_net_1\, B => N_620_4, Y => 
        N_1536_i);
    
    \REG_1[47]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I15_Y, CLR => 
        CLEAR_19, Q => \REG[47]\);
    
    \REG_1[32]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I0_S, CLR => 
        CLEAR_18, Q => \REG[32]\);
    
    un4_bnc_res_1 : XOR2
      port map(A => \BNC_CNT[1]_net_1\, B => REG_405, Y => 
        un4_bnc_res_1_i_i);
    
    \CNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => N_78, CLR => CLEAR_6, Q => 
        \CNT[2]_net_1\);
    
    \un2_i2c_chain_0_0_0_0[1]\ : OAI21TTF
      port map(A => N_218, B => N_1774, C => N_1630_i, Y => 
        \un2_i2c_chain_0_0_0_0_i[1]\);
    
    \STATE1_ns_0_0_0_a2_2[3]\ : OR3FTT
      port map(A => N_1771, B => \STATE1_d[7]\, C => 
        \STATE1[3]_net_1\, Y => N_1734);
    
    un2_i2c_chain_0_0_0_3_113 : OA21TTF
      port map(A => N_1770, B => 
        \un2_i2c_chain_0_0_0_a2_1_0[3]_net_1\, C => N_194, Y => 
        N_7192_i);
    
    \STATE1_ns_1_iv_0_0_3[2]\ : AOI21TTF
      port map(A => N_1587, B => 
        \STATE1_ns_1_iv_0_0_a2_4_1[2]_net_1\, C => 
        \STATE1_ns_1_iv_0_0_1[2]_net_1\, Y => 
        \STATE1_ns_1_iv_0_0_3[2]_net_1\);
    
    \EVENT_DWORD_17_i_0_a2_0[11]\ : NOR2
      port map(A => \EVENT_DWORD[11]_net_1\, B => N_1229_i_1, Y
         => N_336);
    
    \BNC_CNT[9]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_225\, CLR => 
        CLEAR_4, Q => \BNC_CNT[9]_net_1\);
    
    un1_STATE1_17_i_0_i4_1_a2_0_i2_0_a2 : OR2FT
      port map(A => \STATE1[0]_net_1\, B => \STATE1_0[3]_net_1\, 
        Y => N_120_i);
    
    \EVNT_NUM[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[3]\, CLR => 
        CLEAR_12, Q => \EVNT_NUM[3]_net_1\);
    
    un4_bnc_res_26 : XOR2
      port map(A => \BNC_CNT[26]_net_1\, B => REG_430, Y => 
        un4_bnc_res_26_i_i);
    
    un4_bnc_res_28 : XOR2
      port map(A => \BNC_CNT[28]_net_1\, B => REG_432, Y => 
        un4_bnc_res_28_i_i);
    
    \OR_RADDR[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \OR_RADDR_206\, CLR => 
        CLEAR_16, Q => \OR_RADDR[2]_net_1\);
    
    un1_ORATETMO_1_I_17_i : NOR2FT
      port map(A => N_193, B => N_252, Y => N_701_i_0);
    
    un2_bnc_cnt_I_196 : XOR2
      port map(A => N_24, B => \BNC_CNT[27]_net_1\, Y => I_196);
    
    un2_bnc_cnt_I_176 : AND2
      port map(A => \BNC_CNT[24]_net_1\, B => \BNC_CNT[25]_net_1\, 
        Y => \DWACT_FINC_E[20]\);
    
    \CRC32_2_i_0[30]\ : NOR2FT
      port map(A => N_532_3_2, B => N_260_i_i_0, Y => N_1294);
    
    \CRC32[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_95\, CLR => CLEAR_8, Q
         => \CRC32[2]_net_1\);
    
    \un2_i2c_chain_0_0_0_a2_0_1[4]\ : OR2FT
      port map(A => \CNT_0[1]_net_1\, B => N_1765, Y => 
        \un2_i2c_chain_0_0_0_a2_0_i[4]\);
    
    \FID_6_iv_0_0_0[15]\ : OAI21
      port map(A => N_1575_0, B => N_57_i_0_i, C => N_1477, Y => 
        \FID_6_iv_0_0_0_i[15]\);
    
    \FID[23]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_193\, CLR => CLEAR_14, Q
         => \FID[23]_net_1\);
    
    un2_bnc_cnt_I_19 : AND2
      port map(A => \BNC_CNT[3]_net_1\, B => \DWACT_FINC_E[0]\, Y
         => N_149);
    
    un1_REG_1_ADD_16x16_slow_I14_un1_CO1_m7_4 : NAND3
      port map(A => ADD_16x16_slow_I14_un1_CO1_m7_1, B => 
        \REG[39]\, C => \REG[41]\, Y => 
        ADD_16x16_slow_I14_un1_CO1_m7_4_i);
    
    un1_ORATETMO_1_I_15 : XOR2
      port map(A => \ORATETMO[2]_net_1\, B => N_701_i_0_0, Y => 
        \DWACT_ADD_CI_0_partial_sum[2]\);
    
    \FID_6_iv_0_0_0[28]\ : OAI21FTT
      port map(A => REG_71, B => N_1574, C => N_1575, Y => 
        \FID_6_iv_0_0_0_i[28]\);
    
    FID_174 : MUX2H
      port map(A => \FID[4]_net_1\, B => \FID_6[4]\, S => N_205, 
        Y => \FID_174\);
    
    \un2_i2c_chain_0_0_0_3[1]\ : AO21TTF
      port map(A => \CNT[1]_net_1\, B => N_1638_1, C => 
        \un2_i2c_chain_0_0_0_1[1]_net_1\, Y => 
        \un2_i2c_chain_0_0_0_3_i[1]\);
    
    READ_PDL_FLAG_92_0_0_0 : AO21TTF
      port map(A => \READ_PDL_FLAG\, B => \STATE1[0]_net_1\, C
         => N_1669_i, Y => \READ_PDL_FLAG_92_0_0_0\);
    
    L2RS : DFFC
      port map(CLK => ALICLK_c, D => \L2RS_1\, CLR => HWRES_c_12, 
        Q => REG_330);
    
    \CNT_8_i[0]\ : AND2
      port map(A => N_185_i, B => \DWACT_ADD_CI_0_partial_sum[0]\, 
        Y => \CNT_8_i[0]_net_1\);
    
    CRC32_100 : MUX2H
      port map(A => \CRC32[7]_net_1\, B => N_1596, S => N_1469, Y
         => \CRC32_100\);
    
    un4_bnc_res_NE_29 : OR3
      port map(A => un4_bnc_res_NE_27_i, B => un4_bnc_res_NE_21_i, 
        C => un4_bnc_res_NE_22_i, Y => un4_bnc_res_NE_29_i);
    
    un2_bnc_cnt_I_8 : AND2
      port map(A => \BNC_CNT[1]_net_1\, B => \BNC_CNT[0]_net_1\, 
        Y => N_157);
    
    un1_REG_1_ADD_16x16_slow_I10_S_0 : XOR2FT
      port map(A => \REG[42]\, B => \un2_evread_1[14]\, Y => 
        ADD_16x16_slow_I10_S_0);
    
    \STATE1_ns_0_0_0_a2[3]\ : OR3FFT
      port map(A => \STATE1_0[3]_net_1\, B => N_230, C => 
        \STATE1_0[2]_net_1\, Y => N_1731);
    
    \BNC_CNT[16]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_232\, CLR => 
        CLEAR_2, Q => \BNC_CNT[16]_net_1\);
    
    \STATE2[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE2_ns[2]\, CLR => 
        CLEAR_19, Q => \STATE2[0]_net_1\);
    
    \EVENT_DWORD_17_r[28]\ : AND3FFT
      port map(A => N_1694, B => \EVENT_DWORD_17_i_0_1[28]_net_1\, 
        C => N_532_3_6, Y => \EVENT_DWORD_17[28]\);
    
    \CRC32[28]\ : DFFC
      port map(CLK => CLK_c_c, D => \CRC32_121\, CLR => CLEAR_8, 
        Q => \CRC32[28]_net_1\);
    
    \BNC_CNT_3[10]\ : AND2
      port map(A => I_56_0, B => un4_bnc_res_i, Y => 
        \BNC_CNT_3[10]_net_1\);
    
    \FID_6_iv_0_0_0[4]\ : OAI21
      port map(A => N_1575_0, B => \FID_2_i[4]\, C => N_342, Y
         => \FID_6_iv_0_0_0_i[4]\);
    
    \FID[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_184\, CLR => CLEAR_13, Q
         => \FID[14]_net_1\);
    
    \EVENT_DWORD_17_i_1[27]\ : OAI21FTF
      port map(A => N_1454, B => OR_RDATA(7), C => 
        \EVENT_DWORD_17_i_0[27]_net_1\, Y => 
        \EVENT_DWORD_17_i_1[27]_net_1\);
    
    un4_bnc_res_2 : XOR2
      port map(A => \BNC_CNT[2]_net_1\, B => REG_406, Y => 
        un4_bnc_res_2_i_i);
    
    un1_STATE1_24_i_i_o2_0 : NOR2FT
      port map(A => \OR_RACK_sync\, B => N_226_i_0, Y => N_242);
    
    \EVENT_DWORD_17_i_0[27]\ : OAI21TTF
      port map(A => N_105_i_0_0, B => PDL_RDATA(3), C => N_1678, 
        Y => \EVENT_DWORD_17_i_0[27]_net_1\);
    
    un4_bnc_res_NE_7 : OR2
      port map(A => un4_bnc_res_10_i_i, B => un4_bnc_res_13_i_i, 
        Y => un4_bnc_res_NE_7_i);
    
    FID_180 : MUX2H
      port map(A => \FID[10]_net_1\, B => \FID_6[10]\, S => 
        N_205_1, Y => \FID_180\);
    
    \FID[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_170\, CLR => CLEAR_13, Q
         => \FID[0]_net_1\);
    
    FAULT_STROBE_2 : NOR2
      port map(A => \CLEAR_PSM_FLAGS\, B => FAULT_STROBE_0_i, Y
         => \FAULT_STROBE_2\);
    
    \REG_1[36]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I4_S, CLR => 
        CLEAR_18, Q => \REG[36]\);
    
    \EVENT_DWORD_17_i_0_o2_0[3]\ : NOR2FT
      port map(A => N_1768_i, B => N_1454_0, Y => N_190_i_0);
    
    \EVENT_DWORD_17_i_0_0[7]\ : OAI21TTF
      port map(A => \EVENT_DWORD[15]_net_1\, B => N_105_i_0, C
         => N_1620, Y => \EVENT_DWORD_17_i_0_0[7]_net_1\);
    
    un2_bnc_cnt_I_76 : AND3
      port map(A => \DWACT_FINC_E[6]\, B => \DWACT_FINC_E[7]\, C
         => \BNC_CNT[12]_net_1\, Y => N_108);
    
    un2_bnc_cnt_I_217 : XOR2
      port map(A => N_9, B => \BNC_CNT[30]_net_1\, Y => I_217);
    
    un1_REG_1_G_18_0_o2 : AO21TTF
      port map(A => I8_un1_CO1, B => \REG[41]\, C => 
        ADD_16x16_slow_I9_CO1_0, Y => N224);
    
    I2C_CHAIN_128 : MUX2H
      port map(A => I2C_CHAIN_net_1, B => N_93, S => 
        I2C_RREQ_1_sqmuxa, Y => \I2C_CHAIN_128\);
    
    CHIP_ADDR_135 : MUX2H
      port map(A => \CHIP_ADDR[2]_net_1\, B => N_96, S => 
        I2C_RREQ_1_sqmuxa, Y => \CHIP_ADDR_135\);
    
    \OR_RADDR_3_i_0_0[3]\ : AND2
      port map(A => N_532_3_3, B => \CNT_0[3]_net_1\, Y => N_683);
    
    un2_bnc_cnt_I_72 : AND2
      port map(A => \DWACT_FINC_E[7]\, B => \DWACT_FINC_E[6]\, Y
         => N_111);
    
    \ORATETMO_7_0_0[1]\ : OR2
      port map(A => N_233, B => I_19, Y => \ORATETMO_7[1]\);
    
    un2_bnc_cnt_I_84 : XOR2
      port map(A => N_103, B => \BNC_CNT[14]_net_1\, Y => I_84_0);
    
    un5_evread_11 : OR3
      port map(A => un5_evread_7, B => \un5_evread_1\, C => 
        un5_evread_6_i, Y => un5_evread_11_i);
    
    \EVENT_DWORD[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_145\, CLR => 
        CLEAR_11, Q => \EVENT_DWORD[7]_net_1\);
    
    \CRC32_2_i_0_x2[22]\ : XOR2FT
      port map(A => \CRC32[22]_net_1\, B => 
        \EVENT_DWORD[22]_net_1\, Y => N_1782_i_0);
    
    un1_STATE1_1_0_a5_0_a2 : NOR2FT
      port map(A => N_1585, B => \STATE1_0[2]_net_1\, Y => N_795);
    
    \STATE1_ns_1_iv_0_1_o2_3_o3_0_0[0]\ : AO21
      port map(A => N_1593, B => \STATE1[1]_net_1\, C => 
        \STATE1[3]_net_1\, Y => 
        \STATE1_ns_1_iv_0_1_o2_3_o3_0[0]_net_1\);
    
    \un2_i2c_chain_0_0_0_0_o2[5]\ : OR2
      port map(A => \CNT_0[2]_net_1\, B => \CNT_0[3]_net_1\, Y
         => N_188);
    
    un1_STATE1_18_0_0 : NAND3FTT
      port map(A => N_1673_i, B => N_1672, C => N_1762, Y => 
        un1_STATE1_18);
    
    \FID_6_iv_0_a2_1[19]\ : NOR2FT
      port map(A => \EVENT_DWORD[19]_net_1\, B => N_620_4_1, Y
         => N_324_i);
    
    \FID[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \FID_175\, CLR => CLEAR_15, Q
         => \FID[5]_net_1\);
    
    \EVENT_DWORD_17_i_0_0[23]\ : OAI21TTF
      port map(A => \EVENT_DWORD[31]_net_1\, B => N_105_i_0_0, C
         => N_1715, Y => \EVENT_DWORD_17_i_0_0[23]_net_1\);
    
    \STATE1_0[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \STATE1_ns[2]\, CLR => 
        CLEAR_0, Q => \STATE1_0[2]_net_1\);
    
    \CRC32_2_i_x2[29]\ : XOR2FT
      port map(A => \CRC32[29]_net_1\, B => 
        \EVENT_DWORD[29]_net_1\, Y => N_248_i_i_0);
    
    un1_I2C_RREQ_1_sqmuxa_0_0_0_o2 : OR2
      port map(A => N_1592, B => N_1593, Y => N_293);
    
    \BNC_CNT_3[17]\ : AND2
      port map(A => I_105, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[17]_net_1\);
    
    un1_ORATETMO_1_I_22 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, Y => I_22);
    
    BNC_CNT_234 : MUX2H
      port map(A => \BNC_CNT[18]_net_1\, B => 
        \BNC_CNT_3[18]_net_1\, S => LBSP_c_1(2), Y => 
        \BNC_CNT_234\);
    
    \FID_6_0_iv_0_a2_1[30]\ : NOR2
      port map(A => \EVENT_DWORD[30]_net_1\, B => N_620_4, Y => 
        N_1516);
    
    \EVENT_DWORD_17_i_a2[19]\ : NOR2
      port map(A => \EVENT_DWORD[29]_net_1\, B => N_190_i_0, Y
         => N_1675);
    
    \EVENT_DWORD_17_i_0_a2[11]\ : NOR2
      port map(A => \EVENT_DWORD[21]_net_1\, B => N_190_i_0, Y
         => N_335);
    
    \EVENT_DWORD[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_148\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[10]_net_1\);
    
    un1_ORATETMO_1_I_1 : AND2
      port map(A => \ORATETMO_i_i[0]\, B => N_701_i_0_0, Y => 
        \DWACT_ADD_CI_0_TMP_2[0]\);
    
    \CRC32_2_i_0_x2[0]\ : XOR2FT
      port map(A => \CRC32[0]_net_1\, B => \EVENT_DWORD[0]_net_1\, 
        Y => N_254_i_i_0);
    
    EVRDYi : DFFC
      port map(CLK => CLK_c_c, D => \EVRDYi_202\, CLR => CLEAR_12, 
        Q => \EVRDY_c\);
    
    \un2_i2c_chain_0_0_0_a2[3]\ : OR3FFT
      port map(A => \CNT_0[2]_net_1\, B => N_1603, C => N_186, Y
         => N_1633);
    
    un2_bnc_cnt_I_139 : AND2
      port map(A => \DWACT_FINC_E[15]\, B => \BNC_CNT[21]_net_1\, 
        Y => \DWACT_FINC_E[16]\);
    
    un1_evread_0 : OR2FT
      port map(A => EVREAD, B => \FIFO_END_EVNT\, Y => 
        \un2_evread_0[14]\);
    
    \FID_6_0_iv_0_0_o2[3]\ : NOR2FT
      port map(A => N_1575_0, B => N_1587, Y => N_235);
    
    un1_REG_1_G_18 : AND2
      port map(A => \FIFO_END_EVNT\, B => 
        ADD_16x16_slow_I6_un4_CO1_5_tz, Y => N_19);
    
    \FID_6_r[1]\ : OA21
      port map(A => N_1503_i, B => \FID_6_0_iv_0_0_0_i[1]\, C => 
        N_532_3_6, Y => \FID_6[1]\);
    
    \FID_6_iv_0_0_1[18]\ : OAI21FTT
      port map(A => REG_61, B => N_1574_1, C => 
        \FID_6_iv_0_0_0[18]_net_1\, Y => \FID_6_iv_0_0_1_i[18]\);
    
    \BNC_CNT_3[11]\ : AND2
      port map(A => I_66_0, B => un4_bnc_res_i_1, Y => 
        \BNC_CNT_3[11]_net_1\);
    
    \BNC_CNT[8]\ : DFFC
      port map(CLK => ALICLK_c, D => \BNC_CNT_224\, CLR => 
        CLEAR_4, Q => \BNC_CNT[8]_net_1\);
    
    \REG_1[38]\ : DFFC
      port map(CLK => CLK_c_c, D => ADD_16x16_slow_I6_S, CLR => 
        CLEAR_18, Q => \REG[38]\);
    
    \un2_i2c_chain_0_0_0_o2_0[4]\ : OR2FT
      port map(A => \CNT_0[1]_net_1\, B => \CNT_0[0]_net_1\, Y
         => N_216);
    
    un2_bnc_cnt_I_37 : AND3
      port map(A => \DWACT_FINC_E[0]\, B => \DWACT_FINC_E[2]\, C
         => \BNC_CNT[6]_net_1\, Y => N_136);
    
    un1_CNT_1_I_23 : XOR2
      port map(A => \CNT[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, Y => I_23);
    
    \FID_6_iv_0_0_a2[9]\ : NOR2
      port map(A => \FID_2[9]_net_1\, B => N_1575, Y => N_1526);
    
    un2_bnc_cnt_I_41 : AND2
      port map(A => \BNC_CNT[6]_net_1\, B => \BNC_CNT[7]_net_1\, 
        Y => \DWACT_FINC_E[3]\);
    
    I2C_RREQ_137 : MUX2H
      port map(A => I2C_RREQ_net_1, B => \STATE1_d_i[7]_net_1\, S
         => un1_I2C_RREQ_1_sqmuxa, Y => \I2C_RREQ_137\);
    
    \EVENT_DWORD_17_r[0]\ : AND3FFT
      port map(A => N_1641, B => \EVENT_DWORD_17_i_0_0[0]_net_1\, 
        C => N_532_3_8, Y => \EVENT_DWORD_17[0]\);
    
    un1_REG_1_ADD_16x16_slow_I12_S : XOR2
      port map(A => N228, B => ADD_16x16_slow_I12_S_0, Y => 
        ADD_16x16_slow_I12_S);
    
    \EVENT_DWORD[21]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_159\, CLR => 
        CLEAR_10, Q => \EVENT_DWORD[21]_net_1\);
    
    \ORATETMO_7_0_0_a2_0[0]\ : AND2FT
      port map(A => \READ_ADC_FLAG\, B => \READ_OR_FLAG\, Y => 
        \ORATETMO_7_0_0_a2_0[0]_net_1\);
    
    \EVENT_DWORD[16]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVENT_DWORD_154\, CLR => 
        CLEAR_9, Q => \EVENT_DWORD[16]_net_1\);
    
    \un2_i2c_chain_0_0_0_a2_4[3]\ : OR3FTT
      port map(A => \CNT_0[4]_net_1\, B => N_1769, C => N_216, Y
         => \un2_i2c_chain_0_0_0_a2_4[3]_net_1\);
    
    L2RF2 : DFFC
      port map(CLK => ALICLK_c, D => \L2RF1\, CLR => HWRES_c_12, 
        Q => \L2RF2\);
    
    \un2_i2c_chain_0_0_0[3]\ : OR3
      port map(A => N_7192_i, B => \un2_i2c_chain_0_0_0_2_i[3]\, 
        C => \un2_i2c_chain_0_0_0_1_i[3]\, Y => N_96);
    
    \EVNT_NUM[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \EVNT_NUM_2[10]\, CLR => 
        CLEAR_11, Q => \EVNT_NUM[10]_net_1\);
    
    \ORATETMO_7_0_0[4]\ : OR2
      port map(A => N_233, B => I_22, Y => \ORATETMO_7[4]\);
    
    \EVENT_DWORD_17_r[13]\ : AND3FFT
      port map(A => N_339, B => \EVENT_DWORD_17_i_0_0[13]_net_1\, 
        C => N_532_3_7, Y => \EVENT_DWORD_17[13]\);
    
    EVNT_NUM_2_I_59 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_11_1[0]\, B => 
        \EVNT_NUM[10]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12_4[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity I2C_INTERF is

    port( PULSE         : in    std_logic_vector(7 to 7);
          I2C_RDATA     : out   std_logic_vector(9 downto 0);
          CHIP_ADDR     : in    std_logic_vector(2 downto 0);
          CHANNEL       : in    std_logic_vector(2 downto 0);
          TICK          : in    std_logic_vector(0 to 0);
          TICK_2        : in    std_logic_vector(0 to 0);
          REG_107       : out   std_logic;
          REG_108       : out   std_logic;
          REG_109       : out   std_logic;
          REG_110       : out   std_logic;
          REG_111       : out   std_logic;
          REG_112       : out   std_logic;
          REG_113       : out   std_logic;
          REG_114       : out   std_logic;
          REG_0         : in    std_logic;
          REG_84        : in    std_logic;
          REG_85        : in    std_logic;
          REG_91        : in    std_logic;
          REG_92        : in    std_logic;
          REG_99        : out   std_logic;
          REG_93        : in    std_logic;
          REG_94        : in    std_logic;
          REG_95        : in    std_logic;
          REG_96        : in    std_logic;
          REG_97        : in    std_logic;
          REG_98        : in    std_logic;
          REG_83        : in    std_logic;
          REG_100       : out   std_logic;
          TICK_1        : in    std_logic_vector(0 to 0);
          TICK_0        : in    std_logic_vector(0 to 0);
          HWRES_c_4     : in    std_logic;
          HWRES_c_7     : in    std_logic;
          HWRES_c_11    : in    std_logic;
          HWRES_c_10    : in    std_logic;
          HWRES_c_5     : in    std_logic;
          HWRES_c_3     : in    std_logic;
          HWRES_c_6     : in    std_logic;
          I2C_RACK      : out   std_logic;
          SDAout_del2   : out   std_logic;
          HWRES_c_9     : in    std_logic;
          HWRES_c_8     : in    std_logic;
          un1_sdaa_0_a3 : out   std_logic;
          RUN_c_0_0     : in    std_logic;
          RUN_c_0       : in    std_logic;
          I2C_CHAIN     : in    std_logic;
          I2C_RREQ      : in    std_logic;
          SDA1_in       : in    std_logic;
          SDA0_in       : in    std_logic;
          un1_sdab_i    : out   std_logic;
          SCLB_i_a3     : out   std_logic;
          SCLA_i_a3     : out   std_logic;
          HWRES_c_10_0  : in    std_logic;
          CLK_c_c       : in    std_logic;
          HWRES_c_7_0   : in    std_logic
        );

end I2C_INTERF;

architecture DEF_ARCH of I2C_INTERF is 

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OA21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component NAND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \REG_0[105]\, \REG_1_105_13\, \sstate2_0[9]_net_1\, 
        \sstate2_ns_e[0]\, \sstate_0[13]_net_1\, \sstate_ns_e[0]\, 
        N_279_0, N_594_0, \sstate2[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \BITCNT[1]_net_1\, \I2C_RACK_2_i\, I2C_RACK_2, 
        \CHAIN_SELECT\, \SCL\, \sstatese_3_i_m2_i\, 
        \sstate[9]_net_1\, N_610, \sstate[10]_net_1\, 
        \sstate2se_6_i_i\, \sstate2[3]_net_1\, N_603, N_279, 
        \sstate2_i_0_i[2]\, \SDAnoe_del2\, \sstate2se_4_i_i\, 
        \sstate2[5]_net_1\, N_571, \sstate2[4]_net_1\, 
        \sstate2se_5_i_i\, N_569, \sstate2se_7_i_i\, N_567, 
        \sstate2se_8_i_i\, N_565, \sstate2[0]_net_1\, 
        \DATA_12_iv[1]\, \DATA_12_iv_0_a3_0_0_i[1]\, N_597, 
        \sstate[1]_net_1\, N_587, \un1_scl5_6_0_a2\, N_400, N_395, 
        \sstate_ns_e[2]\, \sstate[11]_net_1\, \sstate[12]_net_1\, 
        \sstate_ns_e[6]\, \sstate[7]_net_1\, \sstate[8]_net_1\, 
        \sstate_ns_e[7]\, \sstate[6]_net_1\, \sstate_ns_e[9]\, 
        \sstate[4]_net_1\, \sstate[5]_net_1\, \sstate_ns_e[10]\, 
        \sstate[3]_net_1\, \sstate_ns_e[12]\, \sstate[2]_net_1\, 
        \sstate_ns_e[13]\, \sstate[0]_net_1\, \sstate_ns_e[11]\, 
        BITCNT_2_sqmuxa, \sstate_ns_e[8]\, N_457, 
        \sstatese_7_0_0\, N_432, N_397, \sstate_ns_e[5]\, N_399, 
        \sstatese_4_0_0\, N_436, \sstate_ns_e[3]\, 
        \COMMAND[2]_net_1\, N_609_1, N_608, \sstate_ns_e[1]\, 
        N_441, N_398, N_600, \sstatese_13_0\, N_442, \PULSE_FL\, 
        \sstate2se_2_i_0\, \sstate2[6]_net_1\, N_108, 
        \sstate2[7]_net_1\, \sstate2se_3_i_0\, N_573, 
        \sstate2_ns_e[2]\, \sstate2[8]_net_1\, N_109, 
        \sstate2_ns_e[1]\, N_133_1, N_111, N_113_i, N_544, 
        \SDAnoe_48\, \SDAnoe\, SDAnoe_8, \SDAnoe_m_3\, N_403, 
        \SDAnoe_m_i\, \SDAnoe_m_1\, N_454, N_581, 
        \AIR_COMMAND_47\, \AIR_COMMAND_19[15]\, 
        \AIR_COMMAND[15]_net_1\, un1_scl5_7, N_128, 
        \AIR_COMMAND_46\, \AIR_COMMAND_19[14]\, 
        \AIR_COMMAND[14]_net_1\, N_545_i_i, N_126_i, N_127_i, 
        \AIR_COMMAND_45\, \AIR_COMMAND_19[13]\, 
        \AIR_COMMAND[13]_net_1\, N_124, \AIR_COMMAND_44\, 
        \AIR_COMMAND_19[12]\, \AIR_COMMAND[12]_net_1\, 
        \sstate2[9]_net_1\, \AIR_COMMAND_43\, 
        \AIR_COMMAND_19[11]\, \AIR_COMMAND[11]_net_1\, N_121, 
        \AIR_COMMAND_42\, \AIR_COMMAND_19[10]\, 
        \AIR_COMMAND[10]_net_1\, 
        \AIR_COMMAND_19_0_iv_0_0[10]_net_1\, N_118_i, 
        \AIR_COMMAND_19_0_iv_0_a2_1_i[10]\, 
        \AIR_COMMAND_19_0_iv_0_a2_0_i[10]\, N_578, 
        \AIR_COMMAND_19_0_iv_0_o2_0[10]_net_1\, \AIR_COMMAND_41\, 
        \AIR_COMMAND_19[9]\, \AIR_COMMAND[9]_net_1\, N_116, N_543, 
        N_548, \AIR_COMMAND_40\, \AIR_COMMAND_19[8]\, 
        \AIR_COMMAND[8]_net_1\, N_145, 
        \AIR_COMMAND_19_0_iv_0_a2_1[8]_net_1\, 
        \AIR_COMMAND_19_0_iv_0_0_i[8]\, \REG[105]\, 
        \AIR_COMMAND_39\, N_542, \AIR_COMMAND[2]_net_1\, N_144, 
        \AIR_COMMAND_19_i_0[2]_net_1\, N_143, N_564_1, 
        \AIR_COMMAND_38\, N_541, \AIR_COMMAND[1]_net_1\, 
        \AIR_COMMAND_19_i_0_i[1]\, N_577, \AIR_COMMAND_37\, N_540, 
        \AIR_COMMAND[0]_net_1\, N_563, N_564_i, 
        un1_scl5_7_0_a2_0_2_i, un1_scl5_7_0_a2_0_0, N_137, 
        \SDAout_36\, \SDAout\, SDAout_12, N_506, 
        \un1_sstate_12_0_0_0\, N_402, \COMMAND[0]_net_1\, 
        SDAout_m_i_i, \COMMAND_m_i[15]\, \SBYTE_m_i[7]\, 
        \SBYTE[7]_net_1\, N_512, \COMMAND[15]_net_1\, 
        \COMMAND[1]_net_1\, SDAout_m_1_i, \SBYTE_35\, 
        \SBYTE_9[7]_net_1\, N_449, \SBYTE[6]_net_1\, \SBYTE_34\, 
        \SBYTE_9[6]_net_1\, \SBYTE[5]_net_1\, \COMMAND[14]_net_1\, 
        \SBYTE_33\, \SBYTE_9[5]_net_1\, \SBYTE[4]_net_1\, 
        \COMMAND[13]_net_1\, \SBYTE_32\, \SBYTE_9[4]_net_1\, 
        \SBYTE[3]_net_1\, \COMMAND[12]_net_1\, \SBYTE_31\, 
        \SBYTE_9[3]_net_1\, \SBYTE[2]_net_1\, \COMMAND[11]_net_1\, 
        \SBYTE_30\, \SBYTE_9[2]_net_1\, \SBYTE[1]_net_1\, 
        \COMMAND[10]_net_1\, \SBYTE_29\, \SBYTE_9[1]_net_1\, 
        \SBYTE[0]_net_1\, \COMMAND[9]_net_1\, \SBYTE_28\, 
        \SBYTE_9[0]\, N_596, N_615, N_626, \COMMAND[8]_net_1\, 
        \un1_sstate_10_0_o2_0_a3_0\, \SCL_27\, N_612, N_598, 
        SCL_1_iv_i_a3_0, \SCL_1_iv_i_a3_0_1\, \START_I2C_26\, 
        \START_I2C\, N_539, \START_I2C_2_iv_i_a2_0_0\, N_135, 
        \AIR_CHAIN_25\, \AIR_CHAIN\, N_538, \AIR_CHAIN_4_iv_i_0\, 
        N_133, \CHAIN_SELECT_24\, N_537, N_130, N_551, 
        \I2C_RDATA_23\, N_586, N_278, N_594, N_623, 
        \I2C_RDATA[9]_net_1\, \I2C_RDATA_22\, N_585, N_621, 
        \I2C_RDATA[8]_net_1\, \I2C_RDATA_21\, N_593, N_638, 
        \I2C_RDATA[7]_net_1\, \I2C_RDATA_20\, N_592, N_636, 
        \I2C_RDATA[6]_net_1\, \I2C_RDATA_19\, N_591, N_634, 
        \I2C_RDATA[5]_net_1\, \I2C_RDATA_18\, N_590, N_632, 
        \I2C_RDATA[4]_net_1\, \I2C_RDATA_17\, N_589, N_630, 
        \I2C_RDATA[3]_net_1\, \I2C_RDATA_16\, N_588, N_628, 
        \I2C_RDATA[2]_net_1\, \I2C_RDATA_15\, N_584, N_595, 
        \REG[120]\, N_619, \I2C_RDATA[1]_net_1\, \I2C_RDATA_14\, 
        N_583, \REG[119]\, N_617, \I2C_RDATA[0]_net_1\, 
        sstate_3_sqmuxa, N_550, \PULSE_FL_12\, \COMMAND_11\, 
        N_562, \COMMAND_10\, N_561, \COMMAND_9\, N_560, 
        \COMMAND_8\, N_559, \sstate[13]_net_1\, \COMMAND_7\, 
        N_558, \COMMAND_6\, N_557, \COMMAND_5\, N_556, 
        \COMMAND_4\, N_555, \COMMAND_3\, N_554, \COMMAND_2\, 
        N_553, \COMMAND_1\, N_552, \BITCNT_8[2]\, I_14, 
        BITCNT_0_sqmuxa_2, \BITCNT_8[1]\, I_13, \BITCNT_8[0]\, 
        \DWACT_ADD_CI_0_partial_sum[0]\, \BITCNT[2]_net_1\, 
        N_517_2, \DATA_12[15]_net_1\, DATA_1_sqmuxa_2_i, 
        \DATA_12[14]_net_1\, \DATA_12[13]_net_1\, \REG[118]\, 
        \DATA_12[12]_net_1\, \REG[117]\, \DATA_12[11]_net_1\, 
        \REG[116]\, \DATA_12[10]_net_1\, \REG[115]\, 
        \DATA_12[9]_net_1\, \REG[114]\, \DATA_12[8]_net_1\, 
        \REG[113]\, \BITCNT[0]_net_1\, \SDAnoe_del\, 
        \SDAnoe_del1\, \SDAout_del\, \SDAout_del1\, \REG[106]\, 
        \GND\, \VCC\ : std_logic;

begin 

    I2C_RDATA(9) <= \I2C_RDATA[9]_net_1\;
    I2C_RDATA(8) <= \I2C_RDATA[8]_net_1\;
    I2C_RDATA(7) <= \I2C_RDATA[7]_net_1\;
    I2C_RDATA(6) <= \I2C_RDATA[6]_net_1\;
    I2C_RDATA(5) <= \I2C_RDATA[5]_net_1\;
    I2C_RDATA(4) <= \I2C_RDATA[4]_net_1\;
    I2C_RDATA(3) <= \I2C_RDATA[3]_net_1\;
    I2C_RDATA(2) <= \I2C_RDATA[2]_net_1\;
    I2C_RDATA(1) <= \I2C_RDATA[1]_net_1\;
    I2C_RDATA(0) <= \I2C_RDATA[0]_net_1\;
    REG_107 <= \REG[113]\;
    REG_108 <= \REG[114]\;
    REG_109 <= \REG[115]\;
    REG_110 <= \REG[116]\;
    REG_111 <= \REG[117]\;
    REG_112 <= \REG[118]\;
    REG_113 <= \REG[119]\;
    REG_114 <= \REG[120]\;
    REG_99 <= \REG[105]\;
    REG_100 <= \REG[106]\;

    sstatese_0_0_a2_0 : OR3FTT
      port map(A => TICK_0(0), B => N_398, C => N_600, Y => N_441);
    
    \SBYTE[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_32\, CLR => HWRES_c_8, 
        Q => \SBYTE[4]_net_1\);
    
    \COMMAND_4_i_m2[11]\ : MUX2H
      port map(A => REG_94, B => \AIR_COMMAND[11]_net_1\, S => 
        RUN_c_0, Y => N_558);
    
    START_I2C : DFFC
      port map(CLK => CLK_c_c, D => \START_I2C_26\, CLR => 
        HWRES_c_9, Q => \START_I2C\);
    
    \SBYTE_9[4]\ : MUX2H
      port map(A => \SBYTE[3]_net_1\, B => \COMMAND[12]_net_1\, S
         => N_399, Y => \SBYTE_9[4]_net_1\);
    
    \DATA_12[15]\ : MUX2H
      port map(A => \SBYTE[7]_net_1\, B => \REG[120]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[15]_net_1\);
    
    \BITCNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_8[0]\, CLR => 
        HWRES_c_4, Q => \BITCNT[0]_net_1\);
    
    \AIR_COMMAND_19_0_iv_0[14]\ : OR3
      port map(A => N_545_i_i, B => N_126_i, C => N_127_i, Y => 
        \AIR_COMMAND_19[14]\);
    
    \AIR_COMMAND_19_0_iv_0_o2_0[12]\ : OR2
      port map(A => \sstate2[3]_net_1\, B => \sstate2[8]_net_1\, 
        Y => N_543);
    
    \I2C_RDATA_9_i_a3[8]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[8]_net_1\, Y => 
        N_621);
    
    SDAnoe : DFFS
      port map(CLK => CLK_c_c, D => \SDAnoe_48\, SET => HWRES_c_8, 
        Q => \SDAnoe\);
    
    \COMMAND_4_i_m2[12]\ : MUX2H
      port map(A => REG_95, B => \AIR_COMMAND[12]_net_1\, S => 
        RUN_c_0, Y => N_559);
    
    un1_scl5_7_0_a2_1 : OR2
      port map(A => N_543, B => \sstate2[5]_net_1\, Y => N_577);
    
    sstatese_13_a2 : AO21TTF
      port map(A => TICK_1(0), B => \PULSE_FL\, C => 
        \sstate_0[13]_net_1\, Y => N_442);
    
    SDAnoe_del1 : DFFC
      port map(CLK => CLK_c_c, D => \SDAnoe_del\, CLR => 
        HWRES_c_8, Q => \SDAnoe_del1\);
    
    SDAnoe_del : DFFC
      port map(CLK => CLK_c_c, D => \SDAnoe\, CLR => HWRES_c_8, Q
         => \SDAnoe_del\);
    
    \AIR_COMMAND[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_46\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[14]_net_1\);
    
    un1_scl5_7_0_a2_0_1 : OR2
      port map(A => \sstate2[4]_net_1\, B => \sstate2[6]_net_1\, 
        Y => N_564_1);
    
    \sstate2[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2se_4_i_i\, CLR => 
        HWRES_c_9, Q => \sstate2[4]_net_1\);
    
    AIR_CHAIN_4_iv_i_0 : OAI21TTF
      port map(A => \AIR_CHAIN\, B => \sstate2[9]_net_1\, C => 
        N_133, Y => \AIR_CHAIN_4_iv_i_0\);
    
    un1_sstate_12_0_0_0 : AO21
      port map(A => \COMMAND[2]_net_1\, B => N_454, C => 
        \sstate[9]_net_1\, Y => \un1_sstate_12_0_0_0\);
    
    un1_scl5_7_0_o2 : OR2FT
      port map(A => \sstate2_0[9]_net_1\, B => I2C_RREQ, Y => 
        N_544);
    
    \I2C_RDATA_9_i_a3[0]\ : NOR2FT
      port map(A => N_595, B => \I2C_RDATA[0]_net_1\, Y => N_617);
    
    \I2C_RDATA_9_i[6]\ : OA21TTF
      port map(A => N_594, B => \REG[117]\, C => N_636, Y => 
        N_592);
    
    sstate2se_0_0_0 : AO21FTF
      port map(A => N_133_1, B => TICK_2(0), C => N_111, Y => 
        \sstate2_ns_e[1]\);
    
    \AIR_COMMAND_19_0_iv_0_a2_1_0[8]\ : NOR3FFT
      port map(A => \sstate2[7]_net_1\, B => N_548, C => 
        \sstate2[6]_net_1\, Y => 
        \AIR_COMMAND_19_0_iv_0_a2_1[8]_net_1\);
    
    \AIR_COMMAND_19_i[2]\ : OA21TTF
      port map(A => N_144, B => \REG[105]\, C => 
        \AIR_COMMAND_19_i_0[2]_net_1\, Y => N_542);
    
    \DATA_12[12]\ : MUX2H
      port map(A => \SBYTE[4]_net_1\, B => \REG[117]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[12]_net_1\);
    
    \AIR_COMMAND[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_47\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[15]_net_1\);
    
    sstatese_5_0_m2 : MUX2H
      port map(A => \sstate[7]_net_1\, B => \sstate[8]_net_1\, S
         => TICK_1(0), Y => \sstate_ns_e[6]\);
    
    \SBYTE[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_30\, CLR => HWRES_c_8, 
        Q => \SBYTE[2]_net_1\);
    
    \DATA[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[9]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[114]\);
    
    \COMMAND[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_5\, CLR => HWRES_c_6, 
        Q => \COMMAND[9]_net_1\);
    
    sstate2se_1_0_0_a2 : NAND2
      port map(A => N_279, B => \sstate2[7]_net_1\, Y => N_109);
    
    \DATA[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[10]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[115]\);
    
    \COMMAND_4_i_m2[15]\ : MUX2H
      port map(A => REG_98, B => \AIR_COMMAND[15]_net_1\, S => 
        RUN_c_0, Y => N_562);
    
    \COMMAND[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_3\, CLR => HWRES_c_5, 
        Q => \COMMAND[2]_net_1\);
    
    REG_1_105_13 : OA21TTF
      port map(A => \REG[105]\, B => sstate_3_sqmuxa, C => N_550, 
        Y => \REG_1_105_13\);
    
    sstate2se_6_i_i_a3 : NAND2
      port map(A => N_279, B => \sstate2_i_0_i[2]\, Y => N_603);
    
    \SBYTE_9[3]\ : MUX2H
      port map(A => \SBYTE[2]_net_1\, B => \COMMAND[11]_net_1\, S
         => N_399, Y => \SBYTE_9[3]_net_1\);
    
    SBYTE_28 : MUX2H
      port map(A => \SBYTE[0]_net_1\, B => \SBYTE_9[0]\, S => 
        N_449, Y => \SBYTE_28\);
    
    \DATA[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[13]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[118]\);
    
    SCL_1_iv_i_a3_0_2 : OR2
      port map(A => \sstate[2]_net_1\, B => \sstate[10]_net_1\, Y
         => SCL_1_iv_i_a3_0);
    
    \COMMAND_4_i_m2[10]\ : MUX2H
      port map(A => REG_93, B => \AIR_COMMAND[10]_net_1\, S => 
        RUN_c_0, Y => N_557);
    
    sstate2se_7_i_i : OAI21FTT
      port map(A => \sstate2_i_0_i[2]\, B => N_279_0, C => N_567, 
        Y => \sstate2se_7_i_i\);
    
    \I2C_RDATA_9_i_a3[7]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[7]_net_1\, Y => 
        N_638);
    
    \I2C_RDATA[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_19\, CLR => 
        HWRES_c_7, Q => \I2C_RDATA[5]_net_1\);
    
    \AIR_COMMAND_19_i_a2_1[1]\ : NOR2
      port map(A => N_577, B => \sstate2[9]_net_1\, Y => N_578);
    
    un1_BITCNT_I_9 : XOR2
      port map(A => \BITCNT[0]_net_1\, B => \un1_scl5_6_0_a2\, Y
         => \DWACT_ADD_CI_0_partial_sum[0]\);
    
    N_513_i_a6_1_2 : AND2
      port map(A => \BITCNT[0]_net_1\, B => \BITCNT[1]_net_1\, Y
         => N_517_2);
    
    \AIR_COMMAND_19_0_iv_0[15]\ : AO21TTF
      port map(A => CHANNEL(2), B => \sstate2[6]_net_1\, C => 
        N_128, Y => \AIR_COMMAND_19[15]\);
    
    un1_BITCNT_I_13 : XOR2
      port map(A => \BITCNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_13);
    
    \I2C_RDATA[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_14\, CLR => 
        HWRES_c_7, Q => \I2C_RDATA[0]_net_1\);
    
    BITCNT_2_sqmuxa_0_a2 : NOR3FTT
      port map(A => TICK_0(0), B => N_395, C => N_397, Y => 
        BITCNT_2_sqmuxa);
    
    un1_scl5_7_0 : NAND3
      port map(A => N_563, B => N_564_i, C => TICK(0), Y => 
        un1_scl5_7);
    
    \COMMAND[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_6\, CLR => HWRES_c_5, 
        Q => \COMMAND[10]_net_1\);
    
    \SBYTE_9[7]\ : MUX2H
      port map(A => \SBYTE[6]_net_1\, B => \COMMAND[15]_net_1\, S
         => N_399, Y => \SBYTE_9[7]_net_1\);
    
    I2C_RDATA_17 : MUX2H
      port map(A => N_589, B => \I2C_RDATA[3]_net_1\, S => N_278, 
        Y => \I2C_RDATA_17\);
    
    un1_scl5_2_i : OAI21
      port map(A => \sstate2[1]_net_1\, B => \sstate2[0]_net_1\, 
        C => TICK_1(0), Y => N_278);
    
    \I2C_RDATA_9_i_a3[9]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[9]_net_1\, Y => 
        N_623);
    
    \I2C_RDATA_9_i[4]\ : OA21TTF
      port map(A => N_594, B => \REG[115]\, C => N_632, Y => 
        N_590);
    
    AIR_COMMAND_37 : MUX2H
      port map(A => N_540, B => \AIR_COMMAND[0]_net_1\, S => 
        un1_scl5_7, Y => \AIR_COMMAND_37\);
    
    N_513_i_a6_0_i_o3 : NAND2
      port map(A => \PULSE_FL\, B => \sstate[13]_net_1\, Y => 
        N_600);
    
    SDAout_m : NOR3FTT
      port map(A => N_600, B => N_454, C => SDAout_m_1_i, Y => 
        SDAout_m_i_i);
    
    N_501_i_a7_1 : AND3
      port map(A => N_517_2, B => \sstate[3]_net_1\, C => 
        \BITCNT[2]_net_1\, Y => N_454);
    
    \DATA[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[11]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[116]\);
    
    AIR_COMMAND_47 : MUX2H
      port map(A => \AIR_COMMAND_19[15]\, B => 
        \AIR_COMMAND[15]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_47\);
    
    \SBYTE[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_33\, CLR => HWRES_c_8, 
        Q => \SBYTE[5]_net_1\);
    
    I2C_RACK_2_0_a3_0_a2 : OR2FT
      port map(A => \sstate2[0]_net_1\, B => N_279_0, Y => 
        I2C_RACK_2);
    
    \COMMAND[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_1\, CLR => HWRES_c_5, 
        Q => \COMMAND[0]_net_1\);
    
    SDAout_12_s : OR3
      port map(A => N_506, B => N_403, C => \un1_sstate_12_0_0_0\, 
        Y => SDAout_12);
    
    \SBYTE_9[1]\ : MUX2H
      port map(A => \SBYTE[0]_net_1\, B => \COMMAND[9]_net_1\, S
         => N_399, Y => \SBYTE_9[1]_net_1\);
    
    SDAnoe_m_1 : AND3FTT
      port map(A => \sstate[9]_net_1\, B => N_581, C => \SDAnoe\, 
        Y => \SDAnoe_m_1\);
    
    COMMAND_8 : MUX2H
      port map(A => \COMMAND[12]_net_1\, B => N_559, S => 
        \sstate[13]_net_1\, Y => \COMMAND_8\);
    
    START_I2C_26 : MUX2H
      port map(A => \START_I2C\, B => N_539, S => TICK(0), Y => 
        \START_I2C_26\);
    
    sstatese_11_i_m2 : MUX2H
      port map(A => \sstate[1]_net_1\, B => \sstate[2]_net_1\, S
         => TICK_2(0), Y => \sstate_ns_e[12]\);
    
    sstatese_7_0_o2 : NAND2
      port map(A => \BITCNT[2]_net_1\, B => N_517_2, Y => N_397);
    
    sstate2se_9_0_a2 : NOR2FT
      port map(A => \sstate2_0[9]_net_1\, B => TICK_0(0), Y => 
        N_113_i);
    
    \I2C_RDATA_9_i[1]\ : OA21TTF
      port map(A => N_595, B => \REG[120]\, C => N_619, Y => 
        N_584);
    
    I2C_RDATA_21 : MUX2H
      port map(A => N_593, B => \I2C_RDATA[7]_net_1\, S => N_278, 
        Y => \I2C_RDATA_21\);
    
    \I2C_RDATA[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_15\, CLR => 
        HWRES_c_7, Q => \I2C_RDATA[1]_net_1\);
    
    \AIR_COMMAND[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_40\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[8]_net_1\);
    
    START_I2C_2_iv_i_a2_0_0 : OR2
      port map(A => \sstate2[8]_net_1\, B => \START_I2C\, Y => 
        \START_I2C_2_iv_i_a2_0_0\);
    
    \sstate2[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2se_2_i_0\, CLR => 
        HWRES_c_10, Q => \sstate2[6]_net_1\);
    
    un1_BITCNT_I_1 : AND2
      port map(A => \BITCNT[0]_net_1\, B => \un1_scl5_6_0_a2\, Y
         => \DWACT_ADD_CI_0_TMP[0]\);
    
    \sstate[13]\ : DFFS
      port map(CLK => CLK_c_c, D => \sstate_ns_e[0]\, SET => 
        HWRES_c_10_0, Q => \sstate[13]_net_1\);
    
    \COMMAND_4_i_m2[13]\ : MUX2H
      port map(A => REG_96, B => \AIR_COMMAND[13]_net_1\, S => 
        RUN_c_0, Y => N_560);
    
    \AIR_COMMAND_19_i_a2[0]\ : NOR2FT
      port map(A => \sstate2_0[9]_net_1\, B => REG_83, Y => N_137);
    
    SDAnoe_m_3 : NOR3FFT
      port map(A => \SDAnoe_m_i\, B => \SDAnoe_m_1\, C => N_454, 
        Y => \SDAnoe_m_3\);
    
    \I2C_RDATA_9_i[5]\ : OA21TTF
      port map(A => N_594, B => \REG[116]\, C => N_634, Y => 
        N_591);
    
    sstate2se_4_i_i : OAI21FTT
      port map(A => \sstate2[5]_net_1\, B => N_279_0, C => N_571, 
        Y => \sstate2se_4_i_i\);
    
    \I2C_RDATA[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_16\, CLR => 
        HWRES_c_7, Q => \I2C_RDATA[2]_net_1\);
    
    AIR_CHAIN : DFFC
      port map(CLK => CLK_c_c, D => \AIR_CHAIN_25\, CLR => 
        HWRES_c_3, Q => \AIR_CHAIN\);
    
    \SCLB_i_a3\ : OR2FT
      port map(A => \CHAIN_SELECT\, B => \SCL\, Y => SCLB_i_a3);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \AIR_COMMAND_19_i[0]\ : OA21TTF
      port map(A => N_144, B => \sstate2_i_0_i[2]\, C => N_137, Y
         => N_540);
    
    un1_sstate_10_0_o2_0_a3_0 : OR2
      port map(A => \COMMAND[0]_net_1\, B => \COMMAND[1]_net_1\, 
        Y => \un1_sstate_10_0_o2_0_a3_0\);
    
    START_I2C_2_iv_i : OA21FTF
      port map(A => \sstate2_0[9]_net_1\, B => 
        \START_I2C_2_iv_i_a2_0_0\, C => N_135, Y => N_539);
    
    \SBYTE_m[7]\ : AND2
      port map(A => \SBYTE[7]_net_1\, B => \sstate[6]_net_1\, Y
         => \SBYTE_m_i[7]\);
    
    SBYTE_34 : MUX2H
      port map(A => \SBYTE[6]_net_1\, B => \SBYTE_9[6]_net_1\, S
         => N_449, Y => \SBYTE_34\);
    
    \I2C_RDATA_9_i[9]\ : OA21TTF
      port map(A => N_594, B => \REG[120]\, C => N_623, Y => 
        N_586);
    
    \COMMAND_m[15]\ : OA21
      port map(A => N_512, B => \sstate[11]_net_1\, C => 
        \COMMAND[15]_net_1\, Y => \COMMAND_m_i[15]\);
    
    \DATA_12[13]\ : MUX2H
      port map(A => \SBYTE[5]_net_1\, B => \REG[118]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[13]_net_1\);
    
    AIR_COMMAND_43 : MUX2H
      port map(A => \AIR_COMMAND_19[11]\, B => 
        \AIR_COMMAND[11]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_43\);
    
    \AIR_COMMAND_19_0_iv_0_o2_0[10]\ : OR2
      port map(A => CHANNEL(1), B => CHANNEL(2), Y => 
        \AIR_COMMAND_19_0_iv_0_o2_0[10]_net_1\);
    
    I2C_RDATA_18 : MUX2H
      port map(A => N_590, B => \I2C_RDATA[4]_net_1\, S => N_278, 
        Y => \I2C_RDATA_18\);
    
    \SBYTE_9_iv_0[0]\ : AO21TTF
      port map(A => N_587, B => \sstate[5]_net_1\, C => N_615, Y
         => \SBYTE_9[0]\);
    
    \COMMAND[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_8\, CLR => HWRES_c_5, 
        Q => \COMMAND[12]_net_1\);
    
    sstatese_8_0_m2 : MUX2H
      port map(A => \sstate[4]_net_1\, B => \sstate[5]_net_1\, S
         => TICK_1(0), Y => \sstate_ns_e[9]\);
    
    \SBYTE[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_34\, CLR => HWRES_c_8, 
        Q => \SBYTE[6]_net_1\);
    
    COMMAND_10 : MUX2H
      port map(A => \COMMAND[14]_net_1\, B => N_561, S => 
        \sstate_0[13]_net_1\, Y => \COMMAND_10\);
    
    \COMMAND[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_9\, CLR => HWRES_c_5, 
        Q => \COMMAND[13]_net_1\);
    
    \AIR_COMMAND_19_0_iv_0[9]\ : AO21TTF
      port map(A => \sstate2[9]_net_1\, B => REG_92, C => N_116, 
        Y => \AIR_COMMAND_19[9]\);
    
    sstate2se_5_i_i_a2 : NAND2
      port map(A => N_279, B => \sstate2[3]_net_1\, Y => N_569);
    
    SBYTE_35 : MUX2H
      port map(A => \SBYTE[7]_net_1\, B => \SBYTE_9[7]_net_1\, S
         => N_449, Y => \SBYTE_35\);
    
    \AIR_COMMAND_19_i_0[1]\ : OA21FTF
      port map(A => \sstate2_0[9]_net_1\, B => REG_84, C => N_578, 
        Y => \AIR_COMMAND_19_i_0_i[1]\);
    
    \BITCNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_8[1]\, CLR => 
        HWRES_c_5, Q => \BITCNT[1]_net_1\);
    
    \I2C_RACK\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RACK_2_i\, CLR => 
        HWRES_c_6, Q => I2C_RACK);
    
    AIR_COMMAND_44 : MUX2H
      port map(A => \AIR_COMMAND_19[12]\, B => 
        \AIR_COMMAND[12]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_44\);
    
    SCL_1_iv_i_o3 : OA21
      port map(A => \sstate_0[13]_net_1\, B => 
        \SCL_1_iv_i_a3_0_1\, C => \SCL\, Y => N_598);
    
    SDAout_del : DFFC
      port map(CLK => CLK_c_c, D => \SDAout\, CLR => HWRES_c_9, Q
         => \SDAout_del\);
    
    I2C_RDATA_22 : MUX2H
      port map(A => N_585, B => \I2C_RDATA[8]_net_1\, S => N_278, 
        Y => \I2C_RDATA_22\);
    
    \I2C_RDATA_9_i[0]\ : OA21TTF
      port map(A => N_595, B => \REG[119]\, C => N_617, Y => 
        N_583);
    
    \sstate[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[9]\, CLR => 
        HWRES_c_11, Q => \sstate[4]_net_1\);
    
    SBYTE_32 : MUX2H
      port map(A => \SBYTE[4]_net_1\, B => \SBYTE_9[4]_net_1\, S
         => N_449, Y => \SBYTE_32\);
    
    \COMMAND_4_i_m2[1]\ : MUX2H
      port map(A => REG_84, B => \AIR_COMMAND[1]_net_1\, S => 
        RUN_c_0_0, Y => N_553);
    
    SBYTE_30 : MUX2H
      port map(A => \SBYTE[2]_net_1\, B => \SBYTE_9[2]_net_1\, S
         => N_449, Y => \SBYTE_30\);
    
    COMMAND_9 : MUX2H
      port map(A => \COMMAND[13]_net_1\, B => N_560, S => 
        \sstate_0[13]_net_1\, Y => \COMMAND_9\);
    
    \sstate2[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2se_3_i_0\, CLR => 
        HWRES_c_9, Q => \sstate2[5]_net_1\);
    
    sstate2se_6_i_i : OAI21FTT
      port map(A => \sstate2[3]_net_1\, B => N_279_0, C => N_603, 
        Y => \sstate2se_6_i_i\);
    
    \SBYTE_9[6]\ : MUX2H
      port map(A => \SBYTE[5]_net_1\, B => \COMMAND[14]_net_1\, S
         => N_399, Y => \SBYTE_9[6]_net_1\);
    
    \DATA[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[8]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[113]\);
    
    COMMAND_5 : MUX2H
      port map(A => \COMMAND[9]_net_1\, B => N_556, S => 
        \sstate[13]_net_1\, Y => \COMMAND_5\);
    
    \SBYTE[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_35\, CLR => HWRES_c_8, 
        Q => \SBYTE[7]_net_1\);
    
    COMMAND_2 : MUX2H
      port map(A => \COMMAND[1]_net_1\, B => N_553, S => 
        \sstate[13]_net_1\, Y => \COMMAND_2\);
    
    \DATA_12_iv_0_a3_0_0[1]\ : NAND2FT
      port map(A => REG_83, B => N_587, Y => 
        \DATA_12_iv_0_a3_0_0_i[1]\);
    
    \sstate[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[2]\, CLR => 
        HWRES_c_10, Q => \sstate[11]_net_1\);
    
    \AIR_COMMAND_19_0_iv_0_0[8]\ : AOI21
      port map(A => \sstate2[9]_net_1\, B => REG_91, C => 
        \sstate2[3]_net_1\, Y => \AIR_COMMAND_19_0_iv_0_0_i[8]\);
    
    \COMMAND[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_11\, CLR => 
        HWRES_c_5, Q => \COMMAND[15]_net_1\);
    
    I2C_RDATA_15 : MUX2H
      port map(A => N_584, B => \I2C_RDATA[1]_net_1\, S => N_278, 
        Y => \I2C_RDATA_15\);
    
    \I2C_RDATA[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_17\, CLR => 
        HWRES_c_7, Q => \I2C_RDATA[3]_net_1\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \sstate[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[10]\, CLR => 
        HWRES_c_10_0, Q => \sstate[3]_net_1\);
    
    \I2C_RDATA[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_18\, CLR => 
        HWRES_c_7, Q => \I2C_RDATA[4]_net_1\);
    
    sstatese_2_0_0 : AO21TTF
      port map(A => \COMMAND[2]_net_1\, B => N_609_1, C => N_608, 
        Y => \sstate_ns_e[3]\);
    
    \sstate[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[13]\, CLR => 
        HWRES_c_10, Q => \sstate[0]_net_1\);
    
    \COMMAND_4_i_m2[9]\ : MUX2H
      port map(A => REG_92, B => \AIR_COMMAND[9]_net_1\, S => 
        RUN_c_0, Y => N_556);
    
    \sstate[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstatese_3_i_m2_i\, CLR => 
        HWRES_c_11, Q => \sstate[9]_net_1\);
    
    un1_scl5_7_0_a2_0 : NAND3FFT
      port map(A => un1_scl5_7_0_a2_0_2_i, B => N_577, C => N_544, 
        Y => N_564_i);
    
    BITCNT_0_sqmuxa_2_0_a2 : OR2FT
      port map(A => TICK_0(0), B => N_400, Y => BITCNT_0_sqmuxa_2);
    
    \I2C_RDATA_9_i_a3[2]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[2]_net_1\, Y => 
        N_628);
    
    \AIR_COMMAND_19_0_iv_0_a2_0_0[10]\ : OR2FT
      port map(A => \sstate2[4]_net_1\, B => \sstate2[6]_net_1\, 
        Y => \AIR_COMMAND_19_0_iv_0_a2_0_i[10]\);
    
    \AIR_COMMAND_19_0_iv_0[8]\ : AO21TTF
      port map(A => N_145, B => 
        \AIR_COMMAND_19_0_iv_0_a2_1[8]_net_1\, C => 
        \AIR_COMMAND_19_0_iv_0_0_i[8]\, Y => \AIR_COMMAND_19[8]\);
    
    sstate2se_2_i_0_a2_0 : NOR2
      port map(A => N_279, B => \sstate2[7]_net_1\, Y => N_108);
    
    \sstate2[9]\ : DFFS
      port map(CLK => CLK_c_c, D => \sstate2_ns_e[0]\, SET => 
        HWRES_c_10, Q => \sstate2[9]_net_1\);
    
    \AIR_COMMAND_19_0_iv_0_a2_0[14]\ : AND2
      port map(A => CHANNEL(1), B => \sstate2[6]_net_1\, Y => 
        N_127_i);
    
    \sstate[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[6]\, CLR => 
        HWRES_c_11, Q => \sstate[7]_net_1\);
    
    sstatese_3_i_m2_i_a3 : NOR2FT
      port map(A => TICK_1(0), B => \sstate[10]_net_1\, Y => 
        N_610);
    
    \I2C_RDATA_9_i[7]\ : OA21TTF
      port map(A => N_594, B => \REG[118]\, C => N_638, Y => 
        N_593);
    
    \sstate2[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2se_7_i_i\, CLR => 
        HWRES_c_9, Q => \sstate2[1]_net_1\);
    
    \DATA[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12_iv[1]\, CLR => 
        HWRES_c_6, Q => \REG[106]\);
    
    \COMMAND_4_i_m2[14]\ : MUX2H
      port map(A => REG_97, B => \AIR_COMMAND[14]_net_1\, S => 
        RUN_c_0, Y => N_561);
    
    START_I2C_2_iv_i_a2 : OA21FTT
      port map(A => \REG_0[105]\, B => \sstate2[0]_net_1\, C => 
        N_145, Y => N_135);
    
    \AIR_COMMAND_19_i[1]\ : OA21FTT
      port map(A => N_145, B => \REG_0[105]\, C => 
        \AIR_COMMAND_19_i_0_i[1]\, Y => N_541);
    
    sstate2se_2_i_0 : OA21FTF
      port map(A => N_279_0, B => \sstate2[6]_net_1\, C => N_108, 
        Y => \sstate2se_2_i_0\);
    
    \I2C_RDATA_9_i[3]\ : OA21TTF
      port map(A => N_594, B => \REG[114]\, C => N_630, Y => 
        N_589);
    
    \DATA[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[14]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[119]\);
    
    un1_BITCNT_I_14 : XOR2
      port map(A => \BITCNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_14);
    
    SCL : DFFS
      port map(CLK => CLK_c_c, D => \SCL_27\, SET => HWRES_c_8, Q
         => \SCL\);
    
    CHAIN_SELECT_4_iv_i_a2 : NOR2FT
      port map(A => RUN_c_0, B => N_551, Y => N_130);
    
    \BITCNT_8_r[1]\ : OA21
      port map(A => BITCNT_2_sqmuxa, B => I_13, C => 
        BITCNT_0_sqmuxa_2, Y => \BITCNT_8[1]\);
    
    PULSE_I2C_i_m2 : MUX2H
      port map(A => PULSE(7), B => \START_I2C\, S => RUN_c_0, Y
         => N_550);
    
    \AIR_COMMAND[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_43\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[11]_net_1\);
    
    BITCNT_2_sqmuxa_0_o2 : NOR2
      port map(A => \sstate[3]_net_1\, B => \sstate[6]_net_1\, Y
         => N_395);
    
    \sstate2[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2_ns_e[2]\, CLR => 
        HWRES_c_10, Q => \sstate2[7]_net_1\);
    
    \sstate[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[12]\, CLR => 
        HWRES_c_10_0, Q => \sstate[1]_net_1\);
    
    AIR_COMMAND_42 : MUX2H
      port map(A => \AIR_COMMAND_19[10]\, B => 
        \AIR_COMMAND[10]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_42\);
    
    \SBYTE[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_29\, CLR => HWRES_c_8, 
        Q => \SBYTE[1]_net_1\);
    
    \DATA_12_iv_0_o3[1]\ : AND2
      port map(A => \sstate[1]_net_1\, B => TICK_1(0), Y => N_597);
    
    \I2C_RDATA[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_21\, CLR => 
        HWRES_c_7_0, Q => \I2C_RDATA[7]_net_1\);
    
    \AIR_COMMAND[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_39\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[2]_net_1\);
    
    SDAin_i_a3 : NOR2FT
      port map(A => \CHAIN_SELECT\, B => SDA1_in, Y => N_626);
    
    \sstate[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[7]\, CLR => 
        HWRES_c_11, Q => \sstate[6]_net_1\);
    
    \sstate2_0[9]\ : DFFS
      port map(CLK => CLK_c_c, D => \sstate2_ns_e[0]\, SET => 
        HWRES_c_10_0, Q => \sstate2_0[9]_net_1\);
    
    \BITCNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_8[2]\, CLR => 
        HWRES_c_5, Q => \BITCNT[2]_net_1\);
    
    sstatese_6_i_m2 : MUX2H
      port map(A => \sstate[6]_net_1\, B => \sstate[7]_net_1\, S
         => TICK_1(0), Y => \sstate_ns_e[7]\);
    
    sstatese_4_0_a2_0 : NAND3
      port map(A => TICK_2(0), B => N_397, C => \sstate[6]_net_1\, 
        Y => N_436);
    
    \AIR_COMMAND_19_0_iv_0_o2[8]\ : NAND2
      port map(A => \sstate2[5]_net_1\, B => \REG[105]\, Y => 
        N_548);
    
    \sstate_0[13]\ : DFFS
      port map(CLK => CLK_c_c, D => \sstate_ns_e[0]\, SET => 
        HWRES_c_10_0, Q => \sstate_0[13]_net_1\);
    
    SDAin_i : OA21TTF
      port map(A => \CHAIN_SELECT\, B => SDA0_in, C => N_626, Y
         => N_587);
    
    \BITCNT_8_r[2]\ : OA21
      port map(A => BITCNT_2_sqmuxa, B => I_14, C => 
        BITCNT_0_sqmuxa_2, Y => \BITCNT_8[2]\);
    
    \AIR_COMMAND_19_0_iv_0[11]\ : AO21TTF
      port map(A => \sstate2[9]_net_1\, B => REG_94, C => N_121, 
        Y => \AIR_COMMAND_19[11]\);
    
    \DATA[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[15]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[120]\);
    
    SBYTE_33 : MUX2H
      port map(A => \SBYTE[5]_net_1\, B => \SBYTE_9[5]_net_1\, S
         => N_449, Y => \SBYTE_33\);
    
    AIR_CHAIN_4_iv_i : OA21TTF
      port map(A => N_544, B => REG_0, C => \AIR_CHAIN_4_iv_i_0\, 
        Y => N_538);
    
    \AIR_COMMAND_19_0_iv_0[13]\ : AO21TTF
      port map(A => CHANNEL(0), B => \sstate2[6]_net_1\, C => 
        N_124, Y => \AIR_COMMAND_19[13]\);
    
    un1_SDAnoe_0_sqmuxa_0_o2_0 : NOR2
      port map(A => \sstate[6]_net_1\, B => \sstate[7]_net_1\, Y
         => N_402);
    
    sstatese_7_0_0 : OA21FTT
      port map(A => \sstate[5]_net_1\, B => TICK_0(0), C => N_432, 
        Y => \sstatese_7_0_0\);
    
    SBYTE_31 : MUX2H
      port map(A => \SBYTE[3]_net_1\, B => \SBYTE_9[3]_net_1\, S
         => N_449, Y => \SBYTE_31\);
    
    \I2C_RDATA_9_i_a3[4]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[4]_net_1\, Y => 
        N_632);
    
    \COMMAND[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_10\, CLR => 
        HWRES_c_5, Q => \COMMAND[14]_net_1\);
    
    \AIR_COMMAND_19_0_iv_0_a2[14]\ : AND2
      port map(A => \sstate2_0[9]_net_1\, B => REG_97, Y => 
        N_126_i);
    
    \DATA_12_iv_0[1]\ : MUX2H
      port map(A => \REG[106]\, B => \DATA_12_iv_0_a3_0_0_i[1]\, 
        S => N_597, Y => \DATA_12_iv[1]\);
    
    \AIR_COMMAND_19_0_iv_0_o2[12]\ : NAND2FT
      port map(A => N_543, B => N_548, Y => N_545_i_i);
    
    \AIR_COMMAND_19_0_iv_0_a2_1_0[10]\ : OAI21
      port map(A => CHANNEL(0), B => 
        \AIR_COMMAND_19_0_iv_0_o2_0[10]_net_1\, C => \REG[105]\, 
        Y => \AIR_COMMAND_19_0_iv_0_a2_1_i[10]\);
    
    N_279_i_i_o2_0_o3 : NAND2
      port map(A => \REG_0[105]\, B => TICK_2(0), Y => N_279);
    
    sstatese_12_i_m2 : MUX2H
      port map(A => \sstate[0]_net_1\, B => \sstate[1]_net_1\, S
         => TICK_2(0), Y => \sstate_ns_e[13]\);
    
    SDAout_m_1 : NAND3
      port map(A => \SDAnoe_m_i\, B => N_581, C => \SDAout\, Y
         => SDAout_m_1_i);
    
    sstatese_1_i_m2 : MUX2H
      port map(A => \sstate[11]_net_1\, B => \sstate[12]_net_1\, 
        S => TICK_1(0), Y => \sstate_ns_e[2]\);
    
    \SCLA_i_a3\ : OR2
      port map(A => \CHAIN_SELECT\, B => \SCL\, Y => SCLA_i_a3);
    
    I2C_RACK_2_i : INV
      port map(A => I2C_RACK_2, Y => \I2C_RACK_2_i\);
    
    \DATA_12[10]\ : MUX2H
      port map(A => \SBYTE[2]_net_1\, B => \REG[115]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[10]_net_1\);
    
    \AIR_COMMAND[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_45\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[13]_net_1\);
    
    \I2C_RDATA_9_i_o3_0[8]\ : NAND2
      port map(A => \sstate2[1]_net_1\, B => \REG_0[105]\, Y => 
        N_594_0);
    
    \AIR_COMMAND_19_i_0[2]\ : OAI21FTF
      port map(A => \sstate2_0[9]_net_1\, B => REG_85, C => N_143, 
        Y => \AIR_COMMAND_19_i_0[2]_net_1\);
    
    sstatese_4_0_0 : OA21FTT
      port map(A => \sstate[8]_net_1\, B => TICK_0(0), C => N_436, 
        Y => \sstatese_4_0_0\);
    
    SCL_1_iv_i_a3_0_1 : OR3
      port map(A => \sstate[11]_net_1\, B => \sstate[9]_net_1\, C
         => \sstate[0]_net_1\, Y => \SCL_1_iv_i_a3_0_1\);
    
    \I2C_RDATA_9_i_a3[5]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[5]_net_1\, Y => 
        N_634);
    
    sstatese_2_0_0_a3_0_1 : AND2
      port map(A => \sstate[0]_net_1\, B => TICK_2(0), Y => 
        N_609_1);
    
    \sstate2[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2se_6_i_i\, CLR => 
        HWRES_c_9, Q => \sstate2_i_0_i[2]\);
    
    \I2C_RDATA_9_i_a3[3]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[3]_net_1\, Y => 
        N_630);
    
    \AIR_COMMAND_19_0_iv_0_a2[11]\ : NAND2
      port map(A => CHIP_ADDR(2), B => N_545_i_i, Y => N_121);
    
    \sstate2[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2se_8_i_i\, CLR => 
        HWRES_c_9, Q => \sstate2[0]_net_1\);
    
    I2C_RDATA_16 : MUX2H
      port map(A => N_588, B => \I2C_RDATA[2]_net_1\, S => N_278, 
        Y => \I2C_RDATA_16\);
    
    \AIR_COMMAND_19_0_iv_0_a2[10]\ : NAND3FFT
      port map(A => \AIR_COMMAND_19_0_iv_0_a2_1_i[10]\, B => 
        \AIR_COMMAND_19_0_iv_0_a2_0_i[10]\, C => N_578, Y => 
        N_118_i);
    
    \SBYTE[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_28\, CLR => HWRES_c_8, 
        Q => \SBYTE[0]_net_1\);
    
    \AIR_COMMAND_19_i_a2_1[0]\ : OR2
      port map(A => \sstate2_0[9]_net_1\, B => \sstate2[1]_net_1\, 
        Y => N_144);
    
    AIR_CHAIN_4_iv_i_a2_0 : NOR2
      port map(A => N_133_1, B => I2C_CHAIN, Y => N_133);
    
    \COMMAND[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_7\, CLR => HWRES_c_5, 
        Q => \COMMAND[11]_net_1\);
    
    BITCNT_0_sqmuxa_2_0_o2 : OA21FTF
      port map(A => N_398, B => N_600, C => \sstate[11]_net_1\, Y
         => N_400);
    
    \COMMAND[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_2\, CLR => HWRES_c_5, 
        Q => \COMMAND[1]_net_1\);
    
    sstate2se_8_i_i_a2 : NAND2
      port map(A => N_279, B => \sstate2[0]_net_1\, Y => N_565);
    
    \I2C_RDATA[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_22\, CLR => 
        HWRES_c_7_0, Q => \I2C_RDATA[8]_net_1\);
    
    sstate2se_8_i_i : OAI21FTT
      port map(A => \sstate2[1]_net_1\, B => N_279_0, C => N_565, 
        Y => \sstate2se_8_i_i\);
    
    COMMAND_4 : MUX2H
      port map(A => \COMMAND[8]_net_1\, B => N_555, S => 
        \sstate[13]_net_1\, Y => \COMMAND_4\);
    
    \I2C_RDATA_9_i_a3[1]\ : NOR2FT
      port map(A => N_595, B => \I2C_RDATA[1]_net_1\, Y => N_619);
    
    \sstate2[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2se_5_i_i\, CLR => 
        HWRES_c_9, Q => \sstate2[3]_net_1\);
    
    \SBYTE_9[2]\ : MUX2H
      port map(A => \SBYTE[1]_net_1\, B => \COMMAND[10]_net_1\, S
         => N_399, Y => \SBYTE_9[2]_net_1\);
    
    sstatese_7_0 : AO21TTF
      port map(A => N_457, B => TICK_2(0), C => \sstatese_7_0_0\, 
        Y => \sstate_ns_e[8]\);
    
    \REG_1_0[105]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_105_13\, SET => 
        HWRES_c_7_0, Q => \REG_0[105]\);
    
    BITCNT_0_sqmuxa_2_0_o2_0 : NAND2FT
      port map(A => \COMMAND[0]_net_1\, B => \COMMAND[1]_net_1\, 
        Y => N_398);
    
    sstatese_7_0_a2_2_0_a3 : NOR2FT
      port map(A => \COMMAND[0]_net_1\, B => N_600, Y => N_457);
    
    \DATA_12[9]\ : MUX2H
      port map(A => \SBYTE[1]_net_1\, B => \REG[114]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[9]_net_1\);
    
    \sstate[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[3]\, CLR => 
        HWRES_c_10, Q => \sstate[10]_net_1\);
    
    SDAout_12_iv : OR3
      port map(A => SDAout_m_i_i, B => \COMMAND_m_i[15]\, C => 
        \SBYTE_m_i[7]\, Y => N_506);
    
    \SBYTE_9_iv_0_a3[0]\ : NAND2
      port map(A => \COMMAND[8]_net_1\, B => N_399, Y => N_615);
    
    sstatese_0_0 : OAI21FTT
      port map(A => \sstate[12]_net_1\, B => TICK_0(0), C => 
        N_441, Y => \sstate_ns_e[1]\);
    
    sstate2se_4_i_i_a2 : NAND2
      port map(A => N_279, B => \sstate2[4]_net_1\, Y => N_571);
    
    \AIR_COMMAND_19_0_iv_0[12]\ : AO21
      port map(A => \sstate2[9]_net_1\, B => REG_95, C => 
        N_545_i_i, Y => \AIR_COMMAND_19[12]\);
    
    \COMMAND_4_i_m2[2]\ : MUX2H
      port map(A => REG_85, B => \AIR_COMMAND[2]_net_1\, S => 
        RUN_c_0_0, Y => N_554);
    
    \I2C_RDATA_9_i[8]\ : OA21TTF
      port map(A => N_594, B => \REG[119]\, C => N_621, Y => 
        N_585);
    
    sstatese_9_i_m2 : MUX2H
      port map(A => \sstate[3]_net_1\, B => \sstate[4]_net_1\, S
         => TICK_1(0), Y => \sstate_ns_e[10]\);
    
    \REG_1[105]\ : DFFS
      port map(CLK => CLK_c_c, D => \REG_1_105_13\, SET => 
        HWRES_c_7_0, Q => \REG[105]\);
    
    \AIR_COMMAND[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_38\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[1]_net_1\);
    
    sstatese_7_0_a2 : NAND3
      port map(A => TICK_2(0), B => N_397, C => \sstate[3]_net_1\, 
        Y => N_432);
    
    \AIR_COMMAND_19_0_iv_0_0[10]\ : AOI21TTF
      port map(A => \sstate2[9]_net_1\, B => REG_93, C => N_118_i, 
        Y => \AIR_COMMAND_19_0_iv_0_0[10]_net_1\);
    
    AIR_COMMAND_45 : MUX2H
      port map(A => \AIR_COMMAND_19[13]\, B => 
        \AIR_COMMAND[13]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_45\);
    
    SBYTE_29 : MUX2H
      port map(A => \SBYTE[1]_net_1\, B => \SBYTE_9[1]_net_1\, S
         => N_449, Y => \SBYTE_29\);
    
    \I2C_RDATA_9_i[2]\ : OA21TTF
      port map(A => N_594, B => \REG[113]\, C => N_628, Y => 
        N_588);
    
    \AIR_COMMAND_19_0_iv_0[10]\ : AO21TTF
      port map(A => CHIP_ADDR(1), B => N_545_i_i, C => 
        \AIR_COMMAND_19_0_iv_0_0[10]_net_1\, Y => 
        \AIR_COMMAND_19[10]\);
    
    un1_scl5_7_0_a2_0_2 : NOR2
      port map(A => \sstate2_i_0_i[2]\, B => \sstate2[7]_net_1\, 
        Y => un1_scl5_7_0_a2_0_0);
    
    I2C_RDATA_20 : MUX2H
      port map(A => N_592, B => \I2C_RDATA[6]_net_1\, S => N_278, 
        Y => \I2C_RDATA_20\);
    
    \sstate[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[5]\, CLR => 
        HWRES_c_11, Q => \sstate[8]_net_1\);
    
    \I2C_RDATA[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_23\, CLR => 
        HWRES_c_7_0, Q => \I2C_RDATA[9]_net_1\);
    
    sstate2se_1_0_0 : AO21TTF
      port map(A => \sstate2[8]_net_1\, B => TICK_2(0), C => 
        N_109, Y => \sstate2_ns_e[2]\);
    
    \AIR_COMMAND[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_42\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[10]_net_1\);
    
    COMMAND_11 : MUX2H
      port map(A => \COMMAND[15]_net_1\, B => N_562, S => 
        \sstate_0[13]_net_1\, Y => \COMMAND_11\);
    
    sstate2se_5_i_i : OAI21FTT
      port map(A => \sstate2[4]_net_1\, B => N_279_0, C => N_569, 
        Y => \sstate2se_5_i_i\);
    
    \AIR_COMMAND_19_i_a2_1[2]\ : NOR2
      port map(A => N_144, B => N_564_1, Y => N_143);
    
    \sstate[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[11]\, CLR => 
        HWRES_c_10_0, Q => \sstate[2]_net_1\);
    
    \I2C_RDATA[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \I2C_RDATA_20\, CLR => 
        HWRES_c_7_0, Q => \I2C_RDATA[6]_net_1\);
    
    AIR_COMMAND_46 : MUX2H
      port map(A => \AIR_COMMAND_19[14]\, B => 
        \AIR_COMMAND[14]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_46\);
    
    \sstate[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[8]\, CLR => 
        HWRES_c_11, Q => \sstate[5]_net_1\);
    
    SDAout_del1 : DFFC
      port map(CLK => CLK_c_c, D => \SDAout_del\, CLR => 
        HWRES_c_9, Q => \SDAout_del1\);
    
    \sstate2[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate2_ns_e[1]\, CLR => 
        HWRES_c_10, Q => \sstate2[8]_net_1\);
    
    \AIR_COMMAND[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_37\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[0]_net_1\);
    
    un1_scl5_4_0_a2_0_a3 : AOI21FTF
      port map(A => N_399, B => N_596, C => TICK(0), Y => N_449);
    
    \I2C_RDATA_9_i_o3[8]\ : NAND2
      port map(A => \sstate2[1]_net_1\, B => \REG[105]\, Y => 
        N_594);
    
    SCL_1_iv_i_a3 : NAND3FFT
      port map(A => N_598, B => SCL_1_iv_i_a3_0, C => N_596, Y
         => N_612);
    
    AIR_COMMAND_38 : MUX2H
      port map(A => N_541, B => \AIR_COMMAND[1]_net_1\, S => 
        un1_scl5_7, Y => \AIR_COMMAND_38\);
    
    AIR_CHAIN_25 : MUX2H
      port map(A => \AIR_CHAIN\, B => N_538, S => TICK(0), Y => 
        \AIR_CHAIN_25\);
    
    \sstate[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns_e[1]\, CLR => 
        HWRES_c_10_0, Q => \sstate[12]_net_1\);
    
    AIR_CHAIN_4_iv_i_a2_0_1 : NAND2
      port map(A => \sstate2[9]_net_1\, B => I2C_RREQ, Y => 
        N_133_1);
    
    un1_sstate_12_0_0_o3 : OAI21TTF
      port map(A => N_397, B => N_402, C => N_457, Y => N_403);
    
    sstate2se_7_i_i_a2 : NAND2
      port map(A => N_279, B => \sstate2[1]_net_1\, Y => N_567);
    
    \I2C_RDATA_9_i_a3[6]\ : NOR2FT
      port map(A => N_594_0, B => \I2C_RDATA[6]_net_1\, Y => 
        N_636);
    
    AIR_COMMAND_39 : MUX2H
      port map(A => N_542, B => \AIR_COMMAND[2]_net_1\, S => 
        un1_scl5_7, Y => \AIR_COMMAND_39\);
    
    \AIR_COMMAND_19_0_iv_0_a2[15]\ : NAND2
      port map(A => \sstate2_0[9]_net_1\, B => REG_98, Y => N_128);
    
    un1_BITCNT_I_15 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \BITCNT[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \I2C_RDATA_9_i_o3[0]\ : OR2FT
      port map(A => \REG_0[105]\, B => \sstate2[1]_net_1\, Y => 
        N_595);
    
    \COMMAND_4_i_m2[0]\ : MUX2H
      port map(A => REG_83, B => \AIR_COMMAND[0]_net_1\, S => 
        RUN_c_0_0, Y => N_552);
    
    \AIR_COMMAND[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_44\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[12]_net_1\);
    
    un1_scl5_6_0_a2 : AOI21TTF
      port map(A => N_400, B => N_395, C => TICK_1(0), Y => 
        \un1_scl5_6_0_a2\);
    
    un1_scl5_7_0_a2 : OR3FTT
      port map(A => N_544, B => \REG_0[105]\, C => 
        \sstate2[8]_net_1\, Y => N_563);
    
    \SBYTE_9[5]\ : MUX2H
      port map(A => \SBYTE[4]_net_1\, B => \COMMAND[13]_net_1\, S
         => N_399, Y => \SBYTE_9[5]_net_1\);
    
    SDAout_36 : MUX2H
      port map(A => \SDAout\, B => SDAout_12, S => TICK(0), Y => 
        \SDAout_36\);
    
    DATA_1_sqmuxa_2_0_a2 : NAND2
      port map(A => N_454, B => TICK(0), Y => DATA_1_sqmuxa_2_i);
    
    \DATA_12[11]\ : MUX2H
      port map(A => \SBYTE[3]_net_1\, B => \REG[116]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[11]_net_1\);
    
    \BITCNT_8_r[0]\ : OA21
      port map(A => BITCNT_2_sqmuxa, B => 
        \DWACT_ADD_CI_0_partial_sum[0]\, C => BITCNT_0_sqmuxa_2, 
        Y => \BITCNT_8[0]\);
    
    PULSE_FL : DFFC
      port map(CLK => CLK_c_c, D => \PULSE_FL_12\, CLR => 
        HWRES_c_7_0, Q => \PULSE_FL\);
    
    sstate2se_9_0 : NAND3FTT
      port map(A => N_113_i, B => I2C_RACK_2, C => N_544, Y => 
        \sstate2_ns_e[0]\);
    
    I2C_RDATA_19 : MUX2H
      port map(A => N_591, B => \I2C_RDATA[5]_net_1\, S => N_278, 
        Y => \I2C_RDATA_19\);
    
    \SBYTE[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \SBYTE_31\, CLR => HWRES_c_8, 
        Q => \SBYTE[3]_net_1\);
    
    I2C_RDATA_23 : MUX2H
      port map(A => N_586, B => \I2C_RDATA[9]_net_1\, S => N_278, 
        Y => \I2C_RDATA_23\);
    
    un1_sstate_10_0_o2_0_o3 : OAI21TTF
      port map(A => \un1_sstate_10_0_o2_0_a3_0\, B => N_600, C
         => \sstate[11]_net_1\, Y => N_399);
    
    sstate2se_0_0_0_a2 : OR2FT
      port map(A => \sstate2[8]_net_1\, B => TICK_0(0), Y => 
        N_111);
    
    SDAnoe_del2 : DFFC
      port map(CLK => CLK_c_c, D => \SDAnoe_del1\, CLR => 
        HWRES_c_9, Q => \SDAnoe_del2\);
    
    \AIR_COMMAND[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \AIR_COMMAND_41\, CLR => 
        HWRES_c_4, Q => \AIR_COMMAND[9]_net_1\);
    
    \SDAout_del2\ : DFFC
      port map(CLK => CLK_c_c, D => \SDAout_del1\, CLR => 
        HWRES_c_9, Q => SDAout_del2);
    
    I2C_RDATA_14 : MUX2H
      port map(A => N_583, B => \I2C_RDATA[0]_net_1\, S => N_278, 
        Y => \I2C_RDATA_14\);
    
    N_513_i_a6_i : NAND2
      port map(A => \COMMAND[2]_net_1\, B => \sstate[0]_net_1\, Y
         => N_581);
    
    SDAnoe_m_i : NOR2
      port map(A => \sstate[11]_net_1\, B => \sstate[6]_net_1\, Y
         => \SDAnoe_m_i\);
    
    \DATA_12[14]\ : MUX2H
      port map(A => \SBYTE[6]_net_1\, B => \REG[119]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[14]_net_1\);
    
    N_511_a3 : NOR3FFT
      port map(A => \sstate_0[13]_net_1\, B => \PULSE_FL\, C => 
        \COMMAND[1]_net_1\, Y => N_512);
    
    \un1_sdab_i\ : NOR2FT
      port map(A => \CHAIN_SELECT\, B => \SDAnoe_del2\, Y => 
        un1_sdab_i);
    
    sstatese_4_0 : AO21TTF
      port map(A => N_399, B => TICK_2(0), C => \sstatese_4_0_0\, 
        Y => \sstate_ns_e[5]\);
    
    COMMAND_1 : MUX2H
      port map(A => \COMMAND[0]_net_1\, B => N_552, S => 
        \sstate[13]_net_1\, Y => \COMMAND_1\);
    
    SDAout : DFFS
      port map(CLK => CLK_c_c, D => \SDAout_36\, SET => HWRES_c_9, 
        Q => \SDAout\);
    
    sstatese_10_0 : OAI21FTF
      port map(A => \sstate[2]_net_1\, B => TICK_0(0), C => 
        BITCNT_2_sqmuxa, Y => \sstate_ns_e[11]\);
    
    \AIR_COMMAND_19_0_iv_0_a2[13]\ : NAND2
      port map(A => \sstate2_0[9]_net_1\, B => REG_96, Y => N_124);
    
    \un1_sdaa_0_a3\ : NOR2
      port map(A => \CHAIN_SELECT\, B => \SDAnoe_del2\, Y => 
        un1_sdaa_0_a3);
    
    CHAIN_SELECT_24 : MUX2H
      port map(A => \CHAIN_SELECT\, B => N_537, S => 
        \sstate_0[13]_net_1\, Y => \CHAIN_SELECT_24\);
    
    sstatese_3_i_m2_i : OA21TTF
      port map(A => \sstate[9]_net_1\, B => TICK_1(0), C => N_610, 
        Y => \sstatese_3_i_m2_i\);
    
    PULSE_FL_12 : AO21
      port map(A => \PULSE_FL\, B => \sstate_0[13]_net_1\, C => 
        N_550, Y => \PULSE_FL_12\);
    
    \COMMAND_4_i_m2[8]\ : MUX2H
      port map(A => REG_91, B => \AIR_COMMAND[8]_net_1\, S => 
        RUN_c_0_0, Y => N_555);
    
    sstate2se_3_i_0 : OA21TTF
      port map(A => N_279, B => \sstate2[6]_net_1\, C => N_573, Y
         => \sstate2se_3_i_0\);
    
    \COMMAND[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \COMMAND_4\, CLR => HWRES_c_6, 
        Q => \COMMAND[8]_net_1\);
    
    N_279_i_i_o2_0_o3_0 : NAND2
      port map(A => \REG_0[105]\, B => TICK_0(0), Y => N_279_0);
    
    sstatese_13 : AO21FTF
      port map(A => \COMMAND[2]_net_1\, B => N_609_1, C => 
        \sstatese_13_0\, Y => \sstate_ns_e[0]\);
    
    \AIR_COMMAND_19_0_iv_0_a2[9]\ : NAND2
      port map(A => CHIP_ADDR(0), B => N_545_i_i, Y => N_116);
    
    un1_scl5_7_0_a2_0_4 : OR3FTT
      port map(A => un1_scl5_7_0_a2_0_0, B => \sstate2[1]_net_1\, 
        C => N_564_1, Y => un1_scl5_7_0_a2_0_2_i);
    
    \DATA[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \DATA_12[12]_net_1\, CLR => 
        HWRES_c_6, Q => \REG[117]\);
    
    \DATA_12[8]\ : MUX2H
      port map(A => \SBYTE[0]_net_1\, B => \REG[113]\, S => 
        DATA_1_sqmuxa_2_i, Y => \DATA_12[8]_net_1\);
    
    COMMAND_7 : MUX2H
      port map(A => \COMMAND[11]_net_1\, B => N_558, S => 
        \sstate[13]_net_1\, Y => \COMMAND_7\);
    
    AIR_COMMAND_41 : MUX2H
      port map(A => \AIR_COMMAND_19[9]\, B => 
        \AIR_COMMAND[9]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_41\);
    
    SDAnoe_8_s : AO21
      port map(A => N_600, B => \SDAnoe_m_3\, C => N_403, Y => 
        SDAnoe_8);
    
    CHAIN_SELECT_4_iv_i : OA21TTF
      port map(A => REG_0, B => RUN_c_0, C => N_130, Y => N_537);
    
    sstate_3_sqmuxa_0_a2 : NOR2FT
      port map(A => \sstate_0[13]_net_1\, B => \PULSE_FL\, Y => 
        sstate_3_sqmuxa);
    
    COMMAND_3 : MUX2H
      port map(A => \COMMAND[2]_net_1\, B => N_554, S => 
        \sstate[13]_net_1\, Y => \COMMAND_3\);
    
    AIR_COMMAND_40 : MUX2H
      port map(A => \AIR_COMMAND_19[8]\, B => 
        \AIR_COMMAND[8]_net_1\, S => un1_scl5_7, Y => 
        \AIR_COMMAND_40\);
    
    sstatese_2_0_0_a3 : OR2FT
      port map(A => \sstate[10]_net_1\, B => TICK_0(0), Y => 
        N_608);
    
    SCL_27 : MUX2H
      port map(A => \SCL\, B => N_612, S => TICK(0), Y => 
        \SCL_27\);
    
    SCL_1_iv_i_o3_0 : NOR2
      port map(A => \sstate[5]_net_1\, B => \sstate[8]_net_1\, Y
         => N_596);
    
    COMMAND_6 : MUX2H
      port map(A => \COMMAND[10]_net_1\, B => N_557, S => 
        \sstate[13]_net_1\, Y => \COMMAND_6\);
    
    CHAIN_SELECT_4_iv_i_m2 : MUX2H
      port map(A => \CHAIN_SELECT\, B => \AIR_CHAIN\, S => 
        I2C_RREQ, Y => N_551);
    
    CHAIN_SELECT : DFFC
      port map(CLK => CLK_c_c, D => \CHAIN_SELECT_24\, CLR => 
        HWRES_c_5, Q => \CHAIN_SELECT\);
    
    sstatese_13_0 : AOI21TTF
      port map(A => \sstate[9]_net_1\, B => TICK_2(0), C => N_442, 
        Y => \sstatese_13_0\);
    
    \AIR_COMMAND_19_0_iv_0_a2_1[8]\ : NOR2
      port map(A => \sstate2[8]_net_1\, B => \sstate2[9]_net_1\, 
        Y => N_145);
    
    sstate2se_3_i_0_a2 : NOR2FT
      port map(A => N_279_0, B => \sstate2[5]_net_1\, Y => N_573);
    
    SDAnoe_48 : MUX2H
      port map(A => \SDAnoe\, B => SDAnoe_8, S => TICK(0), Y => 
        \SDAnoe_48\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity MONOSTABLE_3 is

    port( LEDint     : out   std_logic_vector(2 to 2);
          TICK_0     : in    std_logic_vector(2 to 2);
          CLK_c_c    : in    std_logic;
          HWRES_c_33 : in    std_logic;
          TMONOS     : in    std_logic
        );

end MONOSTABLE_3;

architecture DEF_ARCH of MONOSTABLE_3 is 

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_36, \LEDint[2]\, \GND\, \VCC\ : std_logic;

begin 

    LEDint(2) <= \LEDint[2]\;

    PWR_i : PWR
      port map(Y => \VCC\);
    
    MONOUT : DFFC
      port map(CLK => CLK_c_c, D => N_36, CLR => HWRES_c_33, Q
         => \LEDint[2]\);
    
    MONOUT_0_i : OA21FTT
      port map(A => TICK_0(2), B => TMONOS, C => \LEDint[2]\, Y
         => N_36);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity MONOSTABLE_2 is

    port( TICK_0     : in    std_logic_vector(2 to 2);
          CLK_c_c    : in    std_logic;
          HWRES_c_33 : in    std_logic;
          TMONOS     : out   std_logic
        );

end MONOSTABLE_2;

architecture DEF_ARCH of MONOSTABLE_2 is 

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal TMONOS_0_0_a2_1, TMONOS_net_1, \GND\, \VCC\
         : std_logic;

begin 

    TMONOS <= TMONOS_net_1;

    TMONOS_0_0_a2 : NOR2FT
      port map(A => TMONOS_net_1, B => TICK_0(2), Y => 
        TMONOS_0_0_a2_1);
    
    \TMONOS\ : DFFC
      port map(CLK => CLK_c_c, D => TMONOS_0_0_a2_1, CLR => 
        HWRES_c_33, Q => TMONOS_net_1);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity MONOSTABLE_1 is

    port( LEDint       : out   std_logic_vector(1 to 1);
          TICK_0       : in    std_logic_vector(2 to 2);
          PULSE        : in    std_logic_vector(2 to 2);
          HWRES_c_33   : in    std_logic;
          CLK_c_c      : in    std_logic;
          HWRES_c_32_0 : in    std_logic;
          EVNT_TRG     : in    std_logic
        );

end MONOSTABLE_1;

architecture DEF_ARCH of MONOSTABLE_1 is 

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_792_i_0, N_39, \TMONOS\, TMONOS_0_0_a2_0, 
        \LEDint[1]\, \GND\, \VCC\ : std_logic;

begin 

    LEDint(1) <= \LEDint[1]\;

    TMONOS_0_0_a2 : NOR2FT
      port map(A => \TMONOS\, B => TICK_0(2), Y => 
        TMONOS_0_0_a2_0);
    
    TMONOS : DFFB
      port map(CLK => CLK_c_c, D => TMONOS_0_0_a2_0, CLR => 
        HWRES_c_33, SET => N_792_i_0, Q => \TMONOS\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    MONOUT : DFFB
      port map(CLK => CLK_c_c, D => N_39, CLR => HWRES_c_32_0, 
        SET => N_792_i_0, Q => \LEDint[1]\);
    
    MONOUT_0_i : OA21FTT
      port map(A => TICK_0(2), B => \TMONOS\, C => \LEDint[1]\, Y
         => N_39);
    
    TMONOS_i_0 : OR2
      port map(A => EVNT_TRG, B => PULSE(2), Y => N_792_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity MONOSTABLE is

    port( LEDint       : out   std_logic_vector(0 to 0);
          TICK_0       : in    std_logic_vector(2 to 2);
          CLK_c_c      : in    std_logic;
          RUN_c        : in    std_logic;
          HWRES_c_32_0 : in    std_logic
        );

end MONOSTABLE;

architecture DEF_ARCH of MONOSTABLE is 

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_42, \TMONOS\, \TMONOS_0_0_a2\, \LEDint[0]\, \GND\, 
        \VCC\ : std_logic;

begin 

    LEDint(0) <= \LEDint[0]\;

    TMONOS_0_0_a2 : NOR2FT
      port map(A => \TMONOS\, B => TICK_0(2), Y => 
        \TMONOS_0_0_a2\);
    
    TMONOS : DFFB
      port map(CLK => CLK_c_c, D => \TMONOS_0_0_a2\, CLR => 
        HWRES_c_32_0, SET => RUN_c, Q => \TMONOS\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    MONOUT : DFFB
      port map(CLK => CLK_c_c, D => N_42, CLR => HWRES_c_32_0, 
        SET => RUN_c, Q => \LEDint[0]\);
    
    MONOUT_0_i : OA21FTT
      port map(A => TICK_0(2), B => \TMONOS\, C => \LEDint[0]\, Y
         => N_42);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity MONOSTABLE_4 is

    port( LEDint     : out   std_logic_vector(4 to 4);
          TICK_0     : in    std_logic_vector(2 to 2);
          TST_c_c    : in    std_logic_vector(3 to 3);
          CLK_c_c    : in    std_logic;
          HWRES_c_33 : in    std_logic
        );

end MONOSTABLE_4;

architecture DEF_ARCH of MONOSTABLE_4 is 

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \TST_c_c_i_0[3]\, N_33, \TMONOS\, TMONOS_0_0_a2_2, 
        \LEDint[4]\, \GND\, \VCC\ : std_logic;

begin 

    LEDint(4) <= \LEDint[4]\;

    TMONOS_0_0_a2 : NOR2FT
      port map(A => \TMONOS\, B => TICK_0(2), Y => 
        TMONOS_0_0_a2_2);
    
    TMONOS : DFFB
      port map(CLK => CLK_c_c, D => TMONOS_0_0_a2_2, CLR => 
        HWRES_c_33, SET => \TST_c_c_i_0[3]\, Q => \TMONOS\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    MONOUT : DFFB
      port map(CLK => CLK_c_c, D => N_33, CLR => HWRES_c_33, SET
         => \TST_c_c_i_0[3]\, Q => \LEDint[4]\);
    
    MONOUT_0_i : OA21FTT
      port map(A => TICK_0(2), B => \TMONOS\, C => \LEDint[4]\, Y
         => N_33);
    
    TMONOS_i_0 : INV
      port map(A => TST_c_c(3), Y => \TST_c_c_i_0[3]\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity MONOSTABLE_5 is

    port( LEDint     : out   std_logic_vector(5 to 5);
          TICK_0     : in    std_logic_vector(2 to 2);
          CLK_c_c    : in    std_logic;
          HWRES_c_33 : in    std_logic;
          nLBRDY_c   : in    std_logic
        );

end MONOSTABLE_5;

architecture DEF_ARCH of MONOSTABLE_5 is 

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal nLBRDY_c_i_0, N_30, \TMONOS\, TMONOS_0_0_a2_3, 
        \LEDint[5]\, \GND\, \VCC\ : std_logic;

begin 

    LEDint(5) <= \LEDint[5]\;

    TMONOS_0_0_a2 : NOR2FT
      port map(A => \TMONOS\, B => TICK_0(2), Y => 
        TMONOS_0_0_a2_3);
    
    TMONOS : DFFB
      port map(CLK => CLK_c_c, D => TMONOS_0_0_a2_3, CLR => 
        HWRES_c_33, SET => nLBRDY_c_i_0, Q => \TMONOS\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    MONOUT : DFFB
      port map(CLK => CLK_c_c, D => N_30, CLR => HWRES_c_33, SET
         => nLBRDY_c_i_0, Q => \LEDint[5]\);
    
    MONOUT_0_i : OA21FTT
      port map(A => TICK_0(2), B => \TMONOS\, C => \LEDint[5]\, Y
         => N_30);
    
    TMONOS_i_0 : INV
      port map(A => nLBRDY_c, Y => nLBRDY_c_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity ctrl is

    port( TST_c_c      : in    std_logic_vector(3 to 3);
          PULSE        : in    std_logic_vector(2 to 2);
          TICK_0       : in    std_logic_vector(2 to 2);
          REG_15       : in    std_logic;
          REG_0        : in    std_logic;
          REG_1        : in    std_logic;
          REG_2        : in    std_logic;
          REG_3        : in    std_logic;
          REG_4        : in    std_logic;
          REG_5        : in    std_logic;
          TICK         : in    std_logic_vector(2 to 2);
          nLBRDY_c     : in    std_logic;
          EVNT_TRG     : in    std_logic;
          HWRES_c_32_0 : in    std_logic;
          RUN_c        : in    std_logic;
          HWRES_c_34   : in    std_logic;
          CLK_c_c      : in    std_logic;
          HWRES_c_33   : in    std_logic;
          N_18         : out   std_logic;
          N_20         : out   std_logic;
          N_22         : out   std_logic;
          N_24         : out   std_logic;
          N_26         : out   std_logic;
          N_28         : out   std_logic
        );

end ctrl;

architecture DEF_ARCH of ctrl is 

  component MONOSTABLE_3
    port( LEDint     : out   std_logic_vector(2 to 2);
          TICK_0     : in    std_logic_vector(2 to 2) := (others => 'U');
          CLK_c_c    : in    std_logic := 'U';
          HWRES_c_33 : in    std_logic := 'U';
          TMONOS     : in    std_logic := 'U'
        );
  end component;

  component OA21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MONOSTABLE_2
    port( TICK_0     : in    std_logic_vector(2 to 2) := (others => 'U');
          CLK_c_c    : in    std_logic := 'U';
          HWRES_c_33 : in    std_logic := 'U';
          TMONOS     : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MONOSTABLE_1
    port( LEDint       : out   std_logic_vector(1 to 1);
          TICK_0       : in    std_logic_vector(2 to 2) := (others => 'U');
          PULSE        : in    std_logic_vector(2 to 2) := (others => 'U');
          HWRES_c_33   : in    std_logic := 'U';
          CLK_c_c      : in    std_logic := 'U';
          HWRES_c_32_0 : in    std_logic := 'U';
          EVNT_TRG     : in    std_logic := 'U'
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MONOSTABLE
    port( LEDint       : out   std_logic_vector(0 to 0);
          TICK_0       : in    std_logic_vector(2 to 2) := (others => 'U');
          CLK_c_c      : in    std_logic := 'U';
          RUN_c        : in    std_logic := 'U';
          HWRES_c_32_0 : in    std_logic := 'U'
        );
  end component;

  component MONOSTABLE_4
    port( LEDint     : out   std_logic_vector(4 to 4);
          TICK_0     : in    std_logic_vector(2 to 2) := (others => 'U');
          TST_c_c    : in    std_logic_vector(3 to 3) := (others => 'U');
          CLK_c_c    : in    std_logic := 'U';
          HWRES_c_33 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component MONOSTABLE_5
    port( LEDint     : out   std_logic_vector(5 to 5);
          TICK_0     : in    std_logic_vector(2 to 2) := (others => 'U');
          CLK_c_c    : in    std_logic := 'U';
          HWRES_c_33 : in    std_logic := 'U';
          nLBRDY_c   : in    std_logic := 'U'
        );
  end component;

    signal \LEDForce\, \LEDint[5]\, N_165, \LEDbus[5]_net_1\, 
        \LEDint[4]\, N_163, \LEDbus[4]_net_1\, \LEDbus[3]_net_1\, 
        N_160, \LEDbus[2]_net_1\, \LEDint[2]\, \LEDint[1]\, N_158, 
        \LEDbus[1]_net_1\, \LEDint[0]\, N_156, \LEDbus[0]_net_1\, 
        \LEDbus_23\, N_155, \tmonos\, \LEDbus_22\, N_154, 
        \LEDbus_21\, N_153, \LEDbus_20\, N_152, \LEDbus_19\, 
        N_151, \LEDbus_18\, N_150, \LEDForce_17\, N_149, 
        \tmonos_16_0_a2\, \TMONOS\, \GND\, \VCC\ : std_logic;

    for all : MONOSTABLE_3
	Use entity work.MONOSTABLE_3(DEF_ARCH);
    for all : MONOSTABLE_2
	Use entity work.MONOSTABLE_2(DEF_ARCH);
    for all : MONOSTABLE_1
	Use entity work.MONOSTABLE_1(DEF_ARCH);
    for all : MONOSTABLE
	Use entity work.MONOSTABLE(DEF_ARCH);
    for all : MONOSTABLE_4
	Use entity work.MONOSTABLE_4(DEF_ARCH);
    for all : MONOSTABLE_5
	Use entity work.MONOSTABLE_5(DEF_ARCH);
begin 


    LED3_DRV : MONOSTABLE_3
      port map(LEDint(2) => \LEDint[2]\, TICK_0(2) => TICK_0(2), 
        CLK_c_c => CLK_c_c, HWRES_c_33 => HWRES_c_33, TMONOS => 
        \TMONOS\);
    
    \LED_i[5]\ : OA21TTF
      port map(A => \LEDForce\, B => \LEDint[5]\, C => N_165, Y
         => N_28);
    
    LEDForce_2_i_a2 : OR2
      port map(A => \tmonos\, B => REG_15, Y => N_149);
    
    \LEDbus_3_i_a2[3]\ : OR2
      port map(A => \tmonos\, B => REG_3, Y => N_153);
    
    \LED_i[2]\ : OA21FTT
      port map(A => \LEDForce\, B => \LEDbus[2]_net_1\, C => 
        N_160, Y => N_22);
    
    \LEDbus[3]\ : DFFS
      port map(CLK => CLK_c_c, D => \LEDbus_21\, SET => 
        HWRES_c_33, Q => \LEDbus[3]_net_1\);
    
    LED2_DRV : MONOSTABLE_2
      port map(TICK_0(2) => TICK_0(2), CLK_c_c => CLK_c_c, 
        HWRES_c_33 => HWRES_c_33, TMONOS => \TMONOS\);
    
    tmonos : DFFS
      port map(CLK => CLK_c_c, D => \tmonos_16_0_a2\, SET => 
        HWRES_c_34, Q => \tmonos\);
    
    LEDbus_19 : MUX2H
      port map(A => \LEDbus[1]_net_1\, B => N_151, S => TICK(2), 
        Y => \LEDbus_19\);
    
    LEDForce : DFFS
      port map(CLK => CLK_c_c, D => \LEDForce_17\, SET => 
        HWRES_c_33, Q => \LEDForce\);
    
    LEDbus_23 : MUX2H
      port map(A => \LEDbus[5]_net_1\, B => N_155, S => TICK(2), 
        Y => \LEDbus_23\);
    
    \LEDbus[5]\ : DFFS
      port map(CLK => CLK_c_c, D => \LEDbus_23\, SET => 
        HWRES_c_34, Q => \LEDbus[5]_net_1\);
    
    LED1_DRV : MONOSTABLE_1
      port map(LEDint(1) => \LEDint[1]\, TICK_0(2) => TICK_0(2), 
        PULSE(2) => PULSE(2), HWRES_c_33 => HWRES_c_33, CLK_c_c
         => CLK_c_c, HWRES_c_32_0 => HWRES_c_32_0, EVNT_TRG => 
        EVNT_TRG);
    
    \LED_i_a2[4]\ : NOR2FT
      port map(A => \LEDForce\, B => \LEDbus[4]_net_1\, Y => 
        N_163);
    
    \LEDbus[1]\ : DFFS
      port map(CLK => CLK_c_c, D => \LEDbus_19\, SET => 
        HWRES_c_33, Q => \LEDbus[1]_net_1\);
    
    \LED_i[3]\ : OA21FTT
      port map(A => \LEDForce\, B => \LEDbus[3]_net_1\, C => 
        N_160, Y => N_24);
    
    \LED_i_a2[2]\ : OR2
      port map(A => \LEDForce\, B => \LEDint[2]\, Y => N_160);
    
    \LEDbus_3_i_a2[0]\ : OR2
      port map(A => \tmonos\, B => REG_0, Y => N_150);
    
    LED0_DRV : MONOSTABLE
      port map(LEDint(0) => \LEDint[0]\, TICK_0(2) => TICK_0(2), 
        CLK_c_c => CLK_c_c, RUN_c => RUN_c, HWRES_c_32_0 => 
        HWRES_c_32_0);
    
    LED4_DRV : MONOSTABLE_4
      port map(LEDint(4) => \LEDint[4]\, TICK_0(2) => TICK_0(2), 
        TST_c_c(3) => TST_c_c(3), CLK_c_c => CLK_c_c, HWRES_c_33
         => HWRES_c_33);
    
    \LEDbus[4]\ : DFFS
      port map(CLK => CLK_c_c, D => \LEDbus_22\, SET => 
        HWRES_c_34, Q => \LEDbus[4]_net_1\);
    
    \LEDbus[2]\ : DFFS
      port map(CLK => CLK_c_c, D => \LEDbus_20\, SET => 
        HWRES_c_33, Q => \LEDbus[2]_net_1\);
    
    LEDbus_22 : MUX2H
      port map(A => \LEDbus[4]_net_1\, B => N_154, S => TICK(2), 
        Y => \LEDbus_22\);
    
    \LED_i[1]\ : OA21TTF
      port map(A => \LEDForce\, B => \LEDint[1]\, C => N_158, Y
         => N_20);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \LED_i_a2[5]\ : NOR2FT
      port map(A => \LEDForce\, B => \LEDbus[5]_net_1\, Y => 
        N_165);
    
    LEDbus_20 : MUX2H
      port map(A => \LEDbus[2]_net_1\, B => N_152, S => TICK(2), 
        Y => \LEDbus_20\);
    
    LEDbus_18 : MUX2H
      port map(A => \LEDbus[0]_net_1\, B => N_150, S => TICK(2), 
        Y => \LEDbus_18\);
    
    \LED_i_a2[0]\ : NOR2FT
      port map(A => \LEDForce\, B => \LEDbus[0]_net_1\, Y => 
        N_156);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \LED_i[4]\ : OA21TTF
      port map(A => \LEDForce\, B => \LEDint[4]\, C => N_163, Y
         => N_26);
    
    LED5_DRV : MONOSTABLE_5
      port map(LEDint(5) => \LEDint[5]\, TICK_0(2) => TICK_0(2), 
        CLK_c_c => CLK_c_c, HWRES_c_33 => HWRES_c_33, nLBRDY_c
         => nLBRDY_c);
    
    \LEDbus_3_i_a2[2]\ : OR2
      port map(A => \tmonos\, B => REG_2, Y => N_152);
    
    tmonos_16_0_a2 : NOR2FT
      port map(A => \tmonos\, B => TICK_0(2), Y => 
        \tmonos_16_0_a2\);
    
    LEDbus_21 : MUX2H
      port map(A => \LEDbus[3]_net_1\, B => N_153, S => TICK(2), 
        Y => \LEDbus_21\);
    
    \LEDbus[0]\ : DFFS
      port map(CLK => CLK_c_c, D => \LEDbus_18\, SET => 
        HWRES_c_33, Q => \LEDbus[0]_net_1\);
    
    \LED_i_a2[1]\ : NOR2FT
      port map(A => \LEDForce\, B => \LEDbus[1]_net_1\, Y => 
        N_158);
    
    \LED_i[0]\ : OA21TTF
      port map(A => \LEDForce\, B => \LEDint[0]\, C => N_156, Y
         => N_18);
    
    \LEDbus_3_i_a2[5]\ : OR2
      port map(A => \tmonos\, B => REG_5, Y => N_155);
    
    \LEDbus_3_i_a2[4]\ : OR2
      port map(A => \tmonos\, B => REG_4, Y => N_154);
    
    \LEDbus_3_i_a2[1]\ : OR2
      port map(A => \tmonos\, B => REG_1, Y => N_151);
    
    LEDForce_17 : MUX2H
      port map(A => \LEDForce\, B => N_149, S => TICK(2), Y => 
        \LEDForce_17\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity DAC_INTERF is

    port( TICK_0        : in    std_logic_vector(2 to 2);
          SYNC_c        : out   std_logic_vector(15 downto 0);
          DACCFG_DT     : in    std_logic_vector(15 downto 0);
          REG           : in    std_logic_vector(264 downto 233);
          PULSE         : in    std_logic_vector(9 to 9);
          DACCFG_RAD    : out   std_logic_vector(3 downto 0);
          HWRES_c_36    : in    std_logic;
          HWRES_c_34    : in    std_logic;
          HWRES_c_35    : in    std_logic;
          RUN_c_0       : in    std_logic;
          DACCFG_nRD    : out   std_logic;
          SCLK_DAC_c    : out   std_logic;
          SDIN_DAC_c    : out   std_logic;
          HWRES_c_0     : in    std_logic;
          HWRES_c_3     : in    std_logic;
          HWRES_c_0_6_0 : in    std_logic;
          HWRES_c_2     : in    std_logic;
          HWRES_c_1     : in    std_logic;
          HWRES_c_36_0  : in    std_logic;
          CLK_c_c       : in    std_logic;
          HWRES_c       : in    std_logic
        );

end DAC_INTERF;

architecture DEF_ARCH of DAC_INTERF is 

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component AO21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \sstate_1[6]_net_1\, \sstate_ns[0]_net_1\, 
        \sstate_0[6]_net_1\, \sstate_2[0]_net_1\, 
        \sstate[1]_net_1\, \sstate_1[0]_net_1\, 
        \sstate_0[0]_net_1\, \sstate_0[5]_net_1\, N_191_i_0, 
        \un1_sstate_16_0\, N_207, sstate_0_sqmuxa_0, N_364, 
        \DWACT_ADD_CI_0_g_array_1[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \BITCNT[1]_net_1\, \DWACT_ADD_CI_0_g_array_12[0]\, 
        \BITCNT[2]_net_1\, \DWACT_ADD_CI_0_g_array_1_0[0]\, 
        \DWACT_ADD_CI_0_TMP_0[0]\, 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, \sstate_ns_i_1_i[1]\, 
        \sstate_ns_i_a3[1]_net_1\, ISI_0_sqmuxa, N_191_1, 
        \sstate[4]_net_1\, N_225_1, un1_hwres_16_i, un1_reg_9_i, 
        un1_hwres_3_i, un1_reg_3_i, un1_hwres_7_i, un1_reg_2_i, 
        un1_hwres_15_i, un1_reg_5_i, un1_hwres_9_i, un1_reg_11_i, 
        un1_hwres_1_i, un1_reg_6_i, un1_hwres_8_i, un1_reg_7_i, 
        un1_hwres_14_i, un1_reg_10_i, un1_hwres_11_i, 
        un1_reg_12_i, un1_hwres_13_i, un1_reg_8_i, un1_hwres_6_i, 
        un1_reg_13_i, un1_hwres_10_i, un1_reg_14_i, 
        un1_hwres_12_i, un1_reg_1_i, un1_hwres_2_i, un1_reg_15_i, 
        un1_hwres_4_i, un1_reg_4_i, un1_hwres_5_i, un1_reg_16_i, 
        \un1_sstate_5_i_a2\, \un1_sstate_17_i_a3\, N_208, 
        \sstate[3]_net_1\, \sstate_ns[4]_net_1\, \un6_bitcnt\, 
        sstate_0_sqmuxa, N_220, \LastDac\, \RefreshCycle\, 
        \LastDac_21\, \sstate_i_0[6]\, \un1_sstate_20\, 
        \sstate[2]_net_1\, LastDac_1_sqmuxa_i, \un15_sync[15]\, 
        \ISI_20\, ISI_6, N_201, \ISI_6_iv_0\, \SWORD[15]_net_1\, 
        \DACCFG_DT_m[15]_net_1\, \SWORD_19\, \SWORD_6[15]_net_1\, 
        N_314, \SWORD[14]_net_1\, \SWORD_18\, \SWORD_6[14]_net_1\, 
        N_363, \SWORD[13]_net_1\, \SWORD_17\, \SWORD_6[13]_net_1\, 
        N_362, \SWORD[12]_net_1\, \SWORD_16\, \SWORD_6[12]_net_1\, 
        N_361, \SWORD[11]_net_1\, \SWORD_15\, \SWORD_6[11]_net_1\, 
        N_360, \SWORD[10]_net_1\, \SWORD_14\, \SWORD_6[10]_net_1\, 
        N_359, \SWORD[9]_net_1\, \SWORD_13\, \SWORD_6[9]_net_1\, 
        N_358, \SWORD[8]_net_1\, \SWORD_12\, \SWORD_6[8]_net_1\, 
        N_357, \SWORD[7]_net_1\, \sstate[5]_net_1\, \SWORD_11\, 
        \SWORD_6[7]_net_1\, un1_sstate_16, N_356, 
        \SWORD[6]_net_1\, \SWORD_10\, \SWORD_6[6]_net_1\, N_355, 
        \SWORD[5]_net_1\, \SWORD_9\, \SWORD_6[5]_net_1\, N_354, 
        \SWORD[4]_net_1\, \SWORD_8\, \SWORD_6[4]_net_1\, N_353, 
        \SWORD[3]_net_1\, \SWORD_7\, \SWORD_6[3]_net_1\, N_352, 
        \SWORD[2]_net_1\, \SWORD_6\, \SWORD_6[2]_net_1\, N_351, 
        \SWORD[1]_net_1\, \SWORD_5\, \SWORD_6[1]_net_1\, N_350, 
        \SWORD[0]_net_1\, \SWORD_4\, \SWORD_6[0]_net_1\, N_349, 
        \RefreshCycle_3\, N_364_i_0, \ISCK_2\, N_199, 
        \DACCFG_nRD_1\, \sstate_i_0[2]\, N_218, \BITCNT_5[3]\, 
        I_17, \BITCNT_5[2]\, I_18, \BITCNT_5[1]\, I_15, 
        \BITCNT_5[0]\, \DWACT_ADD_CI_0_partial_sum[0]\, 
        \ISI_0_sqmuxa_0_a2_2\, \BITCNT[3]_net_1\, 
        \BITCNT[0]_net_1\, \DACRdPnt_2[3]_net_1\, I_17_0, 
        \DACRdPnt_2[2]_net_1\, I_18_0, \DACRdPnt_2[1]_net_1\, 
        I_15_0, \DACRdPnt_2[0]_net_1\, 
        \DWACT_ADD_CI_0_partial_sum_0[0]\, \SYNC_5[15]_net_1\, 
        N_296, N_278, \un15_sync_1[15]\, \un15_sync_2[15]\, 
        \SYNC_5[14]_net_1\, N_295, N_277, \un15_sync[14]\, 
        \un15_sync_1[14]\, \SYNC_5[13]_net_1\, N_294, N_276, 
        \un15_sync[13]\, \un15_sync_1[13]\, \SYNC_5[12]_net_1\, 
        N_293, N_275, \un15_sync[12]\, \un15_sync_1[12]\, 
        \DACCFG_RAD[2]\, \SYNC_5[11]_net_1\, N_292, N_274, 
        \un15_sync[11]\, \un15_sync_1[11]\, \SYNC_5[10]_net_1\, 
        N_291, N_273, \un15_sync[10]\, \SYNC_5[9]_net_1\, N_290, 
        N_272, \un15_sync[9]\, \SYNC_5[8]_net_1\, N_289, N_271, 
        \un15_sync[8]\, \DACCFG_RAD[3]\, \SYNC_5[7]_net_1\, N_288, 
        N_270, \un15_sync[7]\, \sstate[6]_net_1\, 
        \un15_sync_1[7]\, \SYNC_5[6]_net_1\, N_287, N_269, 
        \un15_sync[6]\, \sstate[0]_net_1\, \SYNC_5[5]_net_1\, 
        N_286, N_268, \un15_sync[5]\, \SYNC_5[4]_net_1\, N_285, 
        N_267, \un15_sync[4]\, \SYNC_5[3]_net_1\, N_284, N_266, 
        \un15_sync[3]\, \un15_sync_1[3]\, \DACCFG_RAD[1]\, 
        \SYNC_5[2]_net_1\, N_283, N_265, \un15_sync[2]\, 
        \DACCFG_RAD[0]\, \SYNC_5[1]_net_1\, N_282, N_264, 
        \un15_sync[1]\, \SYNC_5[0]_net_1\, N_281, N_263, 
        \un15_sync[0]\, \SYNC_c[0]\, \SYNC_c[1]\, \SYNC_c[2]\, 
        \SYNC_c[3]\, \SYNC_c[4]\, \SYNC_c[5]\, \SYNC_c[6]\, 
        \SYNC_c[7]\, \SYNC_c[8]\, \SYNC_c[9]\, \SYNC_c[10]\, 
        \SYNC_c[11]\, \SYNC_c[12]\, \SYNC_c[13]\, \SYNC_c[14]\, 
        \SYNC_c[15]\, \SDIN_DAC_c\, \SCLK_DAC_c\, 
        DACCFG_nRD_net_1, \GND\, \VCC\ : std_logic;

begin 

    SYNC_c(15) <= \SYNC_c[15]\;
    SYNC_c(14) <= \SYNC_c[14]\;
    SYNC_c(13) <= \SYNC_c[13]\;
    SYNC_c(12) <= \SYNC_c[12]\;
    SYNC_c(11) <= \SYNC_c[11]\;
    SYNC_c(10) <= \SYNC_c[10]\;
    SYNC_c(9) <= \SYNC_c[9]\;
    SYNC_c(8) <= \SYNC_c[8]\;
    SYNC_c(7) <= \SYNC_c[7]\;
    SYNC_c(6) <= \SYNC_c[6]\;
    SYNC_c(5) <= \SYNC_c[5]\;
    SYNC_c(4) <= \SYNC_c[4]\;
    SYNC_c(3) <= \SYNC_c[3]\;
    SYNC_c(2) <= \SYNC_c[2]\;
    SYNC_c(1) <= \SYNC_c[1]\;
    SYNC_c(0) <= \SYNC_c[0]\;
    DACCFG_RAD(3) <= \DACCFG_RAD[3]\;
    DACCFG_RAD(2) <= \DACCFG_RAD[2]\;
    DACCFG_RAD(1) <= \DACCFG_RAD[1]\;
    DACCFG_RAD(0) <= \DACCFG_RAD[0]\;
    DACCFG_nRD <= DACCFG_nRD_net_1;
    SCLK_DAC_c <= \SCLK_DAC_c\;
    SDIN_DAC_c <= \SDIN_DAC_c\;

    un1_hwres_11 : NOR2FT
      port map(A => HWRES_c_1, B => REG(238), Y => un1_hwres_11_i);
    
    \SWORD_6_0[11]\ : MUX2H
      port map(A => REG(260), B => DACCFG_DT(11), S => 
        \sstate_0[0]_net_1\, Y => N_360);
    
    \SYNC_5_0[5]\ : MUX2H
      port map(A => \SYNC_c[5]\, B => REG(238), S => 
        \sstate[6]_net_1\, Y => N_268);
    
    \SWORD_6_0[7]\ : MUX2H
      port map(A => REG(256), B => DACCFG_DT(7), S => 
        \sstate_1[0]_net_1\, Y => N_356);
    
    \BITCNT[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_5[0]\, CLR => 
        HWRES_c_34, Q => \BITCNT[0]_net_1\);
    
    \SWORD_6[5]\ : MUX2H
      port map(A => N_354, B => \SWORD[4]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[5]_net_1\);
    
    SWORD_15 : MUX2H
      port map(A => \SWORD[11]_net_1\, B => \SWORD_6[11]_net_1\, 
        S => \un1_sstate_16_0\, Y => \SWORD_15\);
    
    un15_sync_14 : NAND2
      port map(A => \un15_sync_1[14]\, B => \un15_sync_2[15]\, Y
         => \un15_sync[14]\);
    
    \DACRdPnt[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACRdPnt_2[3]_net_1\, CLR
         => HWRES_c_34, Q => \DACCFG_RAD[3]\);
    
    un1_BITCNT_I_19 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \BITCNT[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \SWORD_6[7]\ : MUX2H
      port map(A => N_356, B => \SWORD[6]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[7]_net_1\);
    
    \SYNC_5_s[5]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_286, Y => 
        \SYNC_5[5]_net_1\);
    
    \sstate_ns_i_1[1]\ : NOR2
      port map(A => \sstate[1]_net_1\, B => \sstate[2]_net_1\, Y
         => N_191_1);
    
    \SYNC_5[12]\ : MUX2H
      port map(A => N_275, B => \un15_sync[12]\, S => 
        \sstate_2[0]_net_1\, Y => N_293);
    
    \SWORD_6[9]\ : MUX2H
      port map(A => N_358, B => \SWORD[8]_net_1\, S => 
        \sstate_0[5]_net_1\, Y => \SWORD_6[9]_net_1\);
    
    ISCK_2 : MUX2H
      port map(A => \sstate[5]_net_1\, B => \SCLK_DAC_c\, S => 
        N_199, Y => \ISCK_2\);
    
    \SYNC_1[4]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[4]_net_1\, CLR => 
        un1_hwres_14_i, SET => un1_reg_10_i, Q => \SYNC_c[4]\);
    
    ISCK : DFFC
      port map(CLK => CLK_c_c, D => \ISCK_2\, CLR => HWRES_c_35, 
        Q => \SCLK_DAC_c\);
    
    \SWORD[14]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_18\, CLR => HWRES_c_35, 
        Q => \SWORD[14]_net_1\);
    
    \SYNC_1[0]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[0]_net_1\, CLR => 
        un1_hwres_8_i, SET => un1_reg_7_i, Q => \SYNC_c[0]\);
    
    \sstate_i[2]\ : INV
      port map(A => \sstate[2]_net_1\, Y => \sstate_i_0[2]\);
    
    \SYNC_1[12]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[12]_net_1\, CLR => 
        un1_hwres_9_i, SET => un1_reg_11_i, Q => \SYNC_c[12]\);
    
    un15_sync_5 : NAND2
      port map(A => \un15_sync_1[7]\, B => \un15_sync_1[13]\, Y
         => \un15_sync[5]\);
    
    \DACCFG_nRD\ : DFFS
      port map(CLK => CLK_c_c, D => \DACCFG_nRD_1\, SET => 
        HWRES_c_34, Q => DACCFG_nRD_net_1);
    
    un15_sync_1 : NAND2
      port map(A => \un15_sync_1[3]\, B => \un15_sync_1[13]\, Y
         => \un15_sync[1]\);
    
    \SWORD_6[4]\ : MUX2H
      port map(A => N_353, B => \SWORD[3]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[4]_net_1\);
    
    un15_sync_7_1 : NOR2FT
      port map(A => \DACCFG_RAD[2]\, B => \DACCFG_RAD[3]\, Y => 
        \un15_sync_1[7]\);
    
    \SYNC_5[13]\ : MUX2H
      port map(A => N_276, B => \un15_sync[13]\, S => 
        \sstate_2[0]_net_1\, Y => N_294);
    
    \SYNC_5_0[11]\ : MUX2H
      port map(A => \SYNC_c[11]\, B => REG(244), S => 
        \sstate_1[6]_net_1\, Y => N_274);
    
    \SYNC_5[10]\ : MUX2H
      port map(A => N_273, B => \un15_sync[10]\, S => 
        \sstate_2[0]_net_1\, Y => N_291);
    
    \SWORD[9]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_13\, CLR => 
        HWRES_c_36_0, Q => \SWORD[9]_net_1\);
    
    LastDac_21_i : INV
      port map(A => \sstate_1[6]_net_1\, Y => \sstate_i_0[6]\);
    
    \SYNC_5[15]\ : MUX2H
      port map(A => N_278, B => \un15_sync[15]\, S => 
        \sstate_2[0]_net_1\, Y => N_296);
    
    \SWORD_6[2]\ : MUX2H
      port map(A => N_351, B => \SWORD[1]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[2]_net_1\);
    
    \SWORD_6_0[1]\ : MUX2H
      port map(A => REG(250), B => DACCFG_DT(1), S => 
        \sstate_1[0]_net_1\, Y => N_350);
    
    SWORD_9 : MUX2H
      port map(A => \SWORD[5]_net_1\, B => \SWORD_6[5]_net_1\, S
         => un1_sstate_16, Y => \SWORD_9\);
    
    \SWORD[6]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_10\, CLR => HWRES_c_36, 
        Q => \SWORD[6]_net_1\);
    
    \DACRdPnt_2[1]\ : NOR2FT
      port map(A => I_15_0, B => \sstate_0[6]_net_1\, Y => 
        \DACRdPnt_2[1]_net_1\);
    
    \SYNC_1[13]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[13]_net_1\, CLR => 
        un1_hwres_3_i, SET => un1_reg_3_i, Q => \SYNC_c[13]\);
    
    un1_hwres_6 : NOR2FT
      port map(A => HWRES_c_0_6_0, B => REG(242), Y => 
        un1_hwres_6_i);
    
    un15_sync_15_2 : AND2
      port map(A => \DACCFG_RAD[2]\, B => \DACCFG_RAD[3]\, Y => 
        \un15_sync_2[15]\);
    
    \SYNC_1[10]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[10]_net_1\, CLR => 
        un1_hwres_10_i, SET => un1_reg_14_i, Q => \SYNC_c[10]\);
    
    \SYNC_1[15]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[15]_net_1\, CLR => 
        un1_hwres_4_i, SET => un1_reg_4_i, Q => \SYNC_c[15]\);
    
    SWORD_6 : MUX2H
      port map(A => \SWORD[2]_net_1\, B => \SWORD_6[2]_net_1\, S
         => un1_sstate_16, Y => \SWORD_6\);
    
    \SWORD_6_0[2]\ : MUX2H
      port map(A => REG(251), B => DACCFG_DT(2), S => 
        \sstate_1[0]_net_1\, Y => N_351);
    
    un15_sync_9 : NAND2
      port map(A => \un15_sync_1[11]\, B => \un15_sync_1[13]\, Y
         => \un15_sync[9]\);
    
    \SYNC_5_s[6]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_287, Y => 
        \SYNC_5[6]_net_1\);
    
    \SWORD[8]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_12\, CLR => HWRES_c_36, 
        Q => \SWORD[8]_net_1\);
    
    \SYNC_1[6]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[6]_net_1\, CLR => 
        un1_hwres_15_i, SET => un1_reg_5_i, Q => \SYNC_c[6]\);
    
    SWORD_19 : MUX2H
      port map(A => \SWORD[15]_net_1\, B => \SWORD_6[15]_net_1\, 
        S => \un1_sstate_16_0\, Y => \SWORD_19\);
    
    \DACRdPnt_2[0]\ : NOR2FT
      port map(A => \DWACT_ADD_CI_0_partial_sum_0[0]\, B => 
        \sstate_0[6]_net_1\, Y => \DACRdPnt_2[0]_net_1\);
    
    un1_DACRdPnt_I_17 : XOR2
      port map(A => \DACCFG_RAD[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12_0[0]\, Y => I_17_0);
    
    \sstate_1[6]\ : DFFS
      port map(CLK => CLK_c_c, D => \sstate_ns[0]_net_1\, SET => 
        HWRES_c, Q => \sstate_1[6]_net_1\);
    
    \SYNC_5_s[15]\ : OR2FT
      port map(A => sstate_0_sqmuxa, B => N_296, Y => 
        \SYNC_5[15]_net_1\);
    
    \SYNC_5_s[7]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_288, Y => 
        \SYNC_5[7]_net_1\);
    
    SWORD_8 : MUX2H
      port map(A => \SWORD[4]_net_1\, B => \SWORD_6[4]_net_1\, S
         => un1_sstate_16, Y => \SWORD_8\);
    
    \SWORD[10]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_14\, CLR => HWRES_c_35, 
        Q => \SWORD[10]_net_1\);
    
    RefreshCycle_3_i : INV
      port map(A => N_364, Y => N_364_i_0);
    
    un15_sync_6 : NAND2
      port map(A => \un15_sync_1[7]\, B => \un15_sync_1[14]\, Y
         => \un15_sync[6]\);
    
    \sstate_1[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[1]_net_1\, CLR => 
        HWRES_c_36_0, Q => \sstate_1[0]_net_1\);
    
    un4_g_sim_on : NAND2
      port map(A => RUN_c_0, B => TICK_0(2), Y => N_364);
    
    un1_sstate_19_i : OAI21
      port map(A => \un1_sstate_5_i_a2\, B => \sstate[3]_net_1\, 
        C => ISI_0_sqmuxa, Y => N_201);
    
    \SWORD_6_0[12]\ : MUX2H
      port map(A => REG(261), B => DACCFG_DT(12), S => 
        \sstate_0[0]_net_1\, Y => N_361);
    
    \SWORD_6_0[6]\ : MUX2H
      port map(A => REG(255), B => DACCFG_DT(6), S => 
        \sstate_1[0]_net_1\, Y => N_355);
    
    un1_reg_4 : AND2
      port map(A => HWRES_c_3, B => REG(248), Y => un1_reg_4_i);
    
    \SYNC_5[7]\ : MUX2H
      port map(A => N_270, B => \un15_sync[7]\, S => 
        \sstate_2[0]_net_1\, Y => N_288);
    
    \SYNC_5_0[13]\ : MUX2H
      port map(A => \SYNC_c[13]\, B => REG(246), S => 
        \sstate_1[6]_net_1\, Y => N_276);
    
    sstate_0_sqmuxa_0_a3 : OR2FT
      port map(A => \sstate_0[6]_net_1\, B => N_364, Y => 
        sstate_0_sqmuxa);
    
    un1_sstate_8_0_a3 : NOR3
      port map(A => \sstate[5]_net_1\, B => \sstate[3]_net_1\, C
         => \sstate[4]_net_1\, Y => N_218);
    
    \SYNC_5_0[3]\ : MUX2H
      port map(A => \SYNC_c[3]\, B => REG(236), S => 
        \sstate[6]_net_1\, Y => N_266);
    
    un15_sync_12_1 : NOR2
      port map(A => \DACCFG_RAD[0]\, B => \DACCFG_RAD[1]\, Y => 
        \un15_sync_1[12]\);
    
    un15_sync_11_1 : NOR2FT
      port map(A => \DACCFG_RAD[3]\, B => \DACCFG_RAD[2]\, Y => 
        \un15_sync_1[11]\);
    
    un1_hwres_5 : NOR2FT
      port map(A => HWRES_c_0, B => REG(236), Y => un1_hwres_5_i);
    
    un1_reg_5 : AND2
      port map(A => HWRES_c_2, B => REG(239), Y => un1_reg_5_i);
    
    \SYNC_5_0[1]\ : MUX2H
      port map(A => \SYNC_c[1]\, B => REG(234), S => 
        \sstate[6]_net_1\, Y => N_264);
    
    un1_reg_1 : AND2
      port map(A => HWRES_c_3, B => REG(235), Y => un1_reg_1_i);
    
    \SWORD[12]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_16\, CLR => HWRES_c_35, 
        Q => \SWORD[12]_net_1\);
    
    ISI_6_iv : AO21TTF
      port map(A => N_208, B => REG(264), C => \ISI_6_iv_0\, Y
         => ISI_6);
    
    un1_sstate_7_i : OR2FT
      port map(A => N_191_1, B => \sstate_0[0]_net_1\, Y => N_199);
    
    un1_BITCNT_I_1 : AND2
      port map(A => \BITCNT[0]_net_1\, B => \un1_sstate_17_i_a3\, 
        Y => \DWACT_ADD_CI_0_TMP[0]\);
    
    \SYNC_5_s[0]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_281, Y => 
        \SYNC_5[0]_net_1\);
    
    un1_DACRdPnt_I_15 : XOR2
      port map(A => \DACCFG_RAD[1]\, B => 
        \DWACT_ADD_CI_0_TMP_0[0]\, Y => I_15_0);
    
    \SWORD[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_8\, CLR => HWRES_c_36, 
        Q => \SWORD[4]_net_1\);
    
    un1_hwres_15 : NOR2FT
      port map(A => HWRES_c_1, B => REG(239), Y => un1_hwres_15_i);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SYNC_5_s[2]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_283, Y => 
        \SYNC_5[2]_net_1\);
    
    \SWORD_6_0[0]\ : MUX2H
      port map(A => REG(249), B => DACCFG_DT(0), S => 
        \sstate_1[0]_net_1\, Y => N_349);
    
    \SYNC_5_s[1]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_282, Y => 
        \SYNC_5[1]_net_1\);
    
    SWORD_4 : MUX2H
      port map(A => \SWORD[0]_net_1\, B => \SWORD_6[0]_net_1\, S
         => un1_sstate_16, Y => \SWORD_4\);
    
    ISI_0_sqmuxa_0_a2 : NAND3
      port map(A => \ISI_0_sqmuxa_0_a2_2\, B => \BITCNT[2]_net_1\, 
        C => \BITCNT[3]_net_1\, Y => ISI_0_sqmuxa);
    
    \SWORD_6_0[14]\ : MUX2H
      port map(A => REG(263), B => DACCFG_DT(14), S => 
        \sstate_0[0]_net_1\, Y => N_363);
    
    \SWORD[15]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_19\, CLR => HWRES_c_35, 
        Q => \SWORD[15]_net_1\);
    
    un1_reg_15 : AND2
      port map(A => HWRES_c_3, B => REG(247), Y => un1_reg_15_i);
    
    \sstate_0[6]\ : DFFS
      port map(CLK => CLK_c_c, D => \sstate_ns[0]_net_1\, SET => 
        HWRES_c, Q => \sstate_0[6]_net_1\);
    
    un1_reg_13 : AND2
      port map(A => HWRES_c_2, B => REG(242), Y => un1_reg_13_i);
    
    SWORD_18 : MUX2H
      port map(A => \SWORD[14]_net_1\, B => \SWORD_6[14]_net_1\, 
        S => \un1_sstate_16_0\, Y => \SWORD_18\);
    
    \SYNC_5_s[10]\ : OR2FT
      port map(A => sstate_0_sqmuxa, B => N_291, Y => 
        \SYNC_5[10]_net_1\);
    
    \sstate_ns_a3[0]\ : OR3FFT
      port map(A => \sstate_0[6]_net_1\, B => N_364, C => 
        PULSE(9), Y => N_220);
    
    \BITCNT_5_r[0]\ : OA21FTT
      port map(A => ISI_0_sqmuxa, B => 
        \DWACT_ADD_CI_0_partial_sum[0]\, C => N_207, Y => 
        \BITCNT_5[0]\);
    
    \SWORD_6[13]\ : MUX2H
      port map(A => N_362, B => \SWORD[12]_net_1\, S => 
        \sstate_0[5]_net_1\, Y => \SWORD_6[13]_net_1\);
    
    \SYNC_5[14]\ : MUX2H
      port map(A => N_277, B => \un15_sync[14]\, S => 
        \sstate_2[0]_net_1\, Y => N_295);
    
    un1_DACRdPnt_I_11 : XOR2
      port map(A => \DACCFG_RAD[0]\, B => \un1_sstate_5_i_a2\, Y
         => \DWACT_ADD_CI_0_partial_sum_0[0]\);
    
    \SYNC_5_s[14]\ : OR2FT
      port map(A => sstate_0_sqmuxa, B => N_295, Y => 
        \SYNC_5[14]_net_1\);
    
    \BITCNT[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_5[1]\, CLR => 
        HWRES_c_34, Q => \BITCNT[1]_net_1\);
    
    un1_DACRdPnt_I_18 : XOR2
      port map(A => \DACCFG_RAD[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1_0[0]\, Y => I_18_0);
    
    \SWORD_6_0[5]\ : MUX2H
      port map(A => REG(254), B => DACCFG_DT(5), S => 
        \sstate_1[0]_net_1\, Y => N_354);
    
    \SWORD_6[3]\ : MUX2H
      port map(A => N_352, B => \SWORD[2]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[3]_net_1\);
    
    \SYNC_1[14]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[14]_net_1\, CLR => 
        un1_hwres_2_i, SET => un1_reg_15_i, Q => \SYNC_c[14]\);
    
    \BITCNT_5_r[3]\ : OA21FTT
      port map(A => ISI_0_sqmuxa, B => I_17, C => N_207, Y => 
        \BITCNT_5[3]\);
    
    \DACRdPnt_2[3]\ : NOR2FT
      port map(A => I_17_0, B => \sstate_0[6]_net_1\, Y => 
        \DACRdPnt_2[3]_net_1\);
    
    un15_sync_15_1 : AND2
      port map(A => \DACCFG_RAD[0]\, B => \DACCFG_RAD[1]\, Y => 
        \un15_sync_1[15]\);
    
    \sstate[4]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[5]_net_1\, CLR => 
        HWRES_c, Q => \sstate[4]_net_1\);
    
    \DACCFG_DT_m[15]\ : NAND2
      port map(A => DACCFG_DT(15), B => \sstate_0[0]_net_1\, Y
         => \DACCFG_DT_m[15]_net_1\);
    
    \SWORD_6[0]\ : NOR2FT
      port map(A => N_349, B => \sstate_0[5]_net_1\, Y => 
        \SWORD_6[0]_net_1\);
    
    \sstate_ns[0]\ : OAI21FTT
      port map(A => \un6_bitcnt\, B => ISI_0_sqmuxa, C => N_220, 
        Y => \sstate_ns[0]_net_1\);
    
    \sstate_0[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[1]_net_1\, CLR => 
        HWRES_c_36_0, Q => \sstate_0[0]_net_1\);
    
    \SYNC_5[5]\ : MUX2H
      port map(A => N_268, B => \un15_sync[5]\, S => 
        \sstate[0]_net_1\, Y => N_286);
    
    \SWORD_6[10]\ : MUX2H
      port map(A => N_359, B => \SWORD[9]_net_1\, S => 
        \sstate_0[5]_net_1\, Y => \SWORD_6[10]_net_1\);
    
    un15_sync_11 : NAND2
      port map(A => \un15_sync_1[11]\, B => \un15_sync_1[15]\, Y
         => \un15_sync[11]\);
    
    \BITCNT_5_r[1]\ : OA21FTT
      port map(A => ISI_0_sqmuxa, B => I_15, C => N_207, Y => 
        \BITCNT_5[1]\);
    
    un1_reg_3 : AND2
      port map(A => HWRES_c_2, B => REG(246), Y => un1_reg_3_i);
    
    un1_sstate_5_i_a2 : OR2
      port map(A => \sstate_0[0]_net_1\, B => \sstate_0[6]_net_1\, 
        Y => \un1_sstate_5_i_a2\);
    
    un1_sstate_20 : OAI21TTF
      port map(A => \sstate[2]_net_1\, B => \sstate_0[6]_net_1\, 
        C => LastDac_1_sqmuxa_i, Y => \un1_sstate_20\);
    
    \SWORD_6_0[10]\ : MUX2H
      port map(A => REG(259), B => DACCFG_DT(10), S => 
        \sstate_0[0]_net_1\, Y => N_359);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    LastDac_21 : MUX2H
      port map(A => \sstate_i_0[6]\, B => \LastDac\, S => 
        \un1_sstate_20\, Y => \LastDac_21\);
    
    un1_DACRdPnt_I_1 : AND2
      port map(A => \DACCFG_RAD[0]\, B => \un1_sstate_5_i_a2\, Y
         => \DWACT_ADD_CI_0_TMP_0[0]\);
    
    \sstate_ns_i_a3[1]\ : AO21
      port map(A => N_364, B => PULSE(9), C => N_225_1, Y => 
        \sstate_ns_i_a3[1]_net_1\);
    
    \sstate[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[4]_net_1\, CLR => 
        HWRES_c_36_0, Q => \sstate[3]_net_1\);
    
    \BITCNT_5_r[2]\ : OA21FTT
      port map(A => ISI_0_sqmuxa, B => I_18, C => N_207, Y => 
        \BITCNT_5[2]\);
    
    \sstate[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[1]_net_1\, CLR => 
        HWRES_c_36_0, Q => \sstate[0]_net_1\);
    
    \SYNC_1[7]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[7]_net_1\, CLR => 
        un1_hwres_7_i, SET => un1_reg_2_i, Q => \SYNC_c[7]\);
    
    \SYNC_5[9]\ : MUX2H
      port map(A => N_272, B => \un15_sync[9]\, S => 
        \sstate_2[0]_net_1\, Y => N_290);
    
    \SYNC_1[9]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[9]_net_1\, CLR => 
        un1_hwres_6_i, SET => un1_reg_13_i, Q => \SYNC_c[9]\);
    
    un1_reg_12 : AND2
      port map(A => HWRES_c_2, B => REG(238), Y => un1_reg_12_i);
    
    un1_hwres_7 : NOR2FT
      port map(A => HWRES_c_1, B => REG(240), Y => un1_hwres_7_i);
    
    un1_hwres_9 : NOR2FT
      port map(A => HWRES_c_1, B => REG(245), Y => un1_hwres_9_i);
    
    \SWORD_6[6]\ : MUX2H
      port map(A => N_355, B => \SWORD[5]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[6]_net_1\);
    
    un1_DACRdPnt_I_19 : AND2
      port map(A => \DWACT_ADD_CI_0_TMP_0[0]\, B => 
        \DACCFG_RAD[1]\, Y => \DWACT_ADD_CI_0_g_array_1_0[0]\);
    
    \SWORD[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_7\, CLR => HWRES_c_36, 
        Q => \SWORD[3]_net_1\);
    
    \SYNC_5[8]\ : MUX2H
      port map(A => N_271, B => \un15_sync[8]\, S => 
        \sstate_2[0]_net_1\, Y => N_289);
    
    \SYNC_5_0[9]\ : MUX2H
      port map(A => \SYNC_c[9]\, B => REG(242), S => 
        \sstate_1[6]_net_1\, Y => N_272);
    
    un15_sync_0 : NAND2
      port map(A => \un15_sync_1[3]\, B => \un15_sync_1[12]\, Y
         => \un15_sync[0]\);
    
    \SYNC_1[3]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[3]_net_1\, CLR => 
        un1_hwres_5_i, SET => un1_reg_16_i, Q => \SYNC_c[3]\);
    
    SWORD_12 : MUX2H
      port map(A => \SWORD[8]_net_1\, B => \SWORD_6[8]_net_1\, S
         => \un1_sstate_16_0\, Y => \SWORD_12\);
    
    un1_BITCNT_I_18 : XOR2
      port map(A => \BITCNT[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_18);
    
    SWORD_17 : MUX2H
      port map(A => \SWORD[13]_net_1\, B => \SWORD_6[13]_net_1\, 
        S => \un1_sstate_16_0\, Y => \SWORD_17\);
    
    un1_reg_11 : AND2
      port map(A => HWRES_c_2, B => REG(245), Y => un1_reg_11_i);
    
    un1_DACRdPnt_I_21 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1_0[0]\, B => 
        \DACCFG_RAD[2]\, Y => \DWACT_ADD_CI_0_g_array_12_0[0]\);
    
    un1_reg_16 : AND2
      port map(A => HWRES_c_3, B => REG(236), Y => un1_reg_16_i);
    
    \SWORD_6[14]\ : MUX2H
      port map(A => N_363, B => \SWORD[13]_net_1\, S => 
        \sstate_0[5]_net_1\, Y => \SWORD_6[14]_net_1\);
    
    \sstate[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[2]_net_1\, CLR => 
        HWRES_c_36_0, Q => \sstate[1]_net_1\);
    
    \DACRdPnt[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACRdPnt_2[1]_net_1\, CLR
         => HWRES_c_34, Q => \DACCFG_RAD[1]\);
    
    \SYNC_5[0]\ : MUX2H
      port map(A => N_263, B => \un15_sync[0]\, S => 
        \sstate[0]_net_1\, Y => N_281);
    
    \DACRdPnt[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACRdPnt_2[2]_net_1\, CLR
         => HWRES_c_34, Q => \DACCFG_RAD[2]\);
    
    \SYNC_5_0[15]\ : MUX2H
      port map(A => \SYNC_c[15]\, B => REG(248), S => 
        \sstate_1[6]_net_1\, Y => N_278);
    
    \sstate[6]\ : DFFS
      port map(CLK => CLK_c_c, D => \sstate_ns[0]_net_1\, SET => 
        HWRES_c, Q => \sstate[6]_net_1\);
    
    \SWORD[7]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_11\, CLR => HWRES_c_36, 
        Q => \SWORD[7]_net_1\);
    
    ISI_0_sqmuxa_0_a2_2 : AND3
      port map(A => \sstate[3]_net_1\, B => \BITCNT[0]_net_1\, C
         => \BITCNT[1]_net_1\, Y => \ISI_0_sqmuxa_0_a2_2\);
    
    un1_hwres_8 : NOR2FT
      port map(A => HWRES_c_1, B => REG(233), Y => un1_hwres_8_i);
    
    \SWORD_6_0[13]\ : MUX2H
      port map(A => REG(262), B => DACCFG_DT(13), S => 
        \sstate_0[0]_net_1\, Y => N_362);
    
    \BITCNT[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_5[2]\, CLR => 
        HWRES_c_34, Q => \BITCNT[2]_net_1\);
    
    un1_hwres_12 : NOR2FT
      port map(A => HWRES_c_0_6_0, B => REG(235), Y => 
        un1_hwres_12_i);
    
    SWORD_7 : MUX2H
      port map(A => \SWORD[3]_net_1\, B => \SWORD_6[3]_net_1\, S
         => un1_sstate_16, Y => \SWORD_7\);
    
    un15_sync_15 : NAND2
      port map(A => \un15_sync_1[15]\, B => \un15_sync_2[15]\, Y
         => \un15_sync[15]\);
    
    \SYNC_5[11]\ : MUX2H
      port map(A => N_274, B => \un15_sync[11]\, S => 
        \sstate_2[0]_net_1\, Y => N_292);
    
    un15_sync_12 : NAND2
      port map(A => \un15_sync_1[12]\, B => \un15_sync_2[15]\, Y
         => \un15_sync[12]\);
    
    \SYNC_5_s[9]\ : OR2FT
      port map(A => sstate_0_sqmuxa, B => N_290, Y => 
        \SYNC_5[9]_net_1\);
    
    \DACRdPnt[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \DACRdPnt_2[0]_net_1\, CLR
         => HWRES_c_34, Q => \DACCFG_RAD[0]\);
    
    \SYNC_5_0[2]\ : MUX2H
      port map(A => \SYNC_c[2]\, B => REG(235), S => 
        \sstate[6]_net_1\, Y => N_265);
    
    \SWORD[5]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_9\, CLR => HWRES_c_36, 
        Q => \SWORD[5]_net_1\);
    
    un15_sync_13_1 : NOR2FT
      port map(A => \DACCFG_RAD[0]\, B => \DACCFG_RAD[1]\, Y => 
        \un15_sync_1[13]\);
    
    un1_sstate_13_0_o3 : NOR2
      port map(A => N_208, B => \sstate_2[0]_net_1\, Y => N_207);
    
    SWORD_5 : MUX2H
      port map(A => \SWORD[1]_net_1\, B => \SWORD_6[1]_net_1\, S
         => un1_sstate_16, Y => \SWORD_5\);
    
    \SYNC_1[11]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[11]_net_1\, CLR => 
        un1_hwres_16_i, SET => un1_reg_9_i, Q => \SYNC_c[11]\);
    
    \SWORD_6_0[4]\ : MUX2H
      port map(A => REG(253), B => DACCFG_DT(4), S => 
        \sstate_1[0]_net_1\, Y => N_353);
    
    \SYNC_5_0[0]\ : MUX2H
      port map(A => \SYNC_c[0]\, B => REG(233), S => 
        \sstate[6]_net_1\, Y => N_263);
    
    \SWORD_6_0[9]\ : MUX2H
      port map(A => REG(258), B => DACCFG_DT(9), S => 
        \sstate_1[0]_net_1\, Y => N_358);
    
    ISI_20 : MUX2H
      port map(A => ISI_6, B => \SDIN_DAC_c\, S => N_201, Y => 
        \ISI_20\);
    
    \SWORD_6_0[8]\ : MUX2H
      port map(A => REG(257), B => DACCFG_DT(8), S => 
        \sstate_1[0]_net_1\, Y => N_357);
    
    \SYNC_5_s[12]\ : OR2FT
      port map(A => sstate_0_sqmuxa, B => N_293, Y => 
        \SYNC_5[12]_net_1\);
    
    \SYNC_1[5]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[5]_net_1\, CLR => 
        un1_hwres_11_i, SET => un1_reg_12_i, Q => \SYNC_c[5]\);
    
    un15_sync_3_1 : NOR2
      port map(A => \DACCFG_RAD[2]\, B => \DACCFG_RAD[3]\, Y => 
        \un15_sync_1[3]\);
    
    \SYNC_5_0[8]\ : MUX2H
      port map(A => \SYNC_c[8]\, B => REG(241), S => 
        \sstate_1[6]_net_1\, Y => N_271);
    
    \SYNC_5_0[10]\ : MUX2H
      port map(A => \SYNC_c[10]\, B => REG(243), S => 
        \sstate_1[6]_net_1\, Y => N_273);
    
    LastDac_1_sqmuxa : AND2
      port map(A => \sstate[2]_net_1\, B => \un15_sync[15]\, Y
         => LastDac_1_sqmuxa_i);
    
    \SYNC_5_s[4]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_285, Y => 
        \SYNC_5[4]_net_1\);
    
    \SYNC_5_0[14]\ : MUX2H
      port map(A => \SYNC_c[14]\, B => REG(247), S => 
        \sstate_1[6]_net_1\, Y => N_277);
    
    \SYNC_1[8]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[8]_net_1\, CLR => 
        un1_hwres_1_i, SET => un1_reg_6_i, Q => \SYNC_c[8]\);
    
    un6_bitcnt : NAND2FT
      port map(A => \LastDac\, B => \RefreshCycle\, Y => 
        \un6_bitcnt\);
    
    \SWORD[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_4\, CLR => HWRES_c_35, 
        Q => \SWORD[0]_net_1\);
    
    \SYNC_5[3]\ : MUX2H
      port map(A => N_266, B => \un15_sync[3]\, S => 
        \sstate[0]_net_1\, Y => N_284);
    
    \SYNC_5_0[4]\ : MUX2H
      port map(A => \SYNC_c[4]\, B => REG(237), S => 
        \sstate[6]_net_1\, Y => N_267);
    
    un15_sync_13 : NAND2
      port map(A => \un15_sync_1[13]\, B => \un15_sync_2[15]\, Y
         => \un15_sync[13]\);
    
    \SWORD[1]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_5\, CLR => HWRES_c_35, 
        Q => \SWORD[1]_net_1\);
    
    un1_reg_9 : AND2
      port map(A => HWRES_c_2, B => REG(244), Y => un1_reg_9_i);
    
    SWORD_0_sqmuxa_0_o2 : AND2
      port map(A => PULSE(9), B => \sstate_0[6]_net_1\, Y => 
        N_208);
    
    un1_hwres_4 : NOR2FT
      port map(A => HWRES_c_0, B => REG(248), Y => un1_hwres_4_i);
    
    SWORD_11 : MUX2H
      port map(A => \SWORD[7]_net_1\, B => \SWORD_6[7]_net_1\, S
         => un1_sstate_16, Y => \SWORD_11\);
    
    \sstate_ns[4]\ : OAI21
      port map(A => ISI_0_sqmuxa, B => \un6_bitcnt\, C => 
        sstate_0_sqmuxa, Y => \sstate_ns[4]_net_1\);
    
    un1_hwres_13 : NOR2FT
      port map(A => HWRES_c_1, B => REG(234), Y => un1_hwres_13_i);
    
    \SYNC_5_0[7]\ : MUX2H
      port map(A => \SYNC_c[7]\, B => REG(240), S => 
        \sstate[6]_net_1\, Y => N_270);
    
    \SWORD_6[12]\ : MUX2H
      port map(A => N_361, B => \SWORD[11]_net_1\, S => 
        \sstate_0[5]_net_1\, Y => \SWORD_6[12]_net_1\);
    
    \SYNC_5[2]\ : MUX2H
      port map(A => N_265, B => \un15_sync[2]\, S => 
        \sstate[0]_net_1\, Y => N_283);
    
    \SWORD[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_6\, CLR => HWRES_c_36, 
        Q => \SWORD[2]_net_1\);
    
    un1_hwres_10 : NOR2FT
      port map(A => HWRES_c_0_6_0, B => REG(243), Y => 
        un1_hwres_10_i);
    
    un15_sync_4 : NAND2
      port map(A => \un15_sync_1[7]\, B => \un15_sync_1[12]\, Y
         => \un15_sync[4]\);
    
    \sstate[2]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate_ns[4]_net_1\, CLR => 
        HWRES_c_36_0, Q => \sstate[2]_net_1\);
    
    SWORD_13 : MUX2H
      port map(A => \SWORD[9]_net_1\, B => \SWORD_6[9]_net_1\, S
         => \un1_sstate_16_0\, Y => \SWORD_13\);
    
    \sstate[5]\ : DFFC
      port map(CLK => CLK_c_c, D => N_191_i_0, CLR => HWRES_c, Q
         => \sstate[5]_net_1\);
    
    ISI : DFFC
      port map(CLK => CLK_c_c, D => \ISI_20\, CLR => HWRES_c_35, 
        Q => \SDIN_DAC_c\);
    
    un1_reg_8 : AND2
      port map(A => HWRES_c_2, B => REG(234), Y => un1_reg_8_i);
    
    \SYNC_5[6]\ : MUX2H
      port map(A => N_269, B => \un15_sync[6]\, S => 
        \sstate[0]_net_1\, Y => N_287);
    
    SWORD_14 : MUX2H
      port map(A => \SWORD[10]_net_1\, B => \SWORD_6[10]_net_1\, 
        S => \un1_sstate_16_0\, Y => \SWORD_14\);
    
    DACCFG_nRD_1 : MUX2H
      port map(A => DACCFG_nRD_net_1, B => \sstate_i_0[2]\, S => 
        N_218, Y => \DACCFG_nRD_1\);
    
    \SYNC_5_s[11]\ : OR2FT
      port map(A => sstate_0_sqmuxa, B => N_292, Y => 
        \SYNC_5[11]_net_1\);
    
    sstate_0_sqmuxa_0_a3_0 : OR2FT
      port map(A => \sstate_0[6]_net_1\, B => N_364, Y => 
        sstate_0_sqmuxa_0);
    
    \SYNC_5[4]\ : MUX2H
      port map(A => N_267, B => \un15_sync[4]\, S => 
        \sstate[0]_net_1\, Y => N_285);
    
    \sstate_ns_i_1_0[1]\ : OR3FTT
      port map(A => N_191_1, B => \sstate_0[5]_net_1\, C => 
        \sstate[4]_net_1\, Y => \sstate_ns_i_1_i[1]\);
    
    \sstate_0[5]\ : DFFC
      port map(CLK => CLK_c_c, D => N_191_i_0, CLR => HWRES_c, Q
         => \sstate_0[5]_net_1\);
    
    \SYNC_5_s[8]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_289, Y => 
        \SYNC_5[8]_net_1\);
    
    \SYNC_5_0[6]\ : MUX2H
      port map(A => \SYNC_c[6]\, B => REG(239), S => 
        \sstate[6]_net_1\, Y => N_269);
    
    \SWORD_6[8]\ : MUX2H
      port map(A => N_357, B => \SWORD[7]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[8]_net_1\);
    
    un1_BITCNT_I_17 : XOR2
      port map(A => \BITCNT[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_17);
    
    un1_sstate_16_0 : OR2FT
      port map(A => N_207, B => \sstate_0[5]_net_1\, Y => 
        un1_sstate_16);
    
    un1_hwres_14 : NOR2FT
      port map(A => HWRES_c_1, B => REG(237), Y => un1_hwres_14_i);
    
    un1_BITCNT_I_15 : XOR2
      port map(A => \BITCNT[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_15);
    
    un1_sstate_17_i_a3_1 : OR2
      port map(A => \sstate_0[0]_net_1\, B => \sstate[3]_net_1\, 
        Y => N_225_1);
    
    un15_sync_2 : NAND2
      port map(A => \un15_sync_1[3]\, B => \un15_sync_1[14]\, Y
         => \un15_sync[2]\);
    
    \sstate_ns_i[1]\ : AND3FTT
      port map(A => \sstate_ns_i_1_i[1]\, B => 
        \sstate_ns_i_a3[1]_net_1\, C => ISI_0_sqmuxa, Y => 
        N_191_i_0);
    
    un1_reg_2 : AND2
      port map(A => HWRES_c_2, B => REG(240), Y => un1_reg_2_i);
    
    un1_hwres_2 : NOR2FT
      port map(A => HWRES_c_0_6_0, B => REG(247), Y => 
        un1_hwres_2_i);
    
    un15_sync_14_1 : NOR2FT
      port map(A => \DACCFG_RAD[1]\, B => \DACCFG_RAD[0]\, Y => 
        \un15_sync_1[14]\);
    
    \SWORD_6_0[15]\ : MUX2H
      port map(A => REG(264), B => DACCFG_DT(15), S => 
        \sstate_0[0]_net_1\, Y => N_314);
    
    un15_sync_7 : NAND2
      port map(A => \un15_sync_1[7]\, B => \un15_sync_1[15]\, Y
         => \un15_sync[7]\);
    
    \SYNC_5_s[13]\ : OR2FT
      port map(A => sstate_0_sqmuxa, B => N_294, Y => 
        \SYNC_5[13]_net_1\);
    
    \SWORD_6[1]\ : MUX2H
      port map(A => N_350, B => \SWORD[0]_net_1\, S => 
        \sstate[5]_net_1\, Y => \SWORD_6[1]_net_1\);
    
    SWORD_16 : MUX2H
      port map(A => \SWORD[12]_net_1\, B => \SWORD_6[12]_net_1\, 
        S => \un1_sstate_16_0\, Y => \SWORD_16\);
    
    \SWORD[13]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_17\, CLR => HWRES_c_35, 
        Q => \SWORD[13]_net_1\);
    
    un1_reg_10 : AND2
      port map(A => HWRES_c_2, B => REG(237), Y => un1_reg_10_i);
    
    \SWORD_6[11]\ : MUX2H
      port map(A => N_360, B => \SWORD[10]_net_1\, S => 
        \sstate_0[5]_net_1\, Y => \SWORD_6[11]_net_1\);
    
    RefreshCycle : DFFC
      port map(CLK => CLK_c_c, D => \RefreshCycle_3\, CLR => 
        HWRES_c_35, Q => \RefreshCycle\);
    
    LastDac : DFFC
      port map(CLK => CLK_c_c, D => \LastDac_21\, CLR => 
        HWRES_c_35, Q => \LastDac\);
    
    un1_sstate_16_0_0 : OR2FT
      port map(A => N_207, B => \sstate_0[5]_net_1\, Y => 
        \un1_sstate_16_0\);
    
    \DACRdPnt_2[2]\ : NOR2FT
      port map(A => I_18_0, B => \sstate_0[6]_net_1\, Y => 
        \DACRdPnt_2[2]_net_1\);
    
    \BITCNT[3]\ : DFFC
      port map(CLK => CLK_c_c, D => \BITCNT_5[3]\, CLR => 
        HWRES_c_34, Q => \BITCNT[3]_net_1\);
    
    un1_BITCNT_I_11 : XOR2
      port map(A => \BITCNT[0]_net_1\, B => \un1_sstate_17_i_a3\, 
        Y => \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \sstate_2[0]\ : DFFC
      port map(CLK => CLK_c_c, D => \sstate[1]_net_1\, CLR => 
        HWRES_c_36_0, Q => \sstate_2[0]_net_1\);
    
    \SYNC_5[1]\ : MUX2H
      port map(A => N_264, B => \un15_sync[1]\, S => 
        \sstate[0]_net_1\, Y => N_282);
    
    SWORD_10 : MUX2H
      port map(A => \SWORD[6]_net_1\, B => \SWORD_6[6]_net_1\, S
         => un1_sstate_16, Y => \SWORD_10\);
    
    \SYNC_5_0[12]\ : MUX2H
      port map(A => \SYNC_c[12]\, B => REG(245), S => 
        \sstate_1[6]_net_1\, Y => N_275);
    
    un1_reg_6 : AND2
      port map(A => HWRES_c_2, B => REG(241), Y => un1_reg_6_i);
    
    un15_sync_8 : NAND2
      port map(A => \un15_sync_1[11]\, B => \un15_sync_1[12]\, Y
         => \un15_sync[8]\);
    
    un1_hwres_3 : NOR2FT
      port map(A => HWRES_c_1, B => REG(246), Y => un1_hwres_3_i);
    
    \SWORD[11]\ : DFFC
      port map(CLK => CLK_c_c, D => \SWORD_15\, CLR => HWRES_c_35, 
        Q => \SWORD[11]_net_1\);
    
    \SWORD_6[15]\ : MUX2H
      port map(A => N_314, B => \SWORD[14]_net_1\, S => 
        \sstate_0[5]_net_1\, Y => \SWORD_6[15]_net_1\);
    
    un15_sync_10 : NAND2
      port map(A => \un15_sync_1[11]\, B => \un15_sync_1[14]\, Y
         => \un15_sync[10]\);
    
    ISI_6_iv_0 : AOI21TTF
      port map(A => \SWORD[15]_net_1\, B => \sstate[3]_net_1\, C
         => \DACCFG_DT_m[15]_net_1\, Y => \ISI_6_iv_0\);
    
    \SYNC_5_s[3]\ : OR2FT
      port map(A => sstate_0_sqmuxa_0, B => N_284, Y => 
        \SYNC_5[3]_net_1\);
    
    un15_sync_3 : NAND2
      port map(A => \un15_sync_1[3]\, B => \un15_sync_1[15]\, Y
         => \un15_sync[3]\);
    
    RefreshCycle_3 : MUX2H
      port map(A => \RefreshCycle\, B => N_364_i_0, S => 
        \sstate_1[6]_net_1\, Y => \RefreshCycle_3\);
    
    \SWORD_6_0[3]\ : MUX2H
      port map(A => REG(252), B => DACCFG_DT(3), S => 
        \sstate_1[0]_net_1\, Y => N_352);
    
    un1_BITCNT_I_21 : AND2
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \BITCNT[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    un1_sstate_17_i_a3 : OR2
      port map(A => N_208, B => N_225_1, Y => 
        \un1_sstate_17_i_a3\);
    
    un1_hwres_16 : NOR2FT
      port map(A => HWRES_c_1, B => REG(244), Y => un1_hwres_16_i);
    
    \SYNC_1[2]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[2]_net_1\, CLR => 
        un1_hwres_12_i, SET => un1_reg_1_i, Q => \SYNC_c[2]\);
    
    un1_reg_14 : AND2
      port map(A => HWRES_c_3, B => REG(243), Y => un1_reg_14_i);
    
    un1_reg_7 : AND2
      port map(A => HWRES_c_2, B => REG(233), Y => un1_reg_7_i);
    
    un1_hwres_1 : NOR2FT
      port map(A => HWRES_c_1, B => REG(241), Y => un1_hwres_1_i);
    
    \SYNC_1[1]\ : DFFB
      port map(CLK => CLK_c_c, D => \SYNC_5[1]_net_1\, CLR => 
        un1_hwres_13_i, SET => un1_reg_8_i, Q => \SYNC_c[1]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity DACCFG is

    port( DACCFG_WDT : in    std_logic_vector(13 downto 4);
          DACCFG_RAD : in    std_logic_vector(3 downto 0);
          DACCFG_DT  : out   std_logic_vector(15 downto 0);
          CROMWAD    : in    std_logic_vector(4 downto 1);
          DACCFG_nRD : in    std_logic;
          DACCFG_nWR : in    std_logic;
          CLK_c_c    : in    std_logic
        );

end DACCFG;

architecture DEF_ARCH of DACCFG is 

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component RAM256x9SSTP
    generic (MEMORYFILE:string := "");

    port( DO8    : out   std_logic;
          DO7    : out   std_logic;
          DO6    : out   std_logic;
          DO5    : out   std_logic;
          DO4    : out   std_logic;
          DO3    : out   std_logic;
          DO2    : out   std_logic;
          DO1    : out   std_logic;
          DO0    : out   std_logic;
          DOS    : out   std_logic;
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          DI8    : in    std_logic := 'U';
          DI7    : in    std_logic := 'U';
          DI6    : in    std_logic := 'U';
          DI5    : in    std_logic := 'U';
          DI4    : in    std_logic := 'U';
          DI3    : in    std_logic := 'U';
          DI2    : in    std_logic := 'U';
          DI1    : in    std_logic := 'U';
          DI0    : in    std_logic := 'U';
          WRB    : in    std_logic := 'U';
          RDB    : in    std_logic := 'U';
          WBLKB  : in    std_logic := 'U';
          RBLKB  : in    std_logic := 'U';
          PARODD : in    std_logic := 'U';
          WCLKS  : in    std_logic := 'U';
          RCLKS  : in    std_logic := 'U';
          DIS    : in    std_logic := 'U'
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \CROMWAD_i_0[4]\, M1_DO8, net00020, \GND\, M0_DO8_0, 
        net00019, \VCC\ : std_logic;

begin 


    PWR_i : PWR
      port map(Y => \VCC\);
    
    M1 : RAM256x9SSTP
      generic map(MEMORYFILE => "DACCFG_M1.mem")

      port map(DO8 => M1_DO8, DO7 => DACCFG_DT(15), DO6 => 
        DACCFG_DT(14), DO5 => DACCFG_DT(13), DO4 => DACCFG_DT(12), 
        DO3 => DACCFG_DT(11), DO2 => DACCFG_DT(10), DO1 => 
        DACCFG_DT(9), DO0 => DACCFG_DT(8), DOS => net00020, 
        WADDR7 => \GND\, WADDR6 => \GND\, WADDR5 => \GND\, WADDR4
         => \GND\, WADDR3 => \CROMWAD_i_0[4]\, WADDR2 => 
        CROMWAD(3), WADDR1 => CROMWAD(2), WADDR0 => CROMWAD(1), 
        RADDR7 => \GND\, RADDR6 => \GND\, RADDR5 => \GND\, RADDR4
         => \GND\, RADDR3 => DACCFG_RAD(3), RADDR2 => 
        DACCFG_RAD(2), RADDR1 => DACCFG_RAD(1), RADDR0 => 
        DACCFG_RAD(0), DI8 => \GND\, DI7 => \GND\, DI6 => \GND\, 
        DI5 => DACCFG_WDT(13), DI4 => DACCFG_WDT(12), DI3 => 
        DACCFG_WDT(11), DI2 => DACCFG_WDT(10), DI1 => 
        DACCFG_WDT(9), DI0 => DACCFG_WDT(8), WRB => DACCFG_nWR, 
        RDB => DACCFG_nRD, WBLKB => \GND\, RBLKB => \GND\, PARODD
         => \GND\, WCLKS => CLK_c_c, RCLKS => CLK_c_c, DIS => 
        \GND\);
    
    M0 : RAM256x9SSTP
      generic map(MEMORYFILE => "DACCFG_M0.mem")

      port map(DO8 => M0_DO8_0, DO7 => DACCFG_DT(7), DO6 => 
        DACCFG_DT(6), DO5 => DACCFG_DT(5), DO4 => DACCFG_DT(4), 
        DO3 => DACCFG_DT(3), DO2 => DACCFG_DT(2), DO1 => 
        DACCFG_DT(1), DO0 => DACCFG_DT(0), DOS => net00019, 
        WADDR7 => \GND\, WADDR6 => \GND\, WADDR5 => \GND\, WADDR4
         => \GND\, WADDR3 => \CROMWAD_i_0[4]\, WADDR2 => 
        CROMWAD(3), WADDR1 => CROMWAD(2), WADDR0 => CROMWAD(1), 
        RADDR7 => \GND\, RADDR6 => \GND\, RADDR5 => \GND\, RADDR4
         => \GND\, RADDR3 => DACCFG_RAD(3), RADDR2 => 
        DACCFG_RAD(2), RADDR1 => DACCFG_RAD(1), RADDR0 => 
        DACCFG_RAD(0), DI8 => \GND\, DI7 => DACCFG_WDT(7), DI6
         => DACCFG_WDT(6), DI5 => DACCFG_WDT(5), DI4 => 
        DACCFG_WDT(4), DI3 => \GND\, DI2 => \GND\, DI1 => \GND\, 
        DI0 => \GND\, WRB => DACCFG_nWR, RDB => DACCFG_nRD, WBLKB
         => \GND\, RBLKB => \GND\, PARODD => \GND\, WCLKS => 
        CLK_c_c, RCLKS => CLK_c_c, DIS => \GND\);
    
    M1_i : INV
      port map(A => CROMWAD(4), Y => \CROMWAD_i_0[4]\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity v1392ltm is

    port( ALICLK      : in    std_logic;
          AMB         : in    std_logic_vector(5 downto 0);
          ASB         : in    std_logic;
          BERRVME     : in    std_logic;
          BNCRES      : in    std_logic;
          DS0B        : in    std_logic;
          DS1B        : in    std_logic;
          EVRES       : in    std_logic;
          F_SO        : in    std_logic;
          GA          : in    std_logic_vector(3 downto 0);
          IACKB       : in    std_logic;
          IACKINB     : in    std_logic;
          L0          : in    std_logic;
          L1A         : in    std_logic;
          L1R         : in    std_logic;
          L2A         : in    std_logic;
          L2R         : in    std_logic;
          LCLK        : in    std_logic;
          LOS         : in    std_logic;
          NLBPCKE     : in    std_logic;
          NLBPCKR     : in    std_logic;
          NPWON       : in    std_logic;
          PSM_SP0     : in    std_logic;
          PSM_SP1     : in    std_logic;
          PSM_SP2     : in    std_logic;
          PSM_SP3     : in    std_logic;
          PSM_SP4     : in    std_logic;
          PSM_SP5     : in    std_logic;
          SPULSE0     : in    std_logic;
          SPULSE1     : in    std_logic;
          SPULSE2     : in    std_logic;
          SYSRESB     : in    std_logic;
          WRITEB      : in    std_logic;
          nLBRDY      : in    std_logic;
          ADLTC       : out   std_logic;
          AE_PDL      : out   std_logic_vector(47 downto 0);
          APACLK0     : out   std_logic;
          DIR_CTTM    : out   std_logic_vector(7 downto 0);
          FCS         : out   std_logic;
          F_SCK       : out   std_logic;
          F_SI        : out   std_logic;
          IACKOUTB    : out   std_logic;
          INTR1       : out   std_logic;
          INTR2       : out   std_logic;
          LED         : out   std_logic_vector(5 downto 0);
          LTM_BUSY    : out   std_logic;
          LTM_DRDY    : out   std_logic;
          MD_PDL      : out   std_logic;
          MYBERR      : out   std_logic;
          NDTKIN      : out   std_logic;
          NLBCLR      : out   std_logic;
          NLBCS       : out   std_logic;
          NLBRD       : out   std_logic;
          NLBRES      : out   std_logic;
          NLBWAIT     : out   std_logic;
          NOE16R      : out   std_logic;
          NOE16W      : out   std_logic;
          NOE32R      : out   std_logic;
          NOE32W      : out   std_logic;
          NOE64R      : out   std_logic;
          NOEAD       : out   std_logic;
          NOEDTK      : out   std_logic;
          NSELCLK     : out   std_logic;
          PSM_RES     : out   std_logic;
          P_PDL       : out   std_logic_vector(7 downto 1);
          RSELA0      : out   std_logic;
          RSELA1      : out   std_logic;
          RSELB0      : out   std_logic;
          RSELB1      : out   std_logic;
          RSELC0      : out   std_logic;
          RSELC1      : out   std_logic;
          RSELD0      : out   std_logic;
          RSELD1      : out   std_logic;
          SCL0        : out   std_logic;
          SCL1        : out   std_logic;
          SCLK_DAC    : out   std_logic;
          SCLK_PDL    : out   std_logic;
          SDIN_DAC    : out   std_logic;
          SELCLK      : out   std_logic;
          SI_PDL      : out   std_logic;
          SYNC        : out   std_logic_vector(15 downto 0);
          TST         : out   std_logic_vector(15 downto 0);
          nLBAS       : out   std_logic;
          LB          : inout std_logic_vector(31 downto 0) := (others => 'Z');
          LBSP        : inout std_logic_vector(31 downto 0) := (others => 'Z');
          LWORDB      : inout std_logic := 'Z';
          NCYC_RELOAD : inout std_logic := 'Z';
          NLBLAST     : out   std_logic;
          SDA0        : inout std_logic := 'Z';
          SDA1        : inout std_logic := 'Z';
          SP_PDL      : inout std_logic_vector(47 downto 0) := (others => 'Z');
          VAD         : inout std_logic_vector(31 downto 1) := (others => 'Z');
          VDB         : inout std_logic_vector(31 downto 0) := (others => 'Z')
        );

end v1392ltm;

architecture DEF_ARCH of v1392ltm is 

  component BFR
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OB33PH
    port( PAD : out   std_logic;
          A   : in    std_logic := 'U'
        );
  end component;

  component IOB33PH
    port( PAD : inout   std_logic;
          A   : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GL33
    port( PAD : in    std_logic := 'U';
          GL  : out   std_logic
        );
  end component;

  component OTB33PH
    port( PAD : out   std_logic;
          A   : in    std_logic := 'U';
          EN  : in    std_logic := 'U'
        );
  end component;

  component IB33
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component PDL_INTERF
    port( PULSE         : in    std_logic_vector(8 to 8) := (others => 'U');
          P_PDL_c       : out   std_logic_vector(7 downto 1);
          PDL_RDATA     : out   std_logic_vector(7 downto 0);
          PDL_RADDR     : in    std_logic_vector(5 downto 0) := (others => 'U');
          PDLCFG_RAD    : out   std_logic_vector(5 downto 0);
          PDLCFG_DT     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PDLCFG_DT_0_0 : in    std_logic_vector(0 to 0) := (others => 'U');
          PDLCFG_DT_3   : in    std_logic_vector(0 to 0) := (others => 'U');
          PDLCFG_DT_1   : in    std_logic_vector(0 to 0) := (others => 'U');
          PDLCFG_DT_2   : in    std_logic_vector(0 to 0) := (others => 'U');
          PDLCFG_DT_0   : in    std_logic_vector(0 to 0) := (others => 'U');
          P0            : out   std_logic_vector(47 downto 0);
          AE_PDL_c      : out   std_logic_vector(47 downto 0);
          SP_PDL_in     : in    std_logic_vector(47 downto 0) := (others => 'U');
          REG_0         : in    std_logic_vector(127 downto 124) := (others => 'U');
          REG_i_0       : in    std_logic_vector(121 to 121) := (others => 'U');
          REG_32        : in    std_logic := 'U';
          REG_33        : in    std_logic := 'U';
          REG_34        : in    std_logic := 'U';
          REG_35        : in    std_logic := 'U';
          REG_36        : in    std_logic := 'U';
          REG_37        : in    std_logic := 'U';
          REG_38        : in    std_logic := 'U';
          REG_39        : in    std_logic := 'U';
          REG_40        : in    std_logic := 'U';
          REG_41        : in    std_logic := 'U';
          REG_42        : in    std_logic := 'U';
          REG_43        : in    std_logic := 'U';
          REG_44        : in    std_logic := 'U';
          REG_45        : in    std_logic := 'U';
          REG_46        : in    std_logic := 'U';
          REG_47        : in    std_logic := 'U';
          REG_48        : in    std_logic := 'U';
          REG_49        : in    std_logic := 'U';
          REG_50        : in    std_logic := 'U';
          REG_51        : in    std_logic := 'U';
          REG_52        : in    std_logic := 'U';
          REG_53        : in    std_logic := 'U';
          REG_54        : in    std_logic := 'U';
          REG_55        : in    std_logic := 'U';
          REG_56        : in    std_logic := 'U';
          REG_57        : in    std_logic := 'U';
          REG_58        : in    std_logic := 'U';
          REG_59        : in    std_logic := 'U';
          REG_60        : in    std_logic := 'U';
          REG_61        : in    std_logic := 'U';
          REG_62        : in    std_logic := 'U';
          REG_63        : in    std_logic := 'U';
          REG_64        : in    std_logic := 'U';
          REG_65        : in    std_logic := 'U';
          REG_66        : in    std_logic := 'U';
          REG_67        : in    std_logic := 'U';
          REG_68        : in    std_logic := 'U';
          REG_69        : in    std_logic := 'U';
          REG_70        : in    std_logic := 'U';
          REG_71        : in    std_logic := 'U';
          REG_72        : in    std_logic := 'U';
          REG_73        : in    std_logic := 'U';
          REG_74        : in    std_logic := 'U';
          REG_75        : in    std_logic := 'U';
          REG_76        : in    std_logic := 'U';
          REG_77        : in    std_logic := 'U';
          REG_78        : in    std_logic := 'U';
          REG_79        : in    std_logic := 'U';
          REG_3         : in    std_logic := 'U';
          REG_6         : in    std_logic := 'U';
          REG_5         : in    std_logic := 'U';
          REG_4         : in    std_logic := 'U';
          REG_2         : in    std_logic := 'U';
          REG_1         : in    std_logic := 'U';
          REG_24        : out   std_logic;
          REG_9         : in    std_logic := 'U';
          REG_16        : out   std_logic;
          REG_10        : in    std_logic := 'U';
          REG_17        : out   std_logic;
          REG_11        : in    std_logic := 'U';
          REG_18        : out   std_logic;
          REG_12        : in    std_logic := 'U';
          REG_19        : out   std_logic;
          REG_13        : in    std_logic := 'U';
          REG_20        : out   std_logic;
          REG_14        : in    std_logic := 'U';
          REG_21        : out   std_logic;
          REG_15        : in    std_logic := 'U';
          REG_22        : out   std_logic;
          REG_23        : out   std_logic;
          REG_0_d0      : in    std_logic := 'U';
          REG_8         : in    std_logic := 'U';
          MD_PDL_c      : out   std_logic;
          PDL_RACK      : out   std_logic;
          PDL_RREQ      : in    std_logic := 'U';
          SI_PDL_c      : out   std_logic;
          PDLCFG_nRD    : out   std_logic;
          SCLK_PDL_c    : out   std_logic;
          HWRES_c_2     : in    std_logic := 'U';
          HWRES_c_1     : in    std_logic := 'U';
          MD_PDL_c_0    : out   std_logic;
          MD_PDL_c_1    : out   std_logic;
          MD_PDL_c_2    : out   std_logic;
          MD_PDL_c_3    : out   std_logic;
          LOAD_RES      : in    std_logic := 'U';
          HWRES_c_0_3   : in    std_logic := 'U';
          HWRES_c_0_2   : in    std_logic := 'U';
          LOAD_RES_3    : in    std_logic := 'U';
          CLK_c_c       : in    std_logic := 'U';
          HWRES_c_23_0  : in    std_logic := 'U';
          HWRES_c_0     : in    std_logic := 'U';
          LOAD_RES_0    : in    std_logic := 'U'
        );
  end component;

  component PDLCFG
    port( CROMWDT       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PDLCFG_RAD    : in    std_logic_vector(5 downto 0) := (others => 'U');
          CROMWAD       : in    std_logic_vector(5 downto 0) := (others => 'U');
          PDLCFG_DT_0   : out   std_logic_vector(0 to 0);
          PDLCFG_DT_1   : out   std_logic_vector(0 to 0);
          PDLCFG_DT_2   : out   std_logic_vector(0 to 0);
          PDLCFG_DT_3   : out   std_logic_vector(0 to 0);
          PDLCFG_DT     : out   std_logic_vector(7 downto 0);
          PDLCFG_DT_0_0 : out   std_logic_vector(0 to 0);
          PDLCFG_nRD    : in    std_logic := 'U';
          PDLCFG_nWR    : in    std_logic := 'U';
          CLK_c_c       : in    std_logic := 'U'
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VINTERF
    port( TICK            : in    std_logic_vector(2 to 2) := (others => 'U');
          RAMDT           : in    std_logic_vector(7 downto 0) := (others => 'U');
          VADm            : out   std_logic_vector(31 downto 0);
          RAMAD_VME       : out   std_logic_vector(8 downto 0);
          AMB_c           : in    std_logic_vector(5 downto 0) := (others => 'U');
          LB_in           : in    std_logic_vector(31 downto 0) := (others => 'U');
          OR_RDATA        : out   std_logic_vector(9 downto 0);
          PULSE_0         : out   std_logic;
          PULSE_1         : out   std_logic;
          PULSE_2         : out   std_logic;
          PULSE_3         : out   std_logic;
          PULSE_6         : out   std_logic;
          PULSE_7         : out   std_logic;
          PULSE_8         : out   std_logic;
          PULSE_9         : out   std_logic;
          PULSE_10        : out   std_logic;
          OR_RADDR        : in    std_logic_vector(5 downto 0) := (others => 'U');
          VDB_in_0        : in    std_logic_vector(15 downto 0) := (others => 'U');
          VDB_in          : in    std_logic_vector(31 downto 0) := (others => 'U');
          LB_i            : out   std_logic_vector(31 downto 0);
          DPR             : in    std_logic_vector(31 downto 0) := (others => 'U');
          FBOUT           : in    std_logic_vector(7 downto 0) := (others => 'U');
          LBSP_c          : in    std_logic_vector(2 to 2) := (others => 'U');
          REGMAP_35       : out   std_logic;
          REGMAP_31       : out   std_logic;
          REG_c_21        : in    std_logic := 'U';
          REG_c_22        : in    std_logic := 'U';
          REG_c_23        : in    std_logic := 'U';
          REG_c_0         : out   std_logic;
          LBSP_in_0       : in    std_logic := 'U';
          LBSP_in_1       : in    std_logic := 'U';
          LBSP_in_15      : in    std_logic := 'U';
          LBSP_in_16      : in    std_logic := 'U';
          LBSP_in_17      : in    std_logic := 'U';
          LBSP_in_18      : in    std_logic := 'U';
          LBSP_in_19      : in    std_logic := 'U';
          LBSP_in_20      : in    std_logic := 'U';
          LBSP_in_21      : in    std_logic := 'U';
          LBSP_in_22      : in    std_logic := 'U';
          LBSP_in_23      : in    std_logic := 'U';
          LBSP_in_24      : in    std_logic := 'U';
          LBSP_in_25      : in    std_logic := 'U';
          LBSP_in_26      : in    std_logic := 'U';
          LBSP_in_27      : in    std_logic := 'U';
          LBSP_in_28      : in    std_logic := 'U';
          LBSP_in_29      : in    std_logic := 'U';
          LBSP_in_30      : in    std_logic := 'U';
          LBSP_in_31      : in    std_logic := 'U';
          VAD_in_0        : in    std_logic := 'U';
          VAD_in_1        : in    std_logic := 'U';
          VAD_in_2        : in    std_logic := 'U';
          VAD_in_3        : in    std_logic := 'U';
          VAD_in_4        : in    std_logic := 'U';
          VAD_in_5        : in    std_logic := 'U';
          VAD_in_6        : in    std_logic := 'U';
          VAD_in_7        : in    std_logic := 'U';
          VAD_in_8        : in    std_logic := 'U';
          VAD_in_9        : in    std_logic := 'U';
          VAD_in_10       : in    std_logic := 'U';
          VAD_in_11       : in    std_logic := 'U';
          VAD_in_12       : in    std_logic := 'U';
          VAD_in_13       : in    std_logic := 'U';
          VAD_in_14       : in    std_logic := 'U';
          VAD_in_27       : in    std_logic := 'U';
          VAD_in_28       : in    std_logic := 'U';
          VAD_in_29       : in    std_logic := 'U';
          VAD_in_30       : in    std_logic := 'U';
          GA_c            : in    std_logic_vector(3 downto 0) := (others => 'U');
          VDBm_0          : out   std_logic;
          VDBm_1          : out   std_logic;
          VDBm_2          : out   std_logic;
          VDBm_3          : out   std_logic;
          VDBm_4          : out   std_logic;
          VDBm_5          : out   std_logic;
          VDBm_6          : out   std_logic;
          VDBm_7          : out   std_logic;
          VDBm_8          : out   std_logic;
          VDBm_9          : out   std_logic;
          VDBm_10         : out   std_logic;
          VDBm_12         : out   std_logic;
          VDBm_13         : out   std_logic;
          VDBm_14         : out   std_logic;
          VDBm_15         : out   std_logic;
          VDBm_16         : out   std_logic;
          VDBm_17         : out   std_logic;
          VDBm_18         : out   std_logic;
          VDBm_19         : out   std_logic;
          VDBm_20         : out   std_logic;
          VDBm_22         : out   std_logic;
          VDBm_23         : out   std_logic;
          VDBm_24         : out   std_logic;
          VDBm_25         : out   std_logic;
          VDBm_26         : out   std_logic;
          VDBm_27         : out   std_logic;
          VDBm_28         : out   std_logic;
          VDBm_29         : out   std_logic;
          VDBm_30         : out   std_logic;
          VDBm_31         : out   std_logic;
          VDBm_i_m2       : out   std_logic_vector(11 to 11);
          REG_126         : out   std_logic;
          REG_125         : out   std_logic;
          REG_124         : out   std_logic;
          REG_123         : out   std_logic;
          REG_344         : out   std_logic;
          REG_345         : out   std_logic;
          REG_359         : out   std_logic;
          REG_360         : out   std_logic;
          REG_361         : out   std_logic;
          REG_362         : out   std_logic;
          REG_363         : out   std_logic;
          REG_364         : out   std_logic;
          REG_365         : out   std_logic;
          REG_366         : out   std_logic;
          REG_367         : out   std_logic;
          REG_368         : out   std_logic;
          REG_369         : out   std_logic;
          REG_370         : out   std_logic;
          REG_371         : out   std_logic;
          REG_372         : out   std_logic;
          REG_373         : out   std_logic;
          REG_374         : out   std_logic;
          REG_375         : out   std_logic;
          REG_408         : out   std_logic;
          REG_480         : out   std_logic;
          REG_80          : out   std_logic;
          REG_81          : out   std_logic;
          REG_82          : out   std_logic;
          REG_83          : out   std_logic;
          REG_84          : out   std_logic;
          REG_85          : out   std_logic;
          REG_86          : out   std_logic;
          REG_87          : out   std_logic;
          REG_88          : out   std_logic;
          REG_89          : out   std_logic;
          REG_90          : out   std_logic;
          REG_96          : out   std_logic;
          REG_97          : out   std_logic;
          REG_98          : out   std_logic;
          REG_99          : out   std_logic;
          REG_100         : out   std_logic;
          REG_101         : out   std_logic;
          REG_102         : out   std_logic;
          REG_103         : out   std_logic;
          REG_376         : out   std_logic;
          REG_120         : out   std_logic;
          REG_152         : out   std_logic;
          REG_232         : out   std_logic;
          REG_248         : out   std_logic;
          REG_168         : out   std_logic;
          REG_184         : out   std_logic;
          REG_104         : in    std_logic := 'U';
          REG_136         : in    std_logic := 'U';
          REG_31          : in    std_logic := 'U';
          REG_47          : out   std_logic;
          REG_440         : out   std_logic;
          REG_456         : in    std_logic := 'U';
          REG_441         : out   std_logic;
          REG_457         : in    std_logic := 'U';
          REG_473         : in    std_logic := 'U';
          REG_121         : out   std_logic;
          REG_153         : out   std_logic;
          REG_233         : out   std_logic;
          REG_249         : out   std_logic;
          REG_169         : out   std_logic;
          REG_185         : out   std_logic;
          REG_105         : in    std_logic := 'U';
          REG_137         : in    std_logic := 'U';
          REG_32          : in    std_logic := 'U';
          REG_16          : in    std_logic := 'U';
          REG_48          : out   std_logic;
          REG_377         : out   std_logic;
          REG_409         : out   std_logic;
          REG_442         : out   std_logic;
          REG_458         : in    std_logic := 'U';
          REG_474         : in    std_logic := 'U';
          REG_378         : out   std_logic;
          REG_410         : out   std_logic;
          REG_154         : out   std_logic;
          REG_170         : out   std_logic;
          REG_122         : out   std_logic;
          REG_250         : out   std_logic;
          REG_138         : in    std_logic := 'U';
          REG_186         : out   std_logic;
          REG_234         : out   std_logic;
          REG_33          : in    std_logic := 'U';
          REG_49          : out   std_logic;
          REG_34          : in    std_logic := 'U';
          REG_50          : out   std_logic;
          REG_155         : out   std_logic;
          REG_171         : out   std_logic;
          REG_251         : out   std_logic;
          REG_139         : in    std_logic := 'U';
          REG_187         : out   std_logic;
          REG_235         : out   std_logic;
          REG_443         : out   std_logic;
          REG_459         : in    std_logic := 'U';
          REG_379         : out   std_logic;
          REG_411         : out   std_logic;
          REG_475         : in    std_logic := 'U';
          REG_51          : out   std_logic;
          REG_35          : in    std_logic := 'U';
          REG_19          : in    std_logic := 'U';
          REG_156         : out   std_logic;
          REG_172         : out   std_logic;
          REG_252         : out   std_logic;
          REG_140         : in    std_logic := 'U';
          REG_188         : out   std_logic;
          REG_236         : out   std_logic;
          REG_332         : in    std_logic := 'U';
          REG_444         : out   std_logic;
          REG_460         : in    std_logic := 'U';
          REG_380         : out   std_logic;
          REG_412         : out   std_logic;
          REG_476         : in    std_logic := 'U';
          REG_445         : out   std_logic;
          REG_461         : in    std_logic := 'U';
          REG_413         : out   std_logic;
          REG_381         : out   std_logic;
          REG_52          : out   std_logic;
          REG_36          : in    std_logic := 'U';
          REG_157         : out   std_logic;
          REG_173         : out   std_logic;
          REG_253         : out   std_logic;
          REG_141         : in    std_logic := 'U';
          REG_189         : out   std_logic;
          REG_237         : out   std_logic;
          REG_333         : in    std_logic := 'U';
          REG_477         : in    std_logic := 'U';
          REG_462         : in    std_logic := 'U';
          REG_478         : in    std_logic := 'U';
          REG_382         : out   std_logic;
          REG_414         : out   std_logic;
          REG_37          : in    std_logic := 'U';
          REG_5           : out   std_logic;
          REG_53          : out   std_logic;
          REG_158         : out   std_logic;
          REG_174         : out   std_logic;
          REG_254         : out   std_logic;
          REG_142         : in    std_logic := 'U';
          REG_190         : out   std_logic;
          REG_238         : out   std_logic;
          REG_334         : in    std_logic := 'U';
          REG_463         : in    std_logic := 'U';
          REG_383         : out   std_logic;
          REG_415         : out   std_logic;
          REG_54          : out   std_logic;
          REG_38          : in    std_logic := 'U';
          REG_159         : out   std_logic;
          REG_175         : out   std_logic;
          REG_255         : out   std_logic;
          REG_143         : in    std_logic := 'U';
          REG_191         : out   std_logic;
          REG_239         : out   std_logic;
          REG_479         : in    std_logic := 'U';
          REG_464         : in    std_logic := 'U';
          REG_416         : out   std_logic;
          REG_39          : in    std_logic := 'U';
          REG_7           : out   std_logic;
          REG_55          : out   std_logic;
          REG_128         : out   std_logic;
          REG_160         : out   std_logic;
          REG_240         : out   std_logic;
          REG_256         : out   std_logic;
          REG_176         : out   std_logic;
          REG_192         : out   std_logic;
          REG_112         : in    std_logic := 'U';
          REG_144         : in    std_logic := 'U';
          REG_465         : in    std_logic := 'U';
          REG_56          : out   std_logic;
          REG_40          : in    std_logic := 'U';
          REG_161         : out   std_logic;
          REG_177         : out   std_logic;
          REG_129         : out   std_logic;
          REG_257         : out   std_logic;
          REG_113         : in    std_logic := 'U';
          REG_193         : out   std_logic;
          REG_241         : out   std_logic;
          REG_417         : out   std_logic;
          REG_466         : in    std_logic := 'U';
          REG_57          : out   std_logic;
          REG_41          : in    std_logic := 'U';
          REG_162         : out   std_logic;
          REG_178         : out   std_logic;
          REG_130         : out   std_logic;
          REG_258         : out   std_logic;
          REG_114         : in    std_logic := 'U';
          REG_194         : out   std_logic;
          REG_242         : out   std_logic;
          REG_418         : out   std_logic;
          REG_467         : in    std_logic := 'U';
          REG_42          : in    std_logic := 'U';
          REG_58          : out   std_logic;
          REG_163         : out   std_logic;
          REG_179         : out   std_logic;
          REG_131         : out   std_logic;
          REG_259         : out   std_logic;
          REG_115         : in    std_logic := 'U';
          REG_195         : out   std_logic;
          REG_243         : out   std_logic;
          REG_419         : out   std_logic;
          REG_468         : in    std_logic := 'U';
          REG_43          : in    std_logic := 'U';
          REG_59          : out   std_logic;
          REG_164         : out   std_logic;
          REG_180         : out   std_logic;
          REG_132         : out   std_logic;
          REG_260         : out   std_logic;
          REG_116         : in    std_logic := 'U';
          REG_196         : out   std_logic;
          REG_244         : out   std_logic;
          REG_420         : out   std_logic;
          REG_469         : in    std_logic := 'U';
          REG_60          : out   std_logic;
          REG_44          : in    std_logic := 'U';
          REG_165         : out   std_logic;
          REG_181         : out   std_logic;
          REG_133         : out   std_logic;
          REG_261         : out   std_logic;
          REG_117         : in    std_logic := 'U';
          REG_197         : out   std_logic;
          REG_245         : out   std_logic;
          REG_421         : out   std_logic;
          REG_470         : in    std_logic := 'U';
          REG_61          : out   std_logic;
          REG_45          : in    std_logic := 'U';
          REG_166         : out   std_logic;
          REG_182         : out   std_logic;
          REG_134         : out   std_logic;
          REG_262         : out   std_logic;
          REG_118         : in    std_logic := 'U';
          REG_198         : out   std_logic;
          REG_246         : out   std_logic;
          REG_422         : out   std_logic;
          REG_455         : out   std_logic;
          REG_471         : in    std_logic := 'U';
          REG_423         : out   std_logic;
          REG_46          : in    std_logic := 'U';
          REG_62          : out   std_logic;
          REG_167         : out   std_logic;
          REG_183         : out   std_logic;
          REG_135         : out   std_logic;
          REG_263         : out   std_logic;
          REG_119         : in    std_logic := 'U';
          REG_199         : out   std_logic;
          REG_247         : out   std_logic;
          REG_63          : out   std_logic;
          REG_424         : out   std_logic;
          REG_64          : out   std_logic;
          REG_425         : out   std_logic;
          REG_65          : out   std_logic;
          REG_426         : out   std_logic;
          REG_66          : out   std_logic;
          REG_427         : out   std_logic;
          REG_67          : out   std_logic;
          REG_428         : out   std_logic;
          REG_68          : out   std_logic;
          REG_429         : out   std_logic;
          REG_69          : out   std_logic;
          REG_430         : out   std_logic;
          REG_70          : out   std_logic;
          REG_431         : out   std_logic;
          REG_71          : out   std_logic;
          REG_432         : out   std_logic;
          REG_72          : out   std_logic;
          REG_433         : out   std_logic;
          REG_73          : out   std_logic;
          REG_434         : out   std_logic;
          REG_74          : out   std_logic;
          REG_435         : out   std_logic;
          REG_75          : out   std_logic;
          REG_436         : out   std_logic;
          REG_76          : out   std_logic;
          REG_437         : out   std_logic;
          REG_77          : out   std_logic;
          REG_438         : out   std_logic;
          REG_78          : out   std_logic;
          REG_439         : out   std_logic;
          REG_4           : out   std_logic;
          REG_79          : out   std_logic;
          TST_c_c         : out   std_logic_vector(3 to 3);
          TST_c_4         : out   std_logic;
          TST_c_0         : out   std_logic;
          TST_c_5         : out   std_logic;
          TST_c_2         : out   std_logic;
          TST_c_1         : out   std_logic;
          REG_i_0_116     : out   std_logic;
          REG_i_0_0       : out   std_logic;
          REG_i_0_75      : out   std_logic;
          REG_i_0_260     : out   std_logic;
          REG_i_0_261     : out   std_logic;
          REG_i_0_275     : out   std_logic;
          REG_i_0_276     : out   std_logic;
          REG_i_0_277     : out   std_logic;
          REG_i_0_278     : out   std_logic;
          REG_i_0_279     : out   std_logic;
          REG_i_0_280     : out   std_logic;
          REG_i_0_281     : out   std_logic;
          REG_i_0_282     : out   std_logic;
          REG_i_0_283     : out   std_logic;
          REG_i_0_284     : out   std_logic;
          REG_i_0_285     : out   std_logic;
          REG_i_0_286     : out   std_logic;
          REG_i_0_287     : out   std_logic;
          REG_i_0_288     : out   std_logic;
          REG_i_0_289     : out   std_logic;
          REG_i_0_290     : out   std_logic;
          REG_i_0_291     : out   std_logic;
          REG_i_0_393     : out   std_logic;
          REG_i_0_391     : out   std_logic;
          REG_i_0_395     : out   std_logic;
          REG_i_0_388     : out   std_logic;
          REG_i_0_389     : out   std_logic;
          REG_i_0_390     : out   std_logic;
          REG_i_0_392     : out   std_logic;
          REG_i_0_394     : out   std_logic;
          REG_0           : out   std_logic_vector(127 downto 124);
          HWRES_c_16      : in    std_logic := 'U';
          HWRES_c_15      : in    std_logic := 'U';
          CLEAR_22        : in    std_logic := 'U';
          CLEAR_21        : in    std_logic := 'U';
          CLEAR_25        : in    std_logic := 'U';
          CLEAR_24        : in    std_logic := 'U';
          CLEAR_23        : in    std_logic := 'U';
          CLEAR_27        : in    std_logic := 'U';
          CLEAR_26        : in    std_logic := 'U';
          HWRES_c_18      : in    std_logic := 'U';
          HWRES_c_22      : in    std_logic := 'U';
          CLEAR_28        : in    std_logic := 'U';
          CLEAR           : in    std_logic := 'U';
          HWRES_c_17      : in    std_logic := 'U';
          HWRES_c_21      : in    std_logic := 'U';
          HWRES_c_12      : in    std_logic := 'U';
          HWRES_c_23      : in    std_logic := 'U';
          RAMRD           : out   std_logic;
          HWRES_c_19      : in    std_logic := 'U';
          OR_RACK         : out   std_logic;
          HWRES_c_14      : in    std_logic := 'U';
          OR_RREQ         : in    std_logic := 'U';
          HWRES_c_20      : in    std_logic := 'U';
          EF              : in    std_logic := 'U';
          CLEAR_20        : in    std_logic := 'U';
          ASB_c           : in    std_logic := 'U';
          un5_noe16ri_0_0 : out   std_logic;
          un7_noe32ri_0_0 : out   std_logic;
          WRITEB_c        : in    std_logic := 'U';
          nLBAS_c         : out   std_logic;
          LB_nOE          : out   std_logic;
          LWORDB_in       : in    std_logic := 'U';
          MYBERR_c        : out   std_logic;
          IACKB_c         : in    std_logic := 'U';
          nLBRDY_c        : in    std_logic := 'U';
          FWIMG2LOAD      : out   std_logic;
          NLBLAST_c       : out   std_logic;
          NLBRD_c         : out   std_logic;
          NLBCLR_c        : in    std_logic := 'U';
          EVREAD          : out   std_logic;
          NRDMEB          : out   std_logic;
          DTEST_FIFO      : in    std_logic := 'U';
          RUN_c           : out   std_logic;
          N_2052          : out   std_logic;
          d_m7            : in    std_logic := 'U';
          EV_RES_c        : in    std_logic := 'U';
          L0_c_c          : in    std_logic := 'U';
          L1A_c_c         : in    std_logic := 'U';
          L1R_c_c         : in    std_logic := 'U';
          L2A_c_c         : in    std_logic := 'U';
          L2R_c_c         : in    std_logic := 'U';
          LOS_c_c         : in    std_logic := 'U';
          N_441           : out   std_logic;
          SPULSE0_c_c     : in    std_logic := 'U';
          SPULSE1_c_c     : in    std_logic := 'U';
          SPULSE2_c_c     : in    std_logic := 'U';
          DS1B_c          : in    std_logic := 'U';
          DS0B_c          : in    std_logic := 'U';
          N_500           : out   std_logic;
          NDTKIN_c        : out   std_logic;
          NOE16W_c        : out   std_logic;
          NOE32W_c        : out   std_logic;
          NOEAD_c         : out   std_logic;
          NSELCLK_c       : out   std_logic;
          NSELCLK_c_i_0   : out   std_logic;
          CLEAR_0         : in    std_logic := 'U';
          EVRDY_c         : in    std_logic := 'U';
          HWRES_c_1       : in    std_logic := 'U';
          NOEAD_c_i_0     : out   std_logic;
          N_2613_0        : out   std_logic;
          RUN_c_0         : out   std_logic;
          HWRES_c_0       : in    std_logic := 'U';
          NOEAD_c_0       : out   std_logic;
          NOEAD_c_1       : out   std_logic;
          HWRES_c_22_0    : in    std_logic := 'U';
          ALICLK_c        : in    std_logic := 'U';
          un7_noe32ri_0   : out   std_logic;
          un5_noe16ri_0   : out   std_logic;
          WDOGTO          : out   std_logic;
          HWRES_c_0_6     : in    std_logic := 'U';
          HWRES_c_0_5     : in    std_logic := 'U';
          HWRES_c_0_4     : in    std_logic := 'U';
          HWRES_c_0_3     : in    std_logic := 'U';
          HWRES_c_23_0    : in    std_logic := 'U';
          HWRES_c_21_0    : in    std_logic := 'U';
          HWRES_c_13_0    : in    std_logic := 'U';
          HWRES_c_0_0     : in    std_logic := 'U';
          NOEAD_c_0_0     : out   std_logic;
          HWRES_c_13      : in    std_logic := 'U';
          CLK_c_c         : in    std_logic := 'U';
          RUN_c_0_0       : out   std_logic;
          HWRES_c_0_6_0   : in    std_logic := 'U'
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CROM
    port( CROMWDT   : in    std_logic_vector(7 downto 0) := (others => 'U');
          RAMAD_VME : in    std_logic_vector(8 downto 0) := (others => 'U');
          CROMWAD   : in    std_logic_vector(8 downto 0) := (others => 'U');
          RAMDT     : out   std_logic_vector(7 downto 0);
          WRCROM    : in    std_logic := 'U';
          RAMRD     : in    std_logic := 'U';
          CLK_c_c   : in    std_logic := 'U'
        );
  end component;

  component RESET_MOD
    port( TICK_2_d0     : out   std_logic;
          TICK_1_d0     : out   std_logic;
          TICK_0_d0     : out   std_logic;
          LBSP_c        : out   std_logic_vector(2 to 2);
          PULSE         : in    std_logic_vector(1 to 1) := (others => 'U');
          LBSP_c_0      : out   std_logic_vector(2 to 2);
          LBSP_c_1      : out   std_logic_vector(2 to 2);
          TST_c         : out   std_logic_vector(15 downto 13);
          TICK_0_2      : out   std_logic;
          TICK_0_0      : out   std_logic;
          TICK_1        : out   std_logic_vector(0 to 0);
          TICK_2        : out   std_logic_vector(0 to 0);
          REG_464       : out   std_logic;
          REG_463       : out   std_logic;
          REG_462       : out   std_logic;
          REG_461       : out   std_logic;
          REG_460       : out   std_logic;
          REG_459       : out   std_logic;
          REG_458       : out   std_logic;
          REG_456       : out   std_logic;
          REG_455       : out   std_logic;
          REG_454       : out   std_logic;
          REG_453       : out   std_logic;
          REG_451       : out   std_logic;
          REG_457       : out   std_logic;
          REG_452       : out   std_logic;
          REG_449       : out   std_logic;
          REG_450       : out   std_logic;
          REG_0         : in    std_logic := 'U';
          PON_LOAD_i    : out   std_logic;
          EV_RES_c      : out   std_logic;
          RUN_c         : in    std_logic := 'U';
          LOAD_RES      : in    std_logic := 'U';
          CLEAR         : out   std_logic;
          BNCRES_c      : in    std_logic := 'U';
          EVRES_c       : in    std_logic := 'U';
          WDOGTO        : in    std_logic := 'U';
          HWRES_c       : out   std_logic;
          HWRES_c_i_0   : out   std_logic;
          CLEAR_i_0     : out   std_logic;
          RUN_c_0       : in    std_logic := 'U';
          ALICLK_c      : in    std_logic := 'U';
          HWRES_c_0     : out   std_logic;
          HWRES_c_1     : out   std_logic;
          HWRES_c_2     : out   std_logic;
          HWRES_c_3     : out   std_logic;
          HWRES_c_4     : out   std_logic;
          HWRES_c_5     : out   std_logic;
          NPWON_c       : in    std_logic := 'U';
          HWRES_c_6     : out   std_logic;
          HWRES_c_7     : out   std_logic;
          HWRES_c_8     : out   std_logic;
          HWRES_c_9     : out   std_logic;
          HWRES_c_10    : out   std_logic;
          HWRES_c_11    : out   std_logic;
          HWRES_c_12    : out   std_logic;
          HWRES_c_13    : out   std_logic;
          HWRES_c_14    : out   std_logic;
          HWRES_c_15    : out   std_logic;
          HWRES_c_16    : out   std_logic;
          HWRES_c_17    : out   std_logic;
          HWRES_c_18    : out   std_logic;
          HWRES_c_19    : out   std_logic;
          HWRES_c_20    : out   std_logic;
          HWRES_c_21    : out   std_logic;
          HWRES_c_22    : out   std_logic;
          HWRES_c_23    : out   std_logic;
          HWRES_c_24    : out   std_logic;
          HWRES_c_25    : out   std_logic;
          HWRES_c_26    : out   std_logic;
          HWRES_c_27    : out   std_logic;
          HWRES_c_28    : out   std_logic;
          HWRES_c_29    : out   std_logic;
          HWRES_c_30    : out   std_logic;
          HWRES_c_31    : out   std_logic;
          HWRES_c_32    : out   std_logic;
          HWRES_c_33    : out   std_logic;
          HWRES_c_34    : out   std_logic;
          HWRES_c_35    : out   std_logic;
          HWRES_c_36    : out   std_logic;
          CLEAR_0       : out   std_logic;
          CLEAR_2       : out   std_logic;
          CLEAR_3       : out   std_logic;
          CLEAR_4       : out   std_logic;
          CLEAR_5       : out   std_logic;
          CLEAR_6       : out   std_logic;
          CLEAR_7       : out   std_logic;
          CLEAR_8       : out   std_logic;
          LOAD_RES_2    : in    std_logic := 'U';
          CLEAR_9       : out   std_logic;
          CLEAR_10      : out   std_logic;
          CLEAR_11      : out   std_logic;
          CLEAR_12      : out   std_logic;
          CLEAR_13      : out   std_logic;
          CLEAR_14      : out   std_logic;
          CLEAR_15      : out   std_logic;
          CLEAR_16      : out   std_logic;
          CLEAR_17      : out   std_logic;
          CLEAR_18      : out   std_logic;
          LOAD_RES_1    : in    std_logic := 'U';
          CLEAR_19      : out   std_logic;
          CLEAR_20      : out   std_logic;
          CLEAR_21      : out   std_logic;
          CLEAR_22      : out   std_logic;
          CLEAR_23      : out   std_logic;
          CLEAR_24      : out   std_logic;
          CLEAR_25      : out   std_logic;
          CLEAR_26      : out   std_logic;
          CLEAR_27      : out   std_logic;
          LOAD_RES_0    : in    std_logic := 'U';
          CLEAR_28      : out   std_logic;
          HWRES_c_36_0  : out   std_logic;
          HWRES_c_32_0  : out   std_logic;
          NPWON_c_1     : in    std_logic := 'U';
          HWRES_c_23_0  : out   std_logic;
          HWRES_c_22_0  : out   std_logic;
          HWRES_c_21_0  : out   std_logic;
          HWRES_c_13_0  : out   std_logic;
          HWRES_c_10_0  : out   std_logic;
          HWRES_c_0_0   : out   std_logic;
          HWRES_c_0_2   : out   std_logic;
          HWRES_c_0_3   : out   std_logic;
          HWRES_c_0_4   : out   std_logic;
          HWRES_c_0_5   : out   std_logic;
          HWRES_c_0_6   : out   std_logic;
          RUN_c_0_0     : in    std_logic := 'U';
          NLBCLR_c      : out   std_logic;
          SYSRESB_c     : in    std_logic := 'U';
          CLK_c_c       : in    std_logic := 'U';
          NPWON_c_2     : in    std_logic := 'U';
          HWRES_c_27_0  : out   std_logic;
          NPWON_c_3     : in    std_logic := 'U';
          HWRES_c_7_0   : out   std_logic;
          NPWON_c_0     : in    std_logic := 'U';
          HWRES_c_0_6_0 : out   std_logic
        );
  end component;

  component SPI_INTERF
    port( CROMWDT        : out   std_logic_vector(7 downto 0);
          DACCFG_WDT     : out   std_logic_vector(13 downto 4);
          TICK           : in    std_logic_vector(1 to 1) := (others => 'U');
          FBOUT          : out   std_logic_vector(7 downto 0);
          REG_i_0        : in    std_logic_vector(80 to 80) := (others => 'U');
          REG_400        : out   std_logic;
          REG_398        : out   std_logic;
          REG_396        : out   std_logic;
          REG_393        : out   std_logic;
          REG_0          : in    std_logic := 'U';
          REG_1          : in    std_logic := 'U';
          REG_2          : in    std_logic := 'U';
          REG_3          : in    std_logic := 'U';
          REG_4          : in    std_logic := 'U';
          REG_5          : in    std_logic := 'U';
          REG_6          : in    std_logic := 'U';
          REG_7          : in    std_logic := 'U';
          REG_8          : in    std_logic := 'U';
          REG_399        : out   std_logic;
          REG_395        : out   std_logic;
          REG_397        : out   std_logic;
          REG_394        : out   std_logic;
          CROMWAD        : out   std_logic_vector(8 downto 0);
          sstate_0_2     : out   std_logic;
          PULSE_6        : in    std_logic := 'U';
          PULSE_0        : in    std_logic := 'U';
          PULSE_10       : in    std_logic := 'U';
          sstate_0_i_0   : in    std_logic_vector(2 to 2) := (others => 'U');
          HWRES_c_30     : in    std_logic := 'U';
          HWRES_c_23_0   : in    std_logic := 'U';
          HWRES_c_28     : in    std_logic := 'U';
          HWRES_c_31     : in    std_logic := 'U';
          HWRES_c_24     : in    std_logic := 'U';
          HWRES_c_25     : in    std_logic := 'U';
          DACCFG_nWR     : out   std_logic;
          PDLCFG_nWR     : out   std_logic;
          HWRES_c_32     : in    std_logic := 'U';
          WRCROM         : out   std_logic;
          HWRES_c_26     : in    std_logic := 'U';
          HWRES_c_27     : in    std_logic := 'U';
          NCYC_RELOAD_in : in    std_logic := 'U';
          HWRES_c_29     : in    std_logic := 'U';
          un1_drive_spi  : out   std_logic;
          F_SO_c         : in    std_logic := 'U';
          LOAD_RES       : out   std_logic;
          DRIVE_RELOAD   : out   std_logic;
          ISCK           : out   std_logic;
          FWIMG2LOAD     : in    std_logic := 'U';
          ISI            : out   std_logic;
          FCS_c          : out   std_logic;
          PON_LOAD_i     : in    std_logic := 'U';
          HWRES_c_32_0   : in    std_logic := 'U';
          LOAD_RES_0     : out   std_logic;
          LOAD_RES_1     : out   std_logic;
          LOAD_RES_2     : out   std_logic;
          CLK_c_c        : in    std_logic := 'U';
          HWRES_c_27_0   : in    std_logic := 'U';
          LOAD_RES_3     : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ROC32
    port( DPR          : out   std_logic_vector(31 downto 0);
          un2_evread_0 : out   std_logic;
          CHANNEL      : out   std_logic_vector(2 downto 0);
          CHIP_ADDR    : out   std_logic_vector(2 downto 0);
          I2C_RDATA    : in    std_logic_vector(9 downto 0) := (others => 'U');
          OR_RDATA     : in    std_logic_vector(9 downto 0) := (others => 'U');
          PDL_RDATA    : in    std_logic_vector(7 downto 0) := (others => 'U');
          GA_c         : in    std_logic_vector(3 downto 0) := (others => 'U');
          OR_RADDR     : out   std_logic_vector(5 downto 0);
          PDL_RADDR    : out   std_logic_vector(5 downto 0);
          LBSP_c       : in    std_logic_vector(2 to 2) := (others => 'U');
          LBSP_c_1     : in    std_logic_vector(2 to 2) := (others => 'U');
          LBSP_c_0     : in    std_logic_vector(2 to 2) := (others => 'U');
          PULSE        : in    std_logic_vector(3 downto 2) := (others => 'U');
          REG_i_0      : in    std_logic_vector(5 to 5) := (others => 'U');
          REG_c        : in    std_logic_vector(23 downto 21) := (others => 'U');
          REG_330      : out   std_logic;
          REG_329      : out   std_logic;
          REG_328      : out   std_logic;
          REG_408      : in    std_logic := 'U';
          REG_410      : in    std_logic := 'U';
          REG_432      : in    std_logic := 'U';
          REG_415      : in    std_logic := 'U';
          REG_406      : in    std_logic := 'U';
          REG_418      : in    std_logic := 'U';
          REG_421      : in    std_logic := 'U';
          REG_430      : in    std_logic := 'U';
          REG_433      : in    std_logic := 'U';
          REG_424      : in    std_logic := 'U';
          REG_427      : in    std_logic := 'U';
          REG_416      : in    std_logic := 'U';
          REG_419      : in    std_logic := 'U';
          REG_412      : in    std_logic := 'U';
          REG_413      : in    std_logic := 'U';
          REG_428      : in    std_logic := 'U';
          REG_431      : in    std_logic := 'U';
          REG_422      : in    std_logic := 'U';
          REG_425      : in    std_logic := 'U';
          REG_414      : in    std_logic := 'U';
          REG_417      : in    std_logic := 'U';
          REG_409      : in    std_logic := 'U';
          REG_411      : in    std_logic := 'U';
          REG_426      : in    std_logic := 'U';
          REG_429      : in    std_logic := 'U';
          REG_420      : in    std_logic := 'U';
          REG_423      : in    std_logic := 'U';
          REG_407      : in    std_logic := 'U';
          REG_434      : in    std_logic := 'U';
          REG_435      : in    std_logic := 'U';
          REG_404      : in    std_logic := 'U';
          REG_405      : in    std_logic := 'U';
          REG_43       : in    std_logic := 'U';
          REG_44       : in    std_logic := 'U';
          REG_45       : in    std_logic := 'U';
          REG_46       : in    std_logic := 'U';
          REG_47       : in    std_logic := 'U';
          REG_48       : in    std_logic := 'U';
          REG_49       : in    std_logic := 'U';
          REG_50       : in    std_logic := 'U';
          REG_51       : in    std_logic := 'U';
          REG_52       : in    std_logic := 'U';
          REG_53       : in    std_logic := 'U';
          REG_54       : in    std_logic := 'U';
          REG_55       : in    std_logic := 'U';
          REG_56       : in    std_logic := 'U';
          REG_57       : in    std_logic := 'U';
          REG_58       : in    std_logic := 'U';
          REG_59       : in    std_logic := 'U';
          REG_60       : in    std_logic := 'U';
          REG_61       : in    std_logic := 'U';
          REG_62       : in    std_logic := 'U';
          REG_63       : in    std_logic := 'U';
          REG_64       : in    std_logic := 'U';
          REG_65       : in    std_logic := 'U';
          REG_66       : in    std_logic := 'U';
          REG_67       : in    std_logic := 'U';
          REG_68       : in    std_logic := 'U';
          REG_69       : in    std_logic := 'U';
          REG_70       : in    std_logic := 'U';
          REG_71       : in    std_logic := 'U';
          REG_72       : in    std_logic := 'U';
          REG_73       : in    std_logic := 'U';
          REG_74       : in    std_logic := 'U';
          REG_41       : out   std_logic;
          REG_42       : out   std_logic;
          REG_0        : in    std_logic := 'U';
          REG_15       : out   std_logic;
          REG_27       : out   std_logic;
          REG_28       : out   std_logic;
          REG_30       : out   std_logic;
          REG_29       : out   std_logic;
          REG_39       : out   std_logic;
          REG_37       : out   std_logic;
          REG_36       : out   std_logic;
          REG_34       : out   std_logic;
          REG_33       : out   std_logic;
          REG_38       : out   std_logic;
          REG_35       : out   std_logic;
          REG_40       : out   std_logic;
          REG_31       : out   std_logic;
          REG_32       : out   std_logic;
          EF           : out   std_logic;
          FF_c         : out   std_logic;
          NRDMEB       : in    std_logic := 'U';
          CLEAR_i_0    : in    std_logic := 'U';
          CLEAR_14     : in    std_logic := 'U';
          CLEAR_13     : in    std_logic := 'U';
          CLEAR_4      : in    std_logic := 'U';
          CLEAR_3      : in    std_logic := 'U';
          CLEAR_2      : in    std_logic := 'U';
          CLEAR_8      : in    std_logic := 'U';
          CLEAR_7      : in    std_logic := 'U';
          CLEAR_6      : in    std_logic := 'U';
          CLEAR_11     : in    std_logic := 'U';
          CLEAR_10     : in    std_logic := 'U';
          CLEAR_19     : in    std_logic := 'U';
          CLEAR_9      : in    std_logic := 'U';
          CLEAR_18     : in    std_logic := 'U';
          CLEAR_12     : in    std_logic := 'U';
          CLEAR_15     : in    std_logic := 'U';
          CLEAR_20     : in    std_logic := 'U';
          CLEAR_5      : in    std_logic := 'U';
          PDL_RACK     : in    std_logic := 'U';
          CLEAR_17     : in    std_logic := 'U';
          OR_RACK      : in    std_logic := 'U';
          CLEAR_16     : in    std_logic := 'U';
          L2R_c_c      : in    std_logic := 'U';
          L2A_c_c      : in    std_logic := 'U';
          HWRES_c_12   : in    std_logic := 'U';
          L1A_c_c      : in    std_logic := 'U';
          ALICLK_c     : in    std_logic := 'U';
          HWRES_c_11   : in    std_logic := 'U';
          DTEST_FIFO   : out   std_logic;
          I2C_CHAIN    : out   std_logic;
          PDL_RREQ     : out   std_logic;
          I2C_RREQ     : out   std_logic;
          EVRDY_c      : out   std_logic;
          OR_RREQ      : out   std_logic;
          I2C_RACK     : in    std_logic := 'U';
          EVNT_TRG     : out   std_logic;
          EVREAD       : in    std_logic := 'U';
          CLK_c_c      : in    std_logic := 'U';
          CLEAR_0      : in    std_logic := 'U';
          I_8          : in    std_logic := 'U';
          I_16         : in    std_logic := 'U'
        );
  end component;

  component I2C_INTERF
    port( PULSE         : in    std_logic_vector(7 to 7) := (others => 'U');
          I2C_RDATA     : out   std_logic_vector(9 downto 0);
          CHIP_ADDR     : in    std_logic_vector(2 downto 0) := (others => 'U');
          CHANNEL       : in    std_logic_vector(2 downto 0) := (others => 'U');
          TICK          : in    std_logic_vector(0 to 0) := (others => 'U');
          TICK_2        : in    std_logic_vector(0 to 0) := (others => 'U');
          REG_107       : out   std_logic;
          REG_108       : out   std_logic;
          REG_109       : out   std_logic;
          REG_110       : out   std_logic;
          REG_111       : out   std_logic;
          REG_112       : out   std_logic;
          REG_113       : out   std_logic;
          REG_114       : out   std_logic;
          REG_0         : in    std_logic := 'U';
          REG_84        : in    std_logic := 'U';
          REG_85        : in    std_logic := 'U';
          REG_91        : in    std_logic := 'U';
          REG_92        : in    std_logic := 'U';
          REG_99        : out   std_logic;
          REG_93        : in    std_logic := 'U';
          REG_94        : in    std_logic := 'U';
          REG_95        : in    std_logic := 'U';
          REG_96        : in    std_logic := 'U';
          REG_97        : in    std_logic := 'U';
          REG_98        : in    std_logic := 'U';
          REG_83        : in    std_logic := 'U';
          REG_100       : out   std_logic;
          TICK_1        : in    std_logic_vector(0 to 0) := (others => 'U');
          TICK_0        : in    std_logic_vector(0 to 0) := (others => 'U');
          HWRES_c_4     : in    std_logic := 'U';
          HWRES_c_7     : in    std_logic := 'U';
          HWRES_c_11    : in    std_logic := 'U';
          HWRES_c_10    : in    std_logic := 'U';
          HWRES_c_5     : in    std_logic := 'U';
          HWRES_c_3     : in    std_logic := 'U';
          HWRES_c_6     : in    std_logic := 'U';
          I2C_RACK      : out   std_logic;
          SDAout_del2   : out   std_logic;
          HWRES_c_9     : in    std_logic := 'U';
          HWRES_c_8     : in    std_logic := 'U';
          un1_sdaa_0_a3 : out   std_logic;
          RUN_c_0_0     : in    std_logic := 'U';
          RUN_c_0       : in    std_logic := 'U';
          I2C_CHAIN     : in    std_logic := 'U';
          I2C_RREQ      : in    std_logic := 'U';
          SDA1_in       : in    std_logic := 'U';
          SDA0_in       : in    std_logic := 'U';
          un1_sdab_i    : out   std_logic;
          SCLB_i_a3     : out   std_logic;
          SCLA_i_a3     : out   std_logic;
          HWRES_c_10_0  : in    std_logic := 'U';
          CLK_c_c       : in    std_logic := 'U';
          HWRES_c_7_0   : in    std_logic := 'U'
        );
  end component;

  component ctrl
    port( TST_c_c      : in    std_logic_vector(3 to 3) := (others => 'U');
          PULSE        : in    std_logic_vector(2 to 2) := (others => 'U');
          TICK_0       : in    std_logic_vector(2 to 2) := (others => 'U');
          REG_15       : in    std_logic := 'U';
          REG_0        : in    std_logic := 'U';
          REG_1        : in    std_logic := 'U';
          REG_2        : in    std_logic := 'U';
          REG_3        : in    std_logic := 'U';
          REG_4        : in    std_logic := 'U';
          REG_5        : in    std_logic := 'U';
          TICK         : in    std_logic_vector(2 to 2) := (others => 'U');
          nLBRDY_c     : in    std_logic := 'U';
          EVNT_TRG     : in    std_logic := 'U';
          HWRES_c_32_0 : in    std_logic := 'U';
          RUN_c        : in    std_logic := 'U';
          HWRES_c_34   : in    std_logic := 'U';
          CLK_c_c      : in    std_logic := 'U';
          HWRES_c_33   : in    std_logic := 'U';
          N_18         : out   std_logic;
          N_20         : out   std_logic;
          N_22         : out   std_logic;
          N_24         : out   std_logic;
          N_26         : out   std_logic;
          N_28         : out   std_logic
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component DAC_INTERF
    port( TICK_0        : in    std_logic_vector(2 to 2) := (others => 'U');
          SYNC_c        : out   std_logic_vector(15 downto 0);
          DACCFG_DT     : in    std_logic_vector(15 downto 0) := (others => 'U');
          REG           : in    std_logic_vector(264 downto 233) := (others => 'U');
          PULSE         : in    std_logic_vector(9 to 9) := (others => 'U');
          DACCFG_RAD    : out   std_logic_vector(3 downto 0);
          HWRES_c_36    : in    std_logic := 'U';
          HWRES_c_34    : in    std_logic := 'U';
          HWRES_c_35    : in    std_logic := 'U';
          RUN_c_0       : in    std_logic := 'U';
          DACCFG_nRD    : out   std_logic;
          SCLK_DAC_c    : out   std_logic;
          SDIN_DAC_c    : out   std_logic;
          HWRES_c_0     : in    std_logic := 'U';
          HWRES_c_3     : in    std_logic := 'U';
          HWRES_c_0_6_0 : in    std_logic := 'U';
          HWRES_c_2     : in    std_logic := 'U';
          HWRES_c_1     : in    std_logic := 'U';
          HWRES_c_36_0  : in    std_logic := 'U';
          CLK_c_c       : in    std_logic := 'U';
          HWRES_c       : in    std_logic := 'U'
        );
  end component;

  component DACCFG
    port( DACCFG_WDT : in    std_logic_vector(13 downto 4) := (others => 'U');
          DACCFG_RAD : in    std_logic_vector(3 downto 0) := (others => 'U');
          DACCFG_DT  : out   std_logic_vector(15 downto 0);
          CROMWAD    : in    std_logic_vector(4 downto 1) := (others => 'U');
          DACCFG_nRD : in    std_logic := 'U';
          DACCFG_nWR : in    std_logic := 'U';
          CLK_c_c    : in    std_logic := 'U'
        );
  end component;

    signal \PULSE[0]\, \PULSE[1]\, \PULSE[2]\, \PULSE[3]\, 
        \PULSE[6]\, \PULSE[7]\, \PULSE[8]\, \PULSE[9]\, 
        \PULSE[10]\, \TICK[0]\, \TICK[1]\, \TICK[2]\, \RAMDT[0]\, 
        \RAMDT[1]\, \RAMDT[2]\, \RAMDT[3]\, \RAMDT[4]\, 
        \RAMDT[5]\, \RAMDT[6]\, \RAMDT[7]\, \CROMWDT[0]\, 
        \CROMWDT[1]\, \CROMWDT[2]\, \CROMWDT[3]\, \CROMWDT[4]\, 
        \CROMWDT[5]\, \CROMWDT[6]\, \CROMWDT[7]\, WRCROM, RAMRD, 
        \CROMWAD[0]\, \CROMWAD[1]\, \CROMWAD[2]\, \CROMWAD[3]\, 
        \CROMWAD[4]\, \CROMWAD[5]\, \CROMWAD[6]\, \CROMWAD[7]\, 
        \CROMWAD[8]\, \RAMAD_VME[0]\, \RAMAD_VME[1]\, 
        \RAMAD_VME[2]\, \RAMAD_VME[3]\, \RAMAD_VME[4]\, 
        \RAMAD_VME[5]\, \RAMAD_VME[6]\, \RAMAD_VME[7]\, 
        \RAMAD_VME[8]\, \DACCFG_DT[0]\, \DACCFG_DT[1]\, 
        \DACCFG_DT[2]\, \DACCFG_DT[3]\, \DACCFG_DT[4]\, 
        \DACCFG_DT[5]\, \DACCFG_DT[6]\, \DACCFG_DT[7]\, 
        \DACCFG_DT[8]\, \DACCFG_DT[9]\, \DACCFG_DT[10]\, 
        \DACCFG_DT[11]\, \DACCFG_DT[12]\, \DACCFG_DT[13]\, 
        \DACCFG_DT[14]\, \DACCFG_DT[15]\, \DACCFG_WDT[4]\, 
        \DACCFG_WDT[5]\, \DACCFG_WDT[6]\, \DACCFG_WDT[7]\, 
        \DACCFG_WDT[8]\, \DACCFG_WDT[9]\, \DACCFG_WDT[10]\, 
        \DACCFG_WDT[11]\, \DACCFG_WDT[12]\, \DACCFG_WDT[13]\, 
        DACCFG_nWR, DACCFG_nRD, \DACCFG_RAD[0]\, \DACCFG_RAD[1]\, 
        \DACCFG_RAD[2]\, \DACCFG_RAD[3]\, \I2C_RDATA[0]\, 
        \I2C_RDATA[1]\, \I2C_RDATA[2]\, \I2C_RDATA[3]\, 
        \I2C_RDATA[4]\, \I2C_RDATA[5]\, \I2C_RDATA[6]\, 
        \I2C_RDATA[7]\, \I2C_RDATA[8]\, \I2C_RDATA[9]\, I2C_RREQ, 
        I2C_RACK, I2C_CHAIN, \CHIP_ADDR[0]\, \CHIP_ADDR[1]\, 
        \CHIP_ADDR[2]\, \CHANNEL[0]\, \CHANNEL[1]\, \CHANNEL[2]\, 
        \PDLCFG_DT[0]\, \PDLCFG_DT[1]\, \PDLCFG_DT[2]\, 
        \PDLCFG_DT[3]\, \PDLCFG_DT[4]\, \PDLCFG_DT[5]\, 
        \PDLCFG_DT[6]\, \PDLCFG_DT[7]\, PDLCFG_nWR, PDLCFG_nRD, 
        \PDLCFG_RAD[0]\, \PDLCFG_RAD[1]\, \PDLCFG_RAD[2]\, 
        \PDLCFG_RAD[3]\, \PDLCFG_RAD[4]\, \PDLCFG_RAD[5]\, 
        LOAD_RES, WDOGTO, CLEAR, \PDL_RDATA[0]\, \PDL_RDATA[1]\, 
        \PDL_RDATA[2]\, \PDL_RDATA[3]\, \PDL_RDATA[4]\, 
        \PDL_RDATA[5]\, \PDL_RDATA[6]\, \PDL_RDATA[7]\, 
        \PDL_RADDR[0]\, \PDL_RADDR[1]\, \PDL_RADDR[2]\, 
        \PDL_RADDR[3]\, \PDL_RADDR[4]\, \PDL_RADDR[5]\, PDL_RREQ, 
        PDL_RACK, \OR_RDATA[0]\, \OR_RDATA[1]\, \OR_RDATA[2]\, 
        \OR_RDATA[3]\, \OR_RDATA[4]\, \OR_RDATA[5]\, 
        \OR_RDATA[6]\, \OR_RDATA[7]\, \OR_RDATA[8]\, 
        \OR_RDATA[9]\, \OR_RADDR[0]\, \OR_RADDR[1]\, 
        \OR_RADDR[2]\, \OR_RADDR[3]\, \OR_RADDR[4]\, 
        \OR_RADDR[5]\, OR_RREQ, OR_RACK, \DPR[0]\, \DPR[1]\, 
        \DPR[2]\, \DPR[3]\, \DPR[4]\, \DPR[5]\, \DPR[6]\, 
        \DPR[7]\, \DPR[8]\, \DPR[9]\, \DPR[10]\, \DPR[11]\, 
        \DPR[12]\, \DPR[13]\, \DPR[14]\, \DPR[15]\, \DPR[16]\, 
        \DPR[17]\, \DPR[18]\, \DPR[19]\, \DPR[20]\, \DPR[21]\, 
        \DPR[22]\, \DPR[23]\, \DPR[24]\, \DPR[25]\, \DPR[26]\, 
        \DPR[27]\, \DPR[28]\, \DPR[29]\, \DPR[30]\, \DPR[31]\, 
        NRDMEB, EF, EVREAD, DTEST_FIFO, \FBOUT[0]\, \FBOUT[1]\, 
        \FBOUT[2]\, \FBOUT[3]\, \FBOUT[4]\, \FBOUT[5]\, 
        \FBOUT[6]\, \FBOUT[7]\, FWIMG2LOAD, \REG[5]\, \REG[6]\, 
        \REG[8]\, \REG[17]\, \REG[20]\, \REG[32]\, \REG[33]\, 
        \REG[34]\, \REG[35]\, \REG[36]\, \REG[37]\, \REG[38]\, 
        \REG[39]\, \REG[40]\, \REG[41]\, \REG[42]\, \REG[43]\, 
        \REG[44]\, \REG[45]\, \REG[46]\, \REG[47]\, \REG[48]\, 
        \REG[49]\, \REG[50]\, \REG[51]\, \REG[52]\, \REG[53]\, 
        \REG[54]\, \REG[55]\, \REG[56]\, \REG[57]\, \REG[58]\, 
        \REG[59]\, \REG[60]\, \REG[61]\, \REG[62]\, \REG[63]\, 
        \REG[64]\, \REG[65]\, \REG[66]\, \REG[67]\, \REG[68]\, 
        \REG[69]\, \REG[70]\, \REG[71]\, \REG[72]\, \REG[73]\, 
        \REG[74]\, \REG[75]\, \REG[76]\, \REG[77]\, \REG[78]\, 
        \REG[79]\, \REG[80]\, \REG[81]\, \REG[82]\, \REG[83]\, 
        \REG[84]\, \REG[85]\, \REG[86]\, \REG[87]\, \REG[88]\, 
        \REG[89]\, \REG[90]\, \REG[91]\, \REG[97]\, \REG[98]\, 
        \REG[99]\, \REG[100]\, \REG[101]\, \REG[102]\, \REG[103]\, 
        \REG[104]\, \REG[105]\, \REG[106]\, \REG[113]\, 
        \REG[114]\, \REG[115]\, \REG[116]\, \REG[117]\, 
        \REG[118]\, \REG[119]\, \REG[120]\, \REG[121]\, 
        \REG[122]\, \REG[123]\, \REG[124]\, \REG[125]\, 
        \REG[126]\, \REG[127]\, \REG[129]\, \REG[130]\, 
        \REG[131]\, \REG[132]\, \REG[133]\, \REG[134]\, 
        \REG[135]\, \REG[136]\, \REG[137]\, \REG[138]\, 
        \REG[139]\, \REG[140]\, \REG[141]\, \REG[142]\, 
        \REG[143]\, \REG[144]\, \REG[145]\, \REG[153]\, 
        \REG[154]\, \REG[155]\, \REG[156]\, \REG[157]\, 
        \REG[158]\, \REG[159]\, \REG[160]\, \REG[161]\, 
        \REG[162]\, \REG[163]\, \REG[164]\, \REG[165]\, 
        \REG[166]\, \REG[167]\, \REG[168]\, \REG[169]\, 
        \REG[170]\, \REG[171]\, \REG[172]\, \REG[173]\, 
        \REG[174]\, \REG[175]\, \REG[176]\, \REG[177]\, 
        \REG[178]\, \REG[179]\, \REG[180]\, \REG[181]\, 
        \REG[182]\, \REG[183]\, \REG[184]\, \REG[185]\, 
        \REG[186]\, \REG[187]\, \REG[188]\, \REG[189]\, 
        \REG[190]\, \REG[191]\, \REG[192]\, \REG[193]\, 
        \REG[194]\, \REG[195]\, \REG[196]\, \REG[197]\, 
        \REG[198]\, \REG[199]\, \REG[200]\, \REG[233]\, 
        \REG[234]\, \REG[235]\, \REG[236]\, \REG[237]\, 
        \REG[238]\, \REG[239]\, \REG[240]\, \REG[241]\, 
        \REG[242]\, \REG[243]\, \REG[244]\, \REG[245]\, 
        \REG[246]\, \REG[247]\, \REG[248]\, \REG[249]\, 
        \REG[250]\, \REG[251]\, \REG[252]\, \REG[253]\, 
        \REG[254]\, \REG[255]\, \REG[256]\, \REG[257]\, 
        \REG[258]\, \REG[259]\, \REG[260]\, \REG[261]\, 
        \REG[262]\, \REG[263]\, \REG[264]\, \REG[333]\, 
        \REG[334]\, \REG[335]\, \REG[345]\, \REG[346]\, 
        \REG[360]\, \REG[361]\, \REG[362]\, \REG[363]\, 
        \REG[364]\, \REG[365]\, \REG[366]\, \REG[367]\, 
        \REG[368]\, \REG[369]\, \REG[370]\, \REG[371]\, 
        \REG[372]\, \REG[373]\, \REG[374]\, \REG[375]\, 
        \REG[376]\, \REG[377]\, \REG[378]\, \REG[379]\, 
        \REG[380]\, \REG[381]\, \REG[382]\, \REG[383]\, 
        \REG[384]\, \REG[409]\, \REG[410]\, \REG[411]\, 
        \REG[412]\, \REG[413]\, \REG[414]\, \REG[415]\, 
        \REG[416]\, \REG[417]\, \REG[418]\, \REG[419]\, 
        \REG[420]\, \REG[421]\, \REG[422]\, \REG[423]\, 
        \REG[424]\, \REG[425]\, \REG[426]\, \REG[427]\, 
        \REG[428]\, \REG[429]\, \REG[430]\, \REG[431]\, 
        \REG[432]\, \REG[433]\, \REG[434]\, \REG[435]\, 
        \REG[436]\, \REG[437]\, \REG[438]\, \REG[439]\, 
        \REG[440]\, \REG[441]\, \REG[442]\, \REG[443]\, 
        \REG[444]\, \REG[445]\, \REG[446]\, \REG[456]\, 
        \REG[457]\, \REG[458]\, \REG[459]\, \REG[460]\, 
        \REG[461]\, \REG[462]\, \REG[463]\, \REG[464]\, 
        \REG[465]\, \REG[466]\, \REG[467]\, \REG[468]\, 
        \REG[469]\, \REG[470]\, \REG[471]\, \REG[472]\, 
        \REG[473]\, \REG[474]\, \REG[475]\, \REG[476]\, 
        \REG[477]\, \REG[478]\, \REG[479]\, \REG[480]\, 
        \REG[481]\, N_18, N_20, N_22, N_24, N_26, N_28, 
        \I3.P0[0]\, \I3.P0[1]\, \I3.P0[2]\, \I3.P0[3]\, 
        \I3.P0[4]\, \I3.P0[5]\, \I3.P0[6]\, \I3.P0[7]\, 
        \I3.P0[8]\, \I3.P0[9]\, \I3.P0[10]\, \I3.P0[11]\, 
        \I3.P0[12]\, \I3.P0[13]\, \I3.P0[14]\, \I3.P0[15]\, 
        \I3.P0[16]\, \I3.P0[17]\, \I3.P0[18]\, \I3.P0[19]\, 
        \I3.P0[20]\, \I3.P0[21]\, \I3.P0[22]\, \I3.P0[23]\, 
        \I3.P0[24]\, \I3.P0[25]\, \I3.P0[26]\, \I3.P0[27]\, 
        \I3.P0[28]\, \I3.P0[29]\, \I3.P0[30]\, \I3.P0[31]\, 
        \I3.P0[32]\, \I3.P0[33]\, \I3.P0[34]\, \I3.P0[35]\, 
        \I3.P0[36]\, \I3.P0[37]\, \I3.P0[38]\, \I3.P0[39]\, 
        \I3.P0[40]\, \I3.P0[41]\, \I3.P0[42]\, \I3.P0[43]\, 
        \I3.P0[44]\, \I3.P0[45]\, \I3.P0[46]\, \I3.P0[47]\, 
        \I2.LB_nOE\, \I2.LB_i[0]\, \I2.LB_i[1]\, \I2.LB_i[2]\, 
        \I2.LB_i[3]\, \I2.LB_i[4]\, \I2.LB_i[5]\, \I2.LB_i[6]\, 
        \I2.LB_i[7]\, \I2.LB_i[8]\, \I2.LB_i[9]\, \I2.LB_i[10]\, 
        \I2.LB_i[11]\, \I2.LB_i[12]\, \I2.LB_i[13]\, 
        \I2.LB_i[14]\, \I2.LB_i[15]\, \I2.LB_i[16]\, 
        \I2.LB_i[17]\, \I2.LB_i[18]\, \I2.LB_i[19]\, 
        \I2.LB_i[20]\, \I2.LB_i[21]\, \I2.LB_i[22]\, 
        \I2.LB_i[23]\, \I2.LB_i[24]\, \I2.LB_i[25]\, 
        \I2.LB_i[26]\, \I2.LB_i[27]\, \I2.LB_i[28]\, 
        \I2.LB_i[29]\, \I2.LB_i[30]\, \I2.LB_i[31]\, 
        \I2.REGMAP[31]\, \I2.VADm[0]\, \I2.VADm[1]\, \I2.VADm[2]\, 
        \I2.VADm[3]\, \I2.VADm[4]\, \I2.VADm[5]\, \I2.VADm[6]\, 
        \I2.VADm[7]\, \I2.VADm[8]\, \I2.VADm[9]\, \I2.VADm[10]\, 
        \I2.VADm[11]\, \I2.VADm[12]\, \I2.VADm[13]\, 
        \I2.VADm[14]\, \I2.VADm[15]\, \I2.VADm[16]\, 
        \I2.VADm[17]\, \I2.VADm[18]\, \I2.VADm[19]\, 
        \I2.VADm[20]\, \I2.VADm[21]\, \I2.VADm[22]\, 
        \I2.VADm[23]\, \I2.VADm[24]\, \I2.VADm[25]\, 
        \I2.VADm[26]\, \I2.VADm[27]\, \I2.VADm[28]\, 
        \I2.VADm[29]\, \I2.VADm[30]\, \I2.VADm[31]\, 
        \I2.REGMAP[35]\, un5_noe16ri_0_0, un7_noe32ri_0_0, 
        \I2.VDBm[0]\, \I2.VDBm[1]\, \I2.VDBm[2]\, \I2.VDBm[3]\, 
        \I2.VDBm[4]\, \I2.VDBm[5]\, \I2.VDBm[6]\, \I2.VDBm[7]\, 
        \I2.VDBm[8]\, \I2.VDBm[9]\, \I2.VDBm[10]\, \I2.VDBm[12]\, 
        \I2.VDBm[13]\, \I2.VDBm[14]\, \I2.VDBm[15]\, 
        \I2.VDBm[16]\, \I2.VDBm[17]\, \I2.VDBm[18]\, 
        \I2.VDBm[19]\, \I2.VDBm[20]\, \I2.VDBm[22]\, 
        \I2.VDBm[23]\, \I2.VDBm[24]\, \I2.VDBm[25]\, 
        \I2.VDBm[26]\, \I2.VDBm[27]\, \I2.VDBm[28]\, 
        \I2.VDBm[29]\, \I2.VDBm[30]\, \I2.VDBm[31]\, 
        \VDBm_i_m2[11]\, \I2.N_500\, un1_drive_spi, 
        \I5.DRIVE_RELOAD\, \I5.ISCK\, \I5.ISI\, \I10.EVNT_TRG\, 
        \I1.SDAout_del2\, un1_sdaa_0_a3, un1_sdab_i, SCLB_i_a3, 
        SCLA_i_a3, ALICLK_c, \AMB_c[0]\, \AMB_c[1]\, \AMB_c[2]\, 
        \AMB_c[3]\, \AMB_c[4]\, \AMB_c[5]\, ASB_c, BNCRES_c, 
        DS0B_c, DS1B_c, EVRES_c, F_SO_c, \GA_c[0]\, \GA_c[1]\, 
        \GA_c[2]\, \GA_c[3]\, IACKB_c, NPWON_c, \REG_c[21]\, 
        \REG_c[22]\, \REG_c[23]\, SYSRESB_c, WRITEB_c, nLBRDY_c, 
        \AE_PDL_c[0]\, \AE_PDL_c[1]\, \AE_PDL_c[2]\, 
        \AE_PDL_c[3]\, \AE_PDL_c[4]\, \AE_PDL_c[5]\, 
        \AE_PDL_c[6]\, \AE_PDL_c[7]\, \AE_PDL_c[8]\, 
        \AE_PDL_c[9]\, \AE_PDL_c[10]\, \AE_PDL_c[11]\, 
        \AE_PDL_c[12]\, \AE_PDL_c[13]\, \AE_PDL_c[14]\, 
        \AE_PDL_c[15]\, \AE_PDL_c[16]\, \AE_PDL_c[17]\, 
        \AE_PDL_c[18]\, \AE_PDL_c[19]\, \AE_PDL_c[20]\, 
        \AE_PDL_c[21]\, \AE_PDL_c[22]\, \AE_PDL_c[23]\, 
        \AE_PDL_c[24]\, \AE_PDL_c[25]\, \AE_PDL_c[26]\, 
        \AE_PDL_c[27]\, \AE_PDL_c[28]\, \AE_PDL_c[29]\, 
        \AE_PDL_c[30]\, \AE_PDL_c[31]\, \AE_PDL_c[32]\, 
        \AE_PDL_c[33]\, \AE_PDL_c[34]\, \AE_PDL_c[35]\, 
        \AE_PDL_c[36]\, \AE_PDL_c[37]\, \AE_PDL_c[38]\, 
        \AE_PDL_c[39]\, \AE_PDL_c[40]\, \AE_PDL_c[41]\, 
        \AE_PDL_c[42]\, \AE_PDL_c[43]\, \AE_PDL_c[44]\, 
        \AE_PDL_c[45]\, \AE_PDL_c[46]\, \AE_PDL_c[47]\, CLK_c_c, 
        FCS_c, EVRDY_c, MD_PDL_c, MYBERR_c, NDTKIN_c, NLBCLR_c, 
        NLBRD_c, HWRES_c, \VCC\, NOE16W_c, NOE32W_c, NOEAD_c, 
        NSELCLK_c, \GND\, \P_PDL_c[1]\, \P_PDL_c[2]\, 
        \P_PDL_c[3]\, \P_PDL_c[4]\, \P_PDL_c[5]\, \P_PDL_c[6]\, 
        \P_PDL_c[7]\, SCLK_DAC_c, SCLK_PDL_c, SDIN_DAC_c, 
        SI_PDL_c, \SYNC_c[0]\, \SYNC_c[1]\, \SYNC_c[2]\, 
        \SYNC_c[3]\, \SYNC_c[4]\, \SYNC_c[5]\, \SYNC_c[6]\, 
        \SYNC_c[7]\, \SYNC_c[8]\, \SYNC_c[9]\, \SYNC_c[10]\, 
        \SYNC_c[11]\, \SYNC_c[12]\, \SYNC_c[13]\, \SYNC_c[14]\, 
        \SYNC_c[15]\, \TST_c[0]\, \TST_c[1]\, \TST_c[2]\, 
        \TST_c_c[3]\, \TST_c[4]\, \TST_c[5]\, \TST_c[13]\, 
        \TST_c[14]\, \TST_c[15]\, nLBAS_c, \LB_in[0]\, \LB_in[1]\, 
        \LB_in[2]\, \LB_in[3]\, \LB_in[4]\, \LB_in[5]\, 
        \LB_in[6]\, \LB_in[7]\, \LB_in[8]\, \LB_in[9]\, 
        \LB_in[10]\, \LB_in[11]\, \LB_in[12]\, \LB_in[13]\, 
        \LB_in[14]\, \LB_in[15]\, \LB_in[16]\, \LB_in[17]\, 
        \LB_in[18]\, \LB_in[19]\, \LB_in[20]\, \LB_in[21]\, 
        \LB_in[22]\, \LB_in[23]\, \LB_in[24]\, \LB_in[25]\, 
        \LB_in[26]\, \LB_in[27]\, \LB_in[28]\, \LB_in[29]\, 
        \LB_in[30]\, \LB_in[31]\, \LBSP_in[0]\, \LBSP_in[1]\, 
        \LBSP_c[2]\, EV_RES_c, L0_c_c, L1A_c_c, L1R_c_c, L2A_c_c, 
        L2R_c_c, RUN_c, LOS_c_c, SPULSE0_c_c, SPULSE1_c_c, 
        SPULSE2_c_c, \REG_c[0]\, \LBSP_in[15]\, \LBSP_in[16]\, 
        \LBSP_in[17]\, \LBSP_in[18]\, \LBSP_in[19]\, 
        \LBSP_in[20]\, \LBSP_in[21]\, \LBSP_in[22]\, 
        \LBSP_in[23]\, \LBSP_in[24]\, \LBSP_in[25]\, 
        \LBSP_in[26]\, \LBSP_in[27]\, \LBSP_in[28]\, 
        \LBSP_in[29]\, \LBSP_in[30]\, \LBSP_in[31]\, LWORDB_in, 
        NCYC_RELOAD_in, NLBLAST_c, SDA0_in, SDA1_in, 
        \SP_PDL_in[0]\, \SP_PDL_in[1]\, \SP_PDL_in[2]\, 
        \SP_PDL_in[3]\, \SP_PDL_in[4]\, \SP_PDL_in[5]\, 
        \SP_PDL_in[6]\, \SP_PDL_in[7]\, \SP_PDL_in[8]\, 
        \SP_PDL_in[9]\, \SP_PDL_in[10]\, \SP_PDL_in[11]\, 
        \SP_PDL_in[12]\, \SP_PDL_in[13]\, \SP_PDL_in[14]\, 
        \SP_PDL_in[15]\, \SP_PDL_in[16]\, \SP_PDL_in[17]\, 
        \SP_PDL_in[18]\, \SP_PDL_in[19]\, \SP_PDL_in[20]\, 
        \SP_PDL_in[21]\, \SP_PDL_in[22]\, \SP_PDL_in[23]\, 
        \SP_PDL_in[24]\, \SP_PDL_in[25]\, \SP_PDL_in[26]\, 
        \SP_PDL_in[27]\, \SP_PDL_in[28]\, \SP_PDL_in[29]\, 
        \SP_PDL_in[30]\, \SP_PDL_in[31]\, \SP_PDL_in[32]\, 
        \SP_PDL_in[33]\, \SP_PDL_in[34]\, \SP_PDL_in[35]\, 
        \SP_PDL_in[36]\, \SP_PDL_in[37]\, \SP_PDL_in[38]\, 
        \SP_PDL_in[39]\, \SP_PDL_in[40]\, \SP_PDL_in[41]\, 
        \SP_PDL_in[42]\, \SP_PDL_in[43]\, \SP_PDL_in[44]\, 
        \SP_PDL_in[45]\, \SP_PDL_in[46]\, \SP_PDL_in[47]\, 
        \VAD_in[1]\, \VAD_in[2]\, \VAD_in[3]\, \VAD_in[4]\, 
        \VAD_in[5]\, \VAD_in[6]\, \VAD_in[7]\, \VAD_in[8]\, 
        \VAD_in[9]\, \VAD_in[10]\, \VAD_in[11]\, \VAD_in[12]\, 
        \VAD_in[13]\, \VAD_in[14]\, \VAD_in[15]\, \VAD_in[28]\, 
        \VAD_in[29]\, \VAD_in[30]\, \VAD_in[31]\, \VDB_in[0]\, 
        \VDB_in[1]\, \VDB_in[2]\, \VDB_in[3]\, \VDB_in[4]\, 
        \VDB_in[5]\, \VDB_in[6]\, \VDB_in[7]\, \VDB_in[8]\, 
        \VDB_in[9]\, \VDB_in[10]\, \VDB_in[11]\, \VDB_in[12]\, 
        \VDB_in[13]\, \VDB_in[14]\, \VDB_in[15]\, \VDB_in[16]\, 
        \VDB_in[17]\, \VDB_in[18]\, \VDB_in[19]\, \VDB_in[20]\, 
        \VDB_in[21]\, \VDB_in[22]\, \VDB_in[23]\, \VDB_in[24]\, 
        \VDB_in[25]\, \VDB_in[26]\, \VDB_in[27]\, \VDB_in[28]\, 
        \VDB_in[29]\, \VDB_in[30]\, \VDB_in[31]\, 
        \I10.un2_evread[14]\, \I2.N_441\, \I2.N_2052\, \d_m7\, 
        d_N_3, d_N_5, d_N_7, PON_LOAD_i, HWRES_c_i_0, CLEAR_i_0, 
        \REG_i_0[80]\, \REG_i_0[121]\, \REG_i_0[265]\, 
        \REG_i_0[266]\, \REG_i_0[280]\, \REG_i_0[281]\, 
        \REG_i_0[282]\, \REG_i_0[283]\, \REG_i_0[284]\, 
        \REG_i_0[285]\, \REG_i_0[286]\, \REG_i_0[287]\, 
        \REG_i_0[288]\, \REG_i_0[289]\, \REG_i_0[290]\, 
        \REG_i_0[291]\, \REG_i_0[292]\, \REG_i_0[293]\, 
        \REG_i_0[294]\, \REG_i_0[295]\, \REG_i_0[296]\, 
        \REG_i_0[398]\, \REG_i_0[396]\, \REG_i_0[400]\, 
        \REG_i_0[5]\, NSELCLK_c_i_0, \REG_i_0[393]\, 
        \REG_i_0[394]\, \REG_i_0[395]\, \REG_i_0[397]\, 
        \REG_i_0[399]\, \I2.un5_noe16ri_i_0\, 
        \I2.un7_noe32ri_i_0\, \I2.LB_nOE_i_0\, NOEAD_c_i_0, 
        \I2.LB_nOE_i_0_0\, \I2.LB_nOE_i_0_1\, \I2.N_2613_0\, 
        \VDB_in_0[15]\, \VDB_in_0[14]\, \VDB_in_0[13]\, 
        \VDB_in_0[12]\, \VDB_in_0[11]\, \VDB_in_0[10]\, 
        \VDB_in_0[9]\, \VDB_in_0[8]\, \VDB_in_0[7]\, 
        \VDB_in_0[6]\, \VDB_in_0[5]\, \VDB_in_0[4]\, 
        \VDB_in_0[3]\, \VDB_in_0[2]\, \VDB_in_0[1]\, 
        \VDB_in_0[0]\, RUN_c_0, \LBSP_c_0[2]\, \LBSP_c_1[2]\, 
        NOEAD_c_0, NOEAD_c_1, HWRES_c_0, HWRES_c_1, HWRES_c_2, 
        HWRES_c_3, HWRES_c_4, HWRES_c_5, HWRES_c_6, HWRES_c_7, 
        HWRES_c_8, HWRES_c_9, HWRES_c_10, HWRES_c_11, HWRES_c_12, 
        HWRES_c_13, HWRES_c_14, HWRES_c_15, HWRES_c_16, 
        HWRES_c_17, HWRES_c_18, HWRES_c_19, HWRES_c_20, 
        HWRES_c_21, HWRES_c_22, HWRES_c_23, HWRES_c_24, 
        HWRES_c_25, HWRES_c_26, HWRES_c_27, HWRES_c_28, 
        HWRES_c_29, HWRES_c_30, HWRES_c_31, HWRES_c_32, 
        HWRES_c_33, HWRES_c_34, HWRES_c_35, HWRES_c_36, 
        MD_PDL_c_0, MD_PDL_c_1, MD_PDL_c_2, MD_PDL_c_3, 
        \I5.sstate_0[2]\, \I2.un7_noe32ri_0\, \I2.un5_noe16ri_0\, 
        \REG_0[127]\, \REG_0[126]\, \REG_0[125]\, \REG_0[124]\, 
        CLEAR_0, CLEAR_2, CLEAR_3, CLEAR_4, CLEAR_5, CLEAR_6, 
        CLEAR_7, CLEAR_8, CLEAR_9, CLEAR_10, CLEAR_11, CLEAR_12, 
        CLEAR_13, CLEAR_14, CLEAR_15, CLEAR_16, CLEAR_17, 
        CLEAR_18, CLEAR_19, CLEAR_20, CLEAR_21, CLEAR_22, 
        CLEAR_23, CLEAR_24, CLEAR_25, CLEAR_26, CLEAR_27, 
        CLEAR_28, \PDLCFG_DT_0[0]\, \PDLCFG_DT_1[0]\, 
        \PDLCFG_DT_2[0]\, \PDLCFG_DT_3[0]\, \TICK_0[2]\, 
        \TICK_0[0]\, \TICK_1[0]\, \TICK_2[0]\, HWRES_c_36_0, 
        HWRES_c_32_0, HWRES_c_23_0, HWRES_c_22_0, HWRES_c_21_0, 
        HWRES_c_13_0, HWRES_c_10_0, HWRES_c_0_0, HWRES_c_0_2, 
        HWRES_c_0_3, HWRES_c_0_4, HWRES_c_0_5, HWRES_c_0_6, 
        NOEAD_c_0_0, NPWON_c_0, NPWON_c_1, NPWON_c_2, NPWON_c_3, 
        LOAD_RES_0, LOAD_RES_1, LOAD_RES_2, LOAD_RES_3, 
        \PDLCFG_DT_0_0[0]\, HWRES_c_27_0, HWRES_c_7_0, RUN_c_0_0, 
        HWRES_c_0_6_0, \I5.sstate_0_i_0[2]\, \I_8\, \I_16\
         : std_logic;

    for all : PDL_INTERF
	Use entity work.PDL_INTERF(DEF_ARCH);
    for all : PDLCFG
	Use entity work.PDLCFG(DEF_ARCH);
    for all : VINTERF
	Use entity work.VINTERF(DEF_ARCH);
    for all : CROM
	Use entity work.CROM(DEF_ARCH);
    for all : RESET_MOD
	Use entity work.RESET_MOD(DEF_ARCH);
    for all : SPI_INTERF
	Use entity work.SPI_INTERF(DEF_ARCH);
    for all : ROC32
	Use entity work.ROC32(DEF_ARCH);
    for all : I2C_INTERF
	Use entity work.I2C_INTERF(DEF_ARCH);
    for all : ctrl
	Use entity work.ctrl(DEF_ARCH);
    for all : DAC_INTERF
	Use entity work.DAC_INTERF(DEF_ARCH);
    for all : DACCFG
	Use entity work.DACCFG(DEF_ARCH);
begin 


    \VDB_pad_0[11]\ : BFR
      port map(A => \VDB_in[11]\, Y => \VDB_in_0[11]\);
    
    \VDB_pad_0[2]\ : BFR
      port map(A => \VDB_in[2]\, Y => \VDB_in_0[2]\);
    
    \AE_PDL_pad[0]\ : OB33PH
      port map(PAD => AE_PDL(0), A => \AE_PDL_c[0]\);
    
    NLBLAST_pad : OB33PH
      port map(PAD => NLBLAST, A => NLBLAST_c);
    
    \VDB_pad[9]\ : IOB33PH
      port map(PAD => VDB(9), A => \I2.VDBm[9]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[9]\);
    
    \P_PDL_pad[1]\ : OB33PH
      port map(PAD => P_PDL(1), A => \P_PDL_c[1]\);
    
    \AE_PDL_pad[20]\ : OB33PH
      port map(PAD => AE_PDL(20), A => \AE_PDL_c[20]\);
    
    \LB_pad[16]\ : IOB33PH
      port map(PAD => LB(16), A => \I2.LB_i[16]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[16]\);
    
    \LB_pad[20]\ : IOB33PH
      port map(PAD => LB(20), A => \I2.LB_i[20]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[20]\);
    
    \LBSP_pad[22]\ : IOB33PH
      port map(PAD => LBSP(22), A => \REG[367]\, EN => 
        \REG_i_0[287]\, Y => \LBSP_in[22]\);
    
    \TST_pad_i[6]\ : INV
      port map(A => \I2.un5_noe16ri_0\, Y => \I2.un5_noe16ri_i_0\);
    
    \SP_PDL_pad[20]\ : IOB33PH
      port map(PAD => SP_PDL(20), A => \I3.P0[20]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[20]\);
    
    \VDB_pad_0[14]\ : BFR
      port map(A => \VDB_in[14]\, Y => \VDB_in_0[14]\);
    
    LCLK_pad : GL33
      port map(PAD => LCLK, GL => CLK_c_c);
    
    APACLK0_pad : OB33PH
      port map(PAD => APACLK0, A => CLK_c_c);
    
    \SP_PDL_pad[22]\ : IOB33PH
      port map(PAD => SP_PDL(22), A => \I3.P0[22]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[22]\);
    
    \LBSP_pad[7]\ : OB33PH
      port map(PAD => LBSP(7), A => L2A_c_c);
    
    NOEDTK_pad : OB33PH
      port map(PAD => NOEDTK, A => \TST_c_c[3]\);
    
    \LB_pad[28]\ : IOB33PH
      port map(PAD => LB(28), A => \I2.LB_i[28]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[28]\);
    
    \VDB_pad[26]\ : IOB33PH
      port map(PAD => VDB(26), A => \I2.VDBm[26]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[26]\);
    
    \SP_PDL_pad[6]\ : IOB33PH
      port map(PAD => SP_PDL(6), A => \I3.P0[6]\, EN => MD_PDL_c, 
        Y => \SP_PDL_in[6]\);
    
    RSELD0_pad : OTB33PH
      port map(PAD => RSELD0, A => \REG[378]\, EN => 
        \REG_i_0[394]\);
    
    \LB_pad[29]\ : IOB33PH
      port map(PAD => LB(29), A => \I2.LB_i[29]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[29]\);
    
    \SYNC_pad[13]\ : OB33PH
      port map(PAD => SYNC(13), A => \SYNC_c[13]\);
    
    \AE_PDL_pad[29]\ : OB33PH
      port map(PAD => AE_PDL(29), A => \AE_PDL_c[29]\);
    
    \VDB_pad[2]\ : IOB33PH
      port map(PAD => VDB(2), A => \I2.VDBm[2]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[2]\);
    
    F_SI_pad : OTB33PH
      port map(PAD => F_SI, A => \I5.ISI\, EN => un1_drive_spi);
    
    \LB_pad[14]\ : IOB33PH
      port map(PAD => LB(14), A => \I2.LB_i[14]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[14]\);
    
    \TST_pad[9]\ : OTB33PH
      port map(PAD => TST(9), A => \GND\, EN => \GND\);
    
    \LB_pad[26]\ : IOB33PH
      port map(PAD => LB(26), A => \I2.LB_i[26]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[26]\);
    
    \LBSP_pad[5]\ : OB33PH
      port map(PAD => LBSP(5), A => L1A_c_c);
    
    SCL0_pad : OB33PH
      port map(PAD => SCL0, A => SCLA_i_a3);
    
    nLBRDY_pad : IB33
      port map(PAD => nLBRDY, Y => nLBRDY_c);
    
    \SP_PDL_pad[47]\ : IOB33PH
      port map(PAD => SP_PDL(47), A => \I3.P0[47]\, EN => 
        MD_PDL_c, Y => \SP_PDL_in[47]\);
    
    BNCRES_pad : IB33
      port map(PAD => BNCRES, Y => BNCRES_c);
    
    \AE_PDL_pad[31]\ : OB33PH
      port map(PAD => AE_PDL(31), A => \AE_PDL_c[31]\);
    
    PSM_SP5_pad : IB33
      port map(PAD => PSM_SP5, Y => \REG_c[23]\);
    
    \LBSP_pad[20]\ : IOB33PH
      port map(PAD => LBSP(20), A => \REG[365]\, EN => 
        \REG_i_0[285]\, Y => \LBSP_in[20]\);
    
    \VDB_pad[17]\ : IOB33PH
      port map(PAD => VDB(17), A => \I2.VDBm[17]\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[17]\);
    
    RSELB1_pad : OTB33PH
      port map(PAD => RSELB1, A => \REG[381]\, EN => 
        \REG_i_0[397]\);
    
    \AE_PDL_pad[9]\ : OB33PH
      port map(PAD => AE_PDL(9), A => \AE_PDL_c[9]\);
    
    \LB_pad[11]\ : IOB33PH
      port map(PAD => LB(11), A => \I2.LB_i[11]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[11]\);
    
    \AE_PDL_pad[5]\ : OB33PH
      port map(PAD => AE_PDL(5), A => \AE_PDL_c[5]\);
    
    LWORDB_pad : IOB33PH
      port map(PAD => LWORDB, A => \I2.VADm[0]\, EN => NOEAD_c_0, 
        Y => LWORDB_in);
    
    \GA_pad[1]\ : IB33
      port map(PAD => GA(1), Y => \GA_c[1]\);
    
    \VDB_pad[25]\ : IOB33PH
      port map(PAD => VDB(25), A => \I2.VDBm[25]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[25]\);
    
    \LB_pad[24]\ : IOB33PH
      port map(PAD => LB(24), A => \I2.LB_i[24]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[24]\);
    
    \VDB_pad_0[15]\ : BFR
      port map(A => \VDB_in[15]\, Y => \VDB_in_0[15]\);
    
    \LBSP_pad[24]\ : IOB33PH
      port map(PAD => LBSP(24), A => \REG[369]\, EN => 
        \REG_i_0[289]\, Y => \LBSP_in[24]\);
    
    \GA_pad[3]\ : IB33
      port map(PAD => GA(3), Y => \GA_c[3]\);
    
    NPWON_pad : IB33
      port map(PAD => NPWON, Y => NPWON_c);
    
    \AE_PDL_pad[10]\ : OB33PH
      port map(PAD => AE_PDL(10), A => \AE_PDL_c[10]\);
    
    \VDB_pad[8]\ : IOB33PH
      port map(PAD => VDB(8), A => \I2.VDBm[8]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[8]\);
    
    \VDB_pad[18]\ : IOB33PH
      port map(PAD => VDB(18), A => \I2.VDBm[18]\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[18]\);
    
    \LB_pad[15]\ : IOB33PH
      port map(PAD => LB(15), A => \I2.LB_i[15]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[15]\);
    
    I3 : PDL_INTERF
      port map(PULSE(8) => \PULSE[8]\, P_PDL_c(7) => \P_PDL_c[7]\, 
        P_PDL_c(6) => \P_PDL_c[6]\, P_PDL_c(5) => \P_PDL_c[5]\, 
        P_PDL_c(4) => \P_PDL_c[4]\, P_PDL_c(3) => \P_PDL_c[3]\, 
        P_PDL_c(2) => \P_PDL_c[2]\, P_PDL_c(1) => \P_PDL_c[1]\, 
        PDL_RDATA(7) => \PDL_RDATA[7]\, PDL_RDATA(6) => 
        \PDL_RDATA[6]\, PDL_RDATA(5) => \PDL_RDATA[5]\, 
        PDL_RDATA(4) => \PDL_RDATA[4]\, PDL_RDATA(3) => 
        \PDL_RDATA[3]\, PDL_RDATA(2) => \PDL_RDATA[2]\, 
        PDL_RDATA(1) => \PDL_RDATA[1]\, PDL_RDATA(0) => 
        \PDL_RDATA[0]\, PDL_RADDR(5) => \PDL_RADDR[5]\, 
        PDL_RADDR(4) => \PDL_RADDR[4]\, PDL_RADDR(3) => 
        \PDL_RADDR[3]\, PDL_RADDR(2) => \PDL_RADDR[2]\, 
        PDL_RADDR(1) => \PDL_RADDR[1]\, PDL_RADDR(0) => 
        \PDL_RADDR[0]\, PDLCFG_RAD(5) => \PDLCFG_RAD[5]\, 
        PDLCFG_RAD(4) => \PDLCFG_RAD[4]\, PDLCFG_RAD(3) => 
        \PDLCFG_RAD[3]\, PDLCFG_RAD(2) => \PDLCFG_RAD[2]\, 
        PDLCFG_RAD(1) => \PDLCFG_RAD[1]\, PDLCFG_RAD(0) => 
        \PDLCFG_RAD[0]\, PDLCFG_DT(7) => \PDLCFG_DT[7]\, 
        PDLCFG_DT(6) => \PDLCFG_DT[6]\, PDLCFG_DT(5) => 
        \PDLCFG_DT[5]\, PDLCFG_DT(4) => \PDLCFG_DT[4]\, 
        PDLCFG_DT(3) => \PDLCFG_DT[3]\, PDLCFG_DT(2) => 
        \PDLCFG_DT[2]\, PDLCFG_DT(1) => \PDLCFG_DT[1]\, 
        PDLCFG_DT(0) => \PDLCFG_DT[0]\, PDLCFG_DT_0_0(0) => 
        \PDLCFG_DT_0_0[0]\, PDLCFG_DT_3(0) => \PDLCFG_DT_3[0]\, 
        PDLCFG_DT_1(0) => \PDLCFG_DT_1[0]\, PDLCFG_DT_2(0) => 
        \PDLCFG_DT_2[0]\, PDLCFG_DT_0(0) => \PDLCFG_DT_0[0]\, 
        P0(47) => \I3.P0[47]\, P0(46) => \I3.P0[46]\, P0(45) => 
        \I3.P0[45]\, P0(44) => \I3.P0[44]\, P0(43) => \I3.P0[43]\, 
        P0(42) => \I3.P0[42]\, P0(41) => \I3.P0[41]\, P0(40) => 
        \I3.P0[40]\, P0(39) => \I3.P0[39]\, P0(38) => \I3.P0[38]\, 
        P0(37) => \I3.P0[37]\, P0(36) => \I3.P0[36]\, P0(35) => 
        \I3.P0[35]\, P0(34) => \I3.P0[34]\, P0(33) => \I3.P0[33]\, 
        P0(32) => \I3.P0[32]\, P0(31) => \I3.P0[31]\, P0(30) => 
        \I3.P0[30]\, P0(29) => \I3.P0[29]\, P0(28) => \I3.P0[28]\, 
        P0(27) => \I3.P0[27]\, P0(26) => \I3.P0[26]\, P0(25) => 
        \I3.P0[25]\, P0(24) => \I3.P0[24]\, P0(23) => \I3.P0[23]\, 
        P0(22) => \I3.P0[22]\, P0(21) => \I3.P0[21]\, P0(20) => 
        \I3.P0[20]\, P0(19) => \I3.P0[19]\, P0(18) => \I3.P0[18]\, 
        P0(17) => \I3.P0[17]\, P0(16) => \I3.P0[16]\, P0(15) => 
        \I3.P0[15]\, P0(14) => \I3.P0[14]\, P0(13) => \I3.P0[13]\, 
        P0(12) => \I3.P0[12]\, P0(11) => \I3.P0[11]\, P0(10) => 
        \I3.P0[10]\, P0(9) => \I3.P0[9]\, P0(8) => \I3.P0[8]\, 
        P0(7) => \I3.P0[7]\, P0(6) => \I3.P0[6]\, P0(5) => 
        \I3.P0[5]\, P0(4) => \I3.P0[4]\, P0(3) => \I3.P0[3]\, 
        P0(2) => \I3.P0[2]\, P0(1) => \I3.P0[1]\, P0(0) => 
        \I3.P0[0]\, AE_PDL_c(47) => \AE_PDL_c[47]\, AE_PDL_c(46)
         => \AE_PDL_c[46]\, AE_PDL_c(45) => \AE_PDL_c[45]\, 
        AE_PDL_c(44) => \AE_PDL_c[44]\, AE_PDL_c(43) => 
        \AE_PDL_c[43]\, AE_PDL_c(42) => \AE_PDL_c[42]\, 
        AE_PDL_c(41) => \AE_PDL_c[41]\, AE_PDL_c(40) => 
        \AE_PDL_c[40]\, AE_PDL_c(39) => \AE_PDL_c[39]\, 
        AE_PDL_c(38) => \AE_PDL_c[38]\, AE_PDL_c(37) => 
        \AE_PDL_c[37]\, AE_PDL_c(36) => \AE_PDL_c[36]\, 
        AE_PDL_c(35) => \AE_PDL_c[35]\, AE_PDL_c(34) => 
        \AE_PDL_c[34]\, AE_PDL_c(33) => \AE_PDL_c[33]\, 
        AE_PDL_c(32) => \AE_PDL_c[32]\, AE_PDL_c(31) => 
        \AE_PDL_c[31]\, AE_PDL_c(30) => \AE_PDL_c[30]\, 
        AE_PDL_c(29) => \AE_PDL_c[29]\, AE_PDL_c(28) => 
        \AE_PDL_c[28]\, AE_PDL_c(27) => \AE_PDL_c[27]\, 
        AE_PDL_c(26) => \AE_PDL_c[26]\, AE_PDL_c(25) => 
        \AE_PDL_c[25]\, AE_PDL_c(24) => \AE_PDL_c[24]\, 
        AE_PDL_c(23) => \AE_PDL_c[23]\, AE_PDL_c(22) => 
        \AE_PDL_c[22]\, AE_PDL_c(21) => \AE_PDL_c[21]\, 
        AE_PDL_c(20) => \AE_PDL_c[20]\, AE_PDL_c(19) => 
        \AE_PDL_c[19]\, AE_PDL_c(18) => \AE_PDL_c[18]\, 
        AE_PDL_c(17) => \AE_PDL_c[17]\, AE_PDL_c(16) => 
        \AE_PDL_c[16]\, AE_PDL_c(15) => \AE_PDL_c[15]\, 
        AE_PDL_c(14) => \AE_PDL_c[14]\, AE_PDL_c(13) => 
        \AE_PDL_c[13]\, AE_PDL_c(12) => \AE_PDL_c[12]\, 
        AE_PDL_c(11) => \AE_PDL_c[11]\, AE_PDL_c(10) => 
        \AE_PDL_c[10]\, AE_PDL_c(9) => \AE_PDL_c[9]\, AE_PDL_c(8)
         => \AE_PDL_c[8]\, AE_PDL_c(7) => \AE_PDL_c[7]\, 
        AE_PDL_c(6) => \AE_PDL_c[6]\, AE_PDL_c(5) => 
        \AE_PDL_c[5]\, AE_PDL_c(4) => \AE_PDL_c[4]\, AE_PDL_c(3)
         => \AE_PDL_c[3]\, AE_PDL_c(2) => \AE_PDL_c[2]\, 
        AE_PDL_c(1) => \AE_PDL_c[1]\, AE_PDL_c(0) => 
        \AE_PDL_c[0]\, SP_PDL_in(47) => \SP_PDL_in[47]\, 
        SP_PDL_in(46) => \SP_PDL_in[46]\, SP_PDL_in(45) => 
        \SP_PDL_in[45]\, SP_PDL_in(44) => \SP_PDL_in[44]\, 
        SP_PDL_in(43) => \SP_PDL_in[43]\, SP_PDL_in(42) => 
        \SP_PDL_in[42]\, SP_PDL_in(41) => \SP_PDL_in[41]\, 
        SP_PDL_in(40) => \SP_PDL_in[40]\, SP_PDL_in(39) => 
        \SP_PDL_in[39]\, SP_PDL_in(38) => \SP_PDL_in[38]\, 
        SP_PDL_in(37) => \SP_PDL_in[37]\, SP_PDL_in(36) => 
        \SP_PDL_in[36]\, SP_PDL_in(35) => \SP_PDL_in[35]\, 
        SP_PDL_in(34) => \SP_PDL_in[34]\, SP_PDL_in(33) => 
        \SP_PDL_in[33]\, SP_PDL_in(32) => \SP_PDL_in[32]\, 
        SP_PDL_in(31) => \SP_PDL_in[31]\, SP_PDL_in(30) => 
        \SP_PDL_in[30]\, SP_PDL_in(29) => \SP_PDL_in[29]\, 
        SP_PDL_in(28) => \SP_PDL_in[28]\, SP_PDL_in(27) => 
        \SP_PDL_in[27]\, SP_PDL_in(26) => \SP_PDL_in[26]\, 
        SP_PDL_in(25) => \SP_PDL_in[25]\, SP_PDL_in(24) => 
        \SP_PDL_in[24]\, SP_PDL_in(23) => \SP_PDL_in[23]\, 
        SP_PDL_in(22) => \SP_PDL_in[22]\, SP_PDL_in(21) => 
        \SP_PDL_in[21]\, SP_PDL_in(20) => \SP_PDL_in[20]\, 
        SP_PDL_in(19) => \SP_PDL_in[19]\, SP_PDL_in(18) => 
        \SP_PDL_in[18]\, SP_PDL_in(17) => \SP_PDL_in[17]\, 
        SP_PDL_in(16) => \SP_PDL_in[16]\, SP_PDL_in(15) => 
        \SP_PDL_in[15]\, SP_PDL_in(14) => \SP_PDL_in[14]\, 
        SP_PDL_in(13) => \SP_PDL_in[13]\, SP_PDL_in(12) => 
        \SP_PDL_in[12]\, SP_PDL_in(11) => \SP_PDL_in[11]\, 
        SP_PDL_in(10) => \SP_PDL_in[10]\, SP_PDL_in(9) => 
        \SP_PDL_in[9]\, SP_PDL_in(8) => \SP_PDL_in[8]\, 
        SP_PDL_in(7) => \SP_PDL_in[7]\, SP_PDL_in(6) => 
        \SP_PDL_in[6]\, SP_PDL_in(5) => \SP_PDL_in[5]\, 
        SP_PDL_in(4) => \SP_PDL_in[4]\, SP_PDL_in(3) => 
        \SP_PDL_in[3]\, SP_PDL_in(2) => \SP_PDL_in[2]\, 
        SP_PDL_in(1) => \SP_PDL_in[1]\, SP_PDL_in(0) => 
        \SP_PDL_in[0]\, REG_0(127) => \REG_0[127]\, REG_0(126)
         => \REG_0[126]\, REG_0(125) => \REG_0[125]\, REG_0(124)
         => \REG_0[124]\, REG_i_0(121) => \REG_i_0[121]\, REG_32
         => \REG[153]\, REG_33 => \REG[154]\, REG_34 => 
        \REG[155]\, REG_35 => \REG[156]\, REG_36 => \REG[157]\, 
        REG_37 => \REG[158]\, REG_38 => \REG[159]\, REG_39 => 
        \REG[160]\, REG_40 => \REG[161]\, REG_41 => \REG[162]\, 
        REG_42 => \REG[163]\, REG_43 => \REG[164]\, REG_44 => 
        \REG[165]\, REG_45 => \REG[166]\, REG_46 => \REG[167]\, 
        REG_47 => \REG[168]\, REG_48 => \REG[169]\, REG_49 => 
        \REG[170]\, REG_50 => \REG[171]\, REG_51 => \REG[172]\, 
        REG_52 => \REG[173]\, REG_53 => \REG[174]\, REG_54 => 
        \REG[175]\, REG_55 => \REG[176]\, REG_56 => \REG[177]\, 
        REG_57 => \REG[178]\, REG_58 => \REG[179]\, REG_59 => 
        \REG[180]\, REG_60 => \REG[181]\, REG_61 => \REG[182]\, 
        REG_62 => \REG[183]\, REG_63 => \REG[184]\, REG_64 => 
        \REG[185]\, REG_65 => \REG[186]\, REG_66 => \REG[187]\, 
        REG_67 => \REG[188]\, REG_68 => \REG[189]\, REG_69 => 
        \REG[190]\, REG_70 => \REG[191]\, REG_71 => \REG[192]\, 
        REG_72 => \REG[193]\, REG_73 => \REG[194]\, REG_74 => 
        \REG[195]\, REG_75 => \REG[196]\, REG_76 => \REG[197]\, 
        REG_77 => \REG[198]\, REG_78 => \REG[199]\, REG_79 => 
        \REG[200]\, REG_3 => \REG[124]\, REG_6 => \REG[127]\, 
        REG_5 => \REG[126]\, REG_4 => \REG[125]\, REG_2 => 
        \REG[123]\, REG_1 => \REG[122]\, REG_24 => \REG[145]\, 
        REG_9 => \REG[130]\, REG_16 => \REG[137]\, REG_10 => 
        \REG[131]\, REG_17 => \REG[138]\, REG_11 => \REG[132]\, 
        REG_18 => \REG[139]\, REG_12 => \REG[133]\, REG_19 => 
        \REG[140]\, REG_13 => \REG[134]\, REG_20 => \REG[141]\, 
        REG_14 => \REG[135]\, REG_21 => \REG[142]\, REG_15 => 
        \REG[136]\, REG_22 => \REG[143]\, REG_23 => \REG[144]\, 
        REG_0_d0 => \REG[121]\, REG_8 => \REG[129]\, MD_PDL_c => 
        MD_PDL_c, PDL_RACK => PDL_RACK, PDL_RREQ => PDL_RREQ, 
        SI_PDL_c => SI_PDL_c, PDLCFG_nRD => PDLCFG_nRD, 
        SCLK_PDL_c => SCLK_PDL_c, HWRES_c_2 => HWRES_c_2, 
        HWRES_c_1 => HWRES_c_1, MD_PDL_c_0 => MD_PDL_c_0, 
        MD_PDL_c_1 => MD_PDL_c_1, MD_PDL_c_2 => MD_PDL_c_2, 
        MD_PDL_c_3 => MD_PDL_c_3, LOAD_RES => LOAD_RES, 
        HWRES_c_0_3 => HWRES_c_0_3, HWRES_c_0_2 => HWRES_c_0_2, 
        LOAD_RES_3 => LOAD_RES_3, CLK_c_c => CLK_c_c, 
        HWRES_c_23_0 => HWRES_c_23_0, HWRES_c_0 => HWRES_c_0, 
        LOAD_RES_0 => LOAD_RES_0);
    
    I11 : PDLCFG
      port map(CROMWDT(7) => \CROMWDT[7]\, CROMWDT(6) => 
        \CROMWDT[6]\, CROMWDT(5) => \CROMWDT[5]\, CROMWDT(4) => 
        \CROMWDT[4]\, CROMWDT(3) => \CROMWDT[3]\, CROMWDT(2) => 
        \CROMWDT[2]\, CROMWDT(1) => \CROMWDT[1]\, CROMWDT(0) => 
        \CROMWDT[0]\, PDLCFG_RAD(5) => \PDLCFG_RAD[5]\, 
        PDLCFG_RAD(4) => \PDLCFG_RAD[4]\, PDLCFG_RAD(3) => 
        \PDLCFG_RAD[3]\, PDLCFG_RAD(2) => \PDLCFG_RAD[2]\, 
        PDLCFG_RAD(1) => \PDLCFG_RAD[1]\, PDLCFG_RAD(0) => 
        \PDLCFG_RAD[0]\, CROMWAD(5) => \CROMWAD[5]\, CROMWAD(4)
         => \CROMWAD[4]\, CROMWAD(3) => \CROMWAD[3]\, CROMWAD(2)
         => \CROMWAD[2]\, CROMWAD(1) => \CROMWAD[1]\, CROMWAD(0)
         => \CROMWAD[0]\, PDLCFG_DT_0(0) => \PDLCFG_DT_0[0]\, 
        PDLCFG_DT_1(0) => \PDLCFG_DT_1[0]\, PDLCFG_DT_2(0) => 
        \PDLCFG_DT_2[0]\, PDLCFG_DT_3(0) => \PDLCFG_DT_3[0]\, 
        PDLCFG_DT(7) => \PDLCFG_DT[7]\, PDLCFG_DT(6) => 
        \PDLCFG_DT[6]\, PDLCFG_DT(5) => \PDLCFG_DT[5]\, 
        PDLCFG_DT(4) => \PDLCFG_DT[4]\, PDLCFG_DT(3) => 
        \PDLCFG_DT[3]\, PDLCFG_DT(2) => \PDLCFG_DT[2]\, 
        PDLCFG_DT(1) => \PDLCFG_DT[1]\, PDLCFG_DT(0) => 
        \PDLCFG_DT[0]\, PDLCFG_DT_0_0(0) => \PDLCFG_DT_0_0[0]\, 
        PDLCFG_nRD => PDLCFG_nRD, PDLCFG_nWR => PDLCFG_nWR, 
        CLK_c_c => CLK_c_c);
    
    \LB_pad[30]\ : IOB33PH
      port map(PAD => LB(30), A => \I2.LB_i[30]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[30]\);
    
    \DIR_CTTM_pad[2]\ : OB33PH
      port map(PAD => DIR_CTTM(2), A => \VCC\);
    
    MD_PDL_pad : OB33PH
      port map(PAD => MD_PDL, A => MD_PDL_c_0);
    
    \LB_pad[21]\ : IOB33PH
      port map(PAD => LB(21), A => \I2.LB_i[21]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[21]\);
    
    \AMB_pad[0]\ : IB33
      port map(PAD => AMB(0), Y => \AMB_c[0]\);
    
    INTR2_pad : OB33PH
      port map(PAD => INTR2, A => \VCC\);
    
    d_m2 : MUX2H
      port map(A => \REG[481]\, B => \REG[409]\, S => 
        \I2.REGMAP[31]\, Y => d_N_3);
    
    \AE_PDL_pad[19]\ : OB33PH
      port map(PAD => AE_PDL(19), A => \AE_PDL_c[19]\);
    
    SYSRESB_pad : IB33
      port map(PAD => SYSRESB, Y => SYSRESB_c);
    
    NCYC_RELOAD_pad : IOB33PH
      port map(PAD => NCYC_RELOAD, A => \VCC\, EN => 
        \I5.DRIVE_RELOAD\, Y => NCYC_RELOAD_in);
    
    \VDB_pad[29]\ : IOB33PH
      port map(PAD => VDB(29), A => \I2.VDBm[29]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[29]\);
    
    DS0B_pad : IB33
      port map(PAD => DS0B, Y => DS0B_c);
    
    \AE_PDL_pad[34]\ : OB33PH
      port map(PAD => AE_PDL(34), A => \AE_PDL_c[34]\);
    
    \LB_pad[0]\ : IOB33PH
      port map(PAD => LB(0), A => \I2.LB_i[0]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[0]\);
    
    \AE_PDL_pad[35]\ : OB33PH
      port map(PAD => AE_PDL(35), A => \AE_PDL_c[35]\);
    
    \VDB_pad_0[7]\ : BFR
      port map(A => \VDB_in[7]\, Y => \VDB_in_0[7]\);
    
    \AMB_pad[2]\ : IB33
      port map(PAD => AMB(2), Y => \AMB_c[2]\);
    
    \SYNC_pad[5]\ : OB33PH
      port map(PAD => SYNC(5), A => \SYNC_c[5]\);
    
    EVRES_pad : IB33
      port map(PAD => EVRES, Y => EVRES_c);
    
    NOE16R_pad : OB33PH
      port map(PAD => NOE16R, A => \I2.un5_noe16ri_i_0\);
    
    \LB_pad[25]\ : IOB33PH
      port map(PAD => LB(25), A => \I2.LB_i[25]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[25]\);
    
    \GA_pad[0]\ : IB33
      port map(PAD => GA(0), Y => \GA_c[0]\);
    
    NLBCLR_pad : OB33PH
      port map(PAD => NLBCLR, A => NLBCLR_c);
    
    WRITEB_pad : IB33
      port map(PAD => WRITEB, Y => WRITEB_c);
    
    RSELD1_pad : OTB33PH
      port map(PAD => RSELD1, A => \REG[377]\, EN => 
        \REG_i_0[393]\);
    
    \VDB_pad_0[8]\ : BFR
      port map(A => \VDB_in[8]\, Y => \VDB_in_0[8]\);
    
    \VDB_pad[10]\ : IOB33PH
      port map(PAD => VDB(10), A => \I2.VDBm[10]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[10]\);
    
    \SP_PDL_pad[27]\ : IOB33PH
      port map(PAD => SP_PDL(27), A => \I3.P0[27]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[27]\);
    
    \AE_PDL_pad[38]\ : OB33PH
      port map(PAD => AE_PDL(38), A => \AE_PDL_c[38]\);
    
    I2 : VINTERF
      port map(TICK(2) => \TICK[2]\, RAMDT(7) => \RAMDT[7]\, 
        RAMDT(6) => \RAMDT[6]\, RAMDT(5) => \RAMDT[5]\, RAMDT(4)
         => \RAMDT[4]\, RAMDT(3) => \RAMDT[3]\, RAMDT(2) => 
        \RAMDT[2]\, RAMDT(1) => \RAMDT[1]\, RAMDT(0) => 
        \RAMDT[0]\, VADm(31) => \I2.VADm[31]\, VADm(30) => 
        \I2.VADm[30]\, VADm(29) => \I2.VADm[29]\, VADm(28) => 
        \I2.VADm[28]\, VADm(27) => \I2.VADm[27]\, VADm(26) => 
        \I2.VADm[26]\, VADm(25) => \I2.VADm[25]\, VADm(24) => 
        \I2.VADm[24]\, VADm(23) => \I2.VADm[23]\, VADm(22) => 
        \I2.VADm[22]\, VADm(21) => \I2.VADm[21]\, VADm(20) => 
        \I2.VADm[20]\, VADm(19) => \I2.VADm[19]\, VADm(18) => 
        \I2.VADm[18]\, VADm(17) => \I2.VADm[17]\, VADm(16) => 
        \I2.VADm[16]\, VADm(15) => \I2.VADm[15]\, VADm(14) => 
        \I2.VADm[14]\, VADm(13) => \I2.VADm[13]\, VADm(12) => 
        \I2.VADm[12]\, VADm(11) => \I2.VADm[11]\, VADm(10) => 
        \I2.VADm[10]\, VADm(9) => \I2.VADm[9]\, VADm(8) => 
        \I2.VADm[8]\, VADm(7) => \I2.VADm[7]\, VADm(6) => 
        \I2.VADm[6]\, VADm(5) => \I2.VADm[5]\, VADm(4) => 
        \I2.VADm[4]\, VADm(3) => \I2.VADm[3]\, VADm(2) => 
        \I2.VADm[2]\, VADm(1) => \I2.VADm[1]\, VADm(0) => 
        \I2.VADm[0]\, RAMAD_VME(8) => \RAMAD_VME[8]\, 
        RAMAD_VME(7) => \RAMAD_VME[7]\, RAMAD_VME(6) => 
        \RAMAD_VME[6]\, RAMAD_VME(5) => \RAMAD_VME[5]\, 
        RAMAD_VME(4) => \RAMAD_VME[4]\, RAMAD_VME(3) => 
        \RAMAD_VME[3]\, RAMAD_VME(2) => \RAMAD_VME[2]\, 
        RAMAD_VME(1) => \RAMAD_VME[1]\, RAMAD_VME(0) => 
        \RAMAD_VME[0]\, AMB_c(5) => \AMB_c[5]\, AMB_c(4) => 
        \AMB_c[4]\, AMB_c(3) => \AMB_c[3]\, AMB_c(2) => 
        \AMB_c[2]\, AMB_c(1) => \AMB_c[1]\, AMB_c(0) => 
        \AMB_c[0]\, LB_in(31) => \LB_in[31]\, LB_in(30) => 
        \LB_in[30]\, LB_in(29) => \LB_in[29]\, LB_in(28) => 
        \LB_in[28]\, LB_in(27) => \LB_in[27]\, LB_in(26) => 
        \LB_in[26]\, LB_in(25) => \LB_in[25]\, LB_in(24) => 
        \LB_in[24]\, LB_in(23) => \LB_in[23]\, LB_in(22) => 
        \LB_in[22]\, LB_in(21) => \LB_in[21]\, LB_in(20) => 
        \LB_in[20]\, LB_in(19) => \LB_in[19]\, LB_in(18) => 
        \LB_in[18]\, LB_in(17) => \LB_in[17]\, LB_in(16) => 
        \LB_in[16]\, LB_in(15) => \LB_in[15]\, LB_in(14) => 
        \LB_in[14]\, LB_in(13) => \LB_in[13]\, LB_in(12) => 
        \LB_in[12]\, LB_in(11) => \LB_in[11]\, LB_in(10) => 
        \LB_in[10]\, LB_in(9) => \LB_in[9]\, LB_in(8) => 
        \LB_in[8]\, LB_in(7) => \LB_in[7]\, LB_in(6) => 
        \LB_in[6]\, LB_in(5) => \LB_in[5]\, LB_in(4) => 
        \LB_in[4]\, LB_in(3) => \LB_in[3]\, LB_in(2) => 
        \LB_in[2]\, LB_in(1) => \LB_in[1]\, LB_in(0) => 
        \LB_in[0]\, OR_RDATA(9) => \OR_RDATA[9]\, OR_RDATA(8) => 
        \OR_RDATA[8]\, OR_RDATA(7) => \OR_RDATA[7]\, OR_RDATA(6)
         => \OR_RDATA[6]\, OR_RDATA(5) => \OR_RDATA[5]\, 
        OR_RDATA(4) => \OR_RDATA[4]\, OR_RDATA(3) => 
        \OR_RDATA[3]\, OR_RDATA(2) => \OR_RDATA[2]\, OR_RDATA(1)
         => \OR_RDATA[1]\, OR_RDATA(0) => \OR_RDATA[0]\, PULSE_0
         => \PULSE[0]\, PULSE_1 => \PULSE[1]\, PULSE_2 => 
        \PULSE[2]\, PULSE_3 => \PULSE[3]\, PULSE_6 => \PULSE[6]\, 
        PULSE_7 => \PULSE[7]\, PULSE_8 => \PULSE[8]\, PULSE_9 => 
        \PULSE[9]\, PULSE_10 => \PULSE[10]\, OR_RADDR(5) => 
        \OR_RADDR[5]\, OR_RADDR(4) => \OR_RADDR[4]\, OR_RADDR(3)
         => \OR_RADDR[3]\, OR_RADDR(2) => \OR_RADDR[2]\, 
        OR_RADDR(1) => \OR_RADDR[1]\, OR_RADDR(0) => 
        \OR_RADDR[0]\, VDB_in_0(15) => \VDB_in_0[15]\, 
        VDB_in_0(14) => \VDB_in_0[14]\, VDB_in_0(13) => 
        \VDB_in_0[13]\, VDB_in_0(12) => \VDB_in_0[12]\, 
        VDB_in_0(11) => \VDB_in_0[11]\, VDB_in_0(10) => 
        \VDB_in_0[10]\, VDB_in_0(9) => \VDB_in_0[9]\, VDB_in_0(8)
         => \VDB_in_0[8]\, VDB_in_0(7) => \VDB_in_0[7]\, 
        VDB_in_0(6) => \VDB_in_0[6]\, VDB_in_0(5) => 
        \VDB_in_0[5]\, VDB_in_0(4) => \VDB_in_0[4]\, VDB_in_0(3)
         => \VDB_in_0[3]\, VDB_in_0(2) => \VDB_in_0[2]\, 
        VDB_in_0(1) => \VDB_in_0[1]\, VDB_in_0(0) => 
        \VDB_in_0[0]\, VDB_in(31) => \VDB_in[31]\, VDB_in(30) => 
        \VDB_in[30]\, VDB_in(29) => \VDB_in[29]\, VDB_in(28) => 
        \VDB_in[28]\, VDB_in(27) => \VDB_in[27]\, VDB_in(26) => 
        \VDB_in[26]\, VDB_in(25) => \VDB_in[25]\, VDB_in(24) => 
        \VDB_in[24]\, VDB_in(23) => \VDB_in[23]\, VDB_in(22) => 
        \VDB_in[22]\, VDB_in(21) => \VDB_in[21]\, VDB_in(20) => 
        \VDB_in[20]\, VDB_in(19) => \VDB_in[19]\, VDB_in(18) => 
        \VDB_in[18]\, VDB_in(17) => \VDB_in[17]\, VDB_in(16) => 
        \VDB_in[16]\, VDB_in(15) => \VDB_in[15]\, VDB_in(14) => 
        \VDB_in[14]\, VDB_in(13) => \VDB_in[13]\, VDB_in(12) => 
        \VDB_in[12]\, VDB_in(11) => \VDB_in[11]\, VDB_in(10) => 
        \VDB_in[10]\, VDB_in(9) => \VDB_in[9]\, VDB_in(8) => 
        \VDB_in[8]\, VDB_in(7) => \VDB_in[7]\, VDB_in(6) => 
        \VDB_in[6]\, VDB_in(5) => \VDB_in[5]\, VDB_in(4) => 
        \VDB_in[4]\, VDB_in(3) => \VDB_in[3]\, VDB_in(2) => 
        \VDB_in[2]\, VDB_in(1) => \VDB_in[1]\, VDB_in(0) => 
        \VDB_in[0]\, LB_i(31) => \I2.LB_i[31]\, LB_i(30) => 
        \I2.LB_i[30]\, LB_i(29) => \I2.LB_i[29]\, LB_i(28) => 
        \I2.LB_i[28]\, LB_i(27) => \I2.LB_i[27]\, LB_i(26) => 
        \I2.LB_i[26]\, LB_i(25) => \I2.LB_i[25]\, LB_i(24) => 
        \I2.LB_i[24]\, LB_i(23) => \I2.LB_i[23]\, LB_i(22) => 
        \I2.LB_i[22]\, LB_i(21) => \I2.LB_i[21]\, LB_i(20) => 
        \I2.LB_i[20]\, LB_i(19) => \I2.LB_i[19]\, LB_i(18) => 
        \I2.LB_i[18]\, LB_i(17) => \I2.LB_i[17]\, LB_i(16) => 
        \I2.LB_i[16]\, LB_i(15) => \I2.LB_i[15]\, LB_i(14) => 
        \I2.LB_i[14]\, LB_i(13) => \I2.LB_i[13]\, LB_i(12) => 
        \I2.LB_i[12]\, LB_i(11) => \I2.LB_i[11]\, LB_i(10) => 
        \I2.LB_i[10]\, LB_i(9) => \I2.LB_i[9]\, LB_i(8) => 
        \I2.LB_i[8]\, LB_i(7) => \I2.LB_i[7]\, LB_i(6) => 
        \I2.LB_i[6]\, LB_i(5) => \I2.LB_i[5]\, LB_i(4) => 
        \I2.LB_i[4]\, LB_i(3) => \I2.LB_i[3]\, LB_i(2) => 
        \I2.LB_i[2]\, LB_i(1) => \I2.LB_i[1]\, LB_i(0) => 
        \I2.LB_i[0]\, DPR(31) => \DPR[31]\, DPR(30) => \DPR[30]\, 
        DPR(29) => \DPR[29]\, DPR(28) => \DPR[28]\, DPR(27) => 
        \DPR[27]\, DPR(26) => \DPR[26]\, DPR(25) => \DPR[25]\, 
        DPR(24) => \DPR[24]\, DPR(23) => \DPR[23]\, DPR(22) => 
        \DPR[22]\, DPR(21) => \DPR[21]\, DPR(20) => \DPR[20]\, 
        DPR(19) => \DPR[19]\, DPR(18) => \DPR[18]\, DPR(17) => 
        \DPR[17]\, DPR(16) => \DPR[16]\, DPR(15) => \DPR[15]\, 
        DPR(14) => \DPR[14]\, DPR(13) => \DPR[13]\, DPR(12) => 
        \DPR[12]\, DPR(11) => \DPR[11]\, DPR(10) => \DPR[10]\, 
        DPR(9) => \DPR[9]\, DPR(8) => \DPR[8]\, DPR(7) => 
        \DPR[7]\, DPR(6) => \DPR[6]\, DPR(5) => \DPR[5]\, DPR(4)
         => \DPR[4]\, DPR(3) => \DPR[3]\, DPR(2) => \DPR[2]\, 
        DPR(1) => \DPR[1]\, DPR(0) => \DPR[0]\, FBOUT(7) => 
        \FBOUT[7]\, FBOUT(6) => \FBOUT[6]\, FBOUT(5) => 
        \FBOUT[5]\, FBOUT(4) => \FBOUT[4]\, FBOUT(3) => 
        \FBOUT[3]\, FBOUT(2) => \FBOUT[2]\, FBOUT(1) => 
        \FBOUT[1]\, FBOUT(0) => \FBOUT[0]\, LBSP_c(2) => 
        \LBSP_c[2]\, REGMAP_35 => \I2.REGMAP[35]\, REGMAP_31 => 
        \I2.REGMAP[31]\, REG_c_21 => \REG_c[21]\, REG_c_22 => 
        \REG_c[22]\, REG_c_23 => \REG_c[23]\, REG_c_0 => 
        \REG_c[0]\, LBSP_in_0 => \LBSP_in[0]\, LBSP_in_1 => 
        \LBSP_in[1]\, LBSP_in_15 => \LBSP_in[15]\, LBSP_in_16 => 
        \LBSP_in[16]\, LBSP_in_17 => \LBSP_in[17]\, LBSP_in_18
         => \LBSP_in[18]\, LBSP_in_19 => \LBSP_in[19]\, 
        LBSP_in_20 => \LBSP_in[20]\, LBSP_in_21 => \LBSP_in[21]\, 
        LBSP_in_22 => \LBSP_in[22]\, LBSP_in_23 => \LBSP_in[23]\, 
        LBSP_in_24 => \LBSP_in[24]\, LBSP_in_25 => \LBSP_in[25]\, 
        LBSP_in_26 => \LBSP_in[26]\, LBSP_in_27 => \LBSP_in[27]\, 
        LBSP_in_28 => \LBSP_in[28]\, LBSP_in_29 => \LBSP_in[29]\, 
        LBSP_in_30 => \LBSP_in[30]\, LBSP_in_31 => \LBSP_in[31]\, 
        VAD_in_0 => \VAD_in[1]\, VAD_in_1 => \VAD_in[2]\, 
        VAD_in_2 => \VAD_in[3]\, VAD_in_3 => \VAD_in[4]\, 
        VAD_in_4 => \VAD_in[5]\, VAD_in_5 => \VAD_in[6]\, 
        VAD_in_6 => \VAD_in[7]\, VAD_in_7 => \VAD_in[8]\, 
        VAD_in_8 => \VAD_in[9]\, VAD_in_9 => \VAD_in[10]\, 
        VAD_in_10 => \VAD_in[11]\, VAD_in_11 => \VAD_in[12]\, 
        VAD_in_12 => \VAD_in[13]\, VAD_in_13 => \VAD_in[14]\, 
        VAD_in_14 => \VAD_in[15]\, VAD_in_27 => \VAD_in[28]\, 
        VAD_in_28 => \VAD_in[29]\, VAD_in_29 => \VAD_in[30]\, 
        VAD_in_30 => \VAD_in[31]\, GA_c(3) => \GA_c[3]\, GA_c(2)
         => \GA_c[2]\, GA_c(1) => \GA_c[1]\, GA_c(0) => \GA_c[0]\, 
        VDBm_0 => \I2.VDBm[0]\, VDBm_1 => \I2.VDBm[1]\, VDBm_2
         => \I2.VDBm[2]\, VDBm_3 => \I2.VDBm[3]\, VDBm_4 => 
        \I2.VDBm[4]\, VDBm_5 => \I2.VDBm[5]\, VDBm_6 => 
        \I2.VDBm[6]\, VDBm_7 => \I2.VDBm[7]\, VDBm_8 => 
        \I2.VDBm[8]\, VDBm_9 => \I2.VDBm[9]\, VDBm_10 => 
        \I2.VDBm[10]\, VDBm_12 => \I2.VDBm[12]\, VDBm_13 => 
        \I2.VDBm[13]\, VDBm_14 => \I2.VDBm[14]\, VDBm_15 => 
        \I2.VDBm[15]\, VDBm_16 => \I2.VDBm[16]\, VDBm_17 => 
        \I2.VDBm[17]\, VDBm_18 => \I2.VDBm[18]\, VDBm_19 => 
        \I2.VDBm[19]\, VDBm_20 => \I2.VDBm[20]\, VDBm_22 => 
        \I2.VDBm[22]\, VDBm_23 => \I2.VDBm[23]\, VDBm_24 => 
        \I2.VDBm[24]\, VDBm_25 => \I2.VDBm[25]\, VDBm_26 => 
        \I2.VDBm[26]\, VDBm_27 => \I2.VDBm[27]\, VDBm_28 => 
        \I2.VDBm[28]\, VDBm_29 => \I2.VDBm[29]\, VDBm_30 => 
        \I2.VDBm[30]\, VDBm_31 => \I2.VDBm[31]\, VDBm_i_m2(11)
         => \VDBm_i_m2[11]\, REG_126 => \REG[127]\, REG_125 => 
        \REG[126]\, REG_124 => \REG[125]\, REG_123 => \REG[124]\, 
        REG_344 => \REG[345]\, REG_345 => \REG[346]\, REG_359 => 
        \REG[360]\, REG_360 => \REG[361]\, REG_361 => \REG[362]\, 
        REG_362 => \REG[363]\, REG_363 => \REG[364]\, REG_364 => 
        \REG[365]\, REG_365 => \REG[366]\, REG_366 => \REG[367]\, 
        REG_367 => \REG[368]\, REG_368 => \REG[369]\, REG_369 => 
        \REG[370]\, REG_370 => \REG[371]\, REG_371 => \REG[372]\, 
        REG_372 => \REG[373]\, REG_373 => \REG[374]\, REG_374 => 
        \REG[375]\, REG_375 => \REG[376]\, REG_408 => \REG[409]\, 
        REG_480 => \REG[481]\, REG_80 => \REG[81]\, REG_81 => 
        \REG[82]\, REG_82 => \REG[83]\, REG_83 => \REG[84]\, 
        REG_84 => \REG[85]\, REG_85 => \REG[86]\, REG_86 => 
        \REG[87]\, REG_87 => \REG[88]\, REG_88 => \REG[89]\, 
        REG_89 => \REG[90]\, REG_90 => \REG[91]\, REG_96 => 
        \REG[97]\, REG_97 => \REG[98]\, REG_98 => \REG[99]\, 
        REG_99 => \REG[100]\, REG_100 => \REG[101]\, REG_101 => 
        \REG[102]\, REG_102 => \REG[103]\, REG_103 => \REG[104]\, 
        REG_376 => \REG[377]\, REG_120 => \REG[121]\, REG_152 => 
        \REG[153]\, REG_232 => \REG[233]\, REG_248 => \REG[249]\, 
        REG_168 => \REG[169]\, REG_184 => \REG[185]\, REG_104 => 
        \REG[105]\, REG_136 => \REG[137]\, REG_31 => \REG[32]\, 
        REG_47 => \REG[48]\, REG_440 => \REG[441]\, REG_456 => 
        \REG[457]\, REG_441 => \REG[442]\, REG_457 => \REG[458]\, 
        REG_473 => \REG[474]\, REG_121 => \REG[122]\, REG_153 => 
        \REG[154]\, REG_233 => \REG[234]\, REG_249 => \REG[250]\, 
        REG_169 => \REG[170]\, REG_185 => \REG[186]\, REG_105 => 
        \REG[106]\, REG_137 => \REG[138]\, REG_32 => \REG[33]\, 
        REG_16 => \REG[17]\, REG_48 => \REG[49]\, REG_377 => 
        \REG[378]\, REG_409 => \REG[410]\, REG_442 => \REG[443]\, 
        REG_458 => \REG[459]\, REG_474 => \REG[475]\, REG_378 => 
        \REG[379]\, REG_410 => \REG[411]\, REG_154 => \REG[155]\, 
        REG_170 => \REG[171]\, REG_122 => \REG[123]\, REG_250 => 
        \REG[251]\, REG_138 => \REG[139]\, REG_186 => \REG[187]\, 
        REG_234 => \REG[235]\, REG_33 => \REG[34]\, REG_49 => 
        \REG[50]\, REG_34 => \REG[35]\, REG_50 => \REG[51]\, 
        REG_155 => \REG[156]\, REG_171 => \REG[172]\, REG_251 => 
        \REG[252]\, REG_139 => \REG[140]\, REG_187 => \REG[188]\, 
        REG_235 => \REG[236]\, REG_443 => \REG[444]\, REG_459 => 
        \REG[460]\, REG_379 => \REG[380]\, REG_411 => \REG[412]\, 
        REG_475 => \REG[476]\, REG_51 => \REG[52]\, REG_35 => 
        \REG[36]\, REG_19 => \REG[20]\, REG_156 => \REG[157]\, 
        REG_172 => \REG[173]\, REG_252 => \REG[253]\, REG_140 => 
        \REG[141]\, REG_188 => \REG[189]\, REG_236 => \REG[237]\, 
        REG_332 => \REG[333]\, REG_444 => \REG[445]\, REG_460 => 
        \REG[461]\, REG_380 => \REG[381]\, REG_412 => \REG[413]\, 
        REG_476 => \REG[477]\, REG_445 => \REG[446]\, REG_461 => 
        \REG[462]\, REG_413 => \REG[414]\, REG_381 => \REG[382]\, 
        REG_52 => \REG[53]\, REG_36 => \REG[37]\, REG_157 => 
        \REG[158]\, REG_173 => \REG[174]\, REG_253 => \REG[254]\, 
        REG_141 => \REG[142]\, REG_189 => \REG[190]\, REG_237 => 
        \REG[238]\, REG_333 => \REG[334]\, REG_477 => \REG[478]\, 
        REG_462 => \REG[463]\, REG_478 => \REG[479]\, REG_382 => 
        \REG[383]\, REG_414 => \REG[415]\, REG_37 => \REG[38]\, 
        REG_5 => \REG[6]\, REG_53 => \REG[54]\, REG_158 => 
        \REG[159]\, REG_174 => \REG[175]\, REG_254 => \REG[255]\, 
        REG_142 => \REG[143]\, REG_190 => \REG[191]\, REG_238 => 
        \REG[239]\, REG_334 => \REG[335]\, REG_463 => \REG[464]\, 
        REG_383 => \REG[384]\, REG_415 => \REG[416]\, REG_54 => 
        \REG[55]\, REG_38 => \REG[39]\, REG_159 => \REG[160]\, 
        REG_175 => \REG[176]\, REG_255 => \REG[256]\, REG_143 => 
        \REG[144]\, REG_191 => \REG[192]\, REG_239 => \REG[240]\, 
        REG_479 => \REG[480]\, REG_464 => \REG[465]\, REG_416 => 
        \REG[417]\, REG_39 => \REG[40]\, REG_7 => \REG[8]\, 
        REG_55 => \REG[56]\, REG_128 => \REG[129]\, REG_160 => 
        \REG[161]\, REG_240 => \REG[241]\, REG_256 => \REG[257]\, 
        REG_176 => \REG[177]\, REG_192 => \REG[193]\, REG_112 => 
        \REG[113]\, REG_144 => \REG[145]\, REG_465 => \REG[466]\, 
        REG_56 => \REG[57]\, REG_40 => \REG[41]\, REG_161 => 
        \REG[162]\, REG_177 => \REG[178]\, REG_129 => \REG[130]\, 
        REG_257 => \REG[258]\, REG_113 => \REG[114]\, REG_193 => 
        \REG[194]\, REG_241 => \REG[242]\, REG_417 => \REG[418]\, 
        REG_466 => \REG[467]\, REG_57 => \REG[58]\, REG_41 => 
        \REG[42]\, REG_162 => \REG[163]\, REG_178 => \REG[179]\, 
        REG_130 => \REG[131]\, REG_258 => \REG[259]\, REG_114 => 
        \REG[115]\, REG_194 => \REG[195]\, REG_242 => \REG[243]\, 
        REG_418 => \REG[419]\, REG_467 => \REG[468]\, REG_42 => 
        \REG[43]\, REG_58 => \REG[59]\, REG_163 => \REG[164]\, 
        REG_179 => \REG[180]\, REG_131 => \REG[132]\, REG_259 => 
        \REG[260]\, REG_115 => \REG[116]\, REG_195 => \REG[196]\, 
        REG_243 => \REG[244]\, REG_419 => \REG[420]\, REG_468 => 
        \REG[469]\, REG_43 => \REG[44]\, REG_59 => \REG[60]\, 
        REG_164 => \REG[165]\, REG_180 => \REG[181]\, REG_132 => 
        \REG[133]\, REG_260 => \REG[261]\, REG_116 => \REG[117]\, 
        REG_196 => \REG[197]\, REG_244 => \REG[245]\, REG_420 => 
        \REG[421]\, REG_469 => \REG[470]\, REG_60 => \REG[61]\, 
        REG_44 => \REG[45]\, REG_165 => \REG[166]\, REG_181 => 
        \REG[182]\, REG_133 => \REG[134]\, REG_261 => \REG[262]\, 
        REG_117 => \REG[118]\, REG_197 => \REG[198]\, REG_245 => 
        \REG[246]\, REG_421 => \REG[422]\, REG_470 => \REG[471]\, 
        REG_61 => \REG[62]\, REG_45 => \REG[46]\, REG_166 => 
        \REG[167]\, REG_182 => \REG[183]\, REG_134 => \REG[135]\, 
        REG_262 => \REG[263]\, REG_118 => \REG[119]\, REG_198 => 
        \REG[199]\, REG_246 => \REG[247]\, REG_422 => \REG[423]\, 
        REG_455 => \REG[456]\, REG_471 => \REG[472]\, REG_423 => 
        \REG[424]\, REG_46 => \REG[47]\, REG_62 => \REG[63]\, 
        REG_167 => \REG[168]\, REG_183 => \REG[184]\, REG_135 => 
        \REG[136]\, REG_263 => \REG[264]\, REG_119 => \REG[120]\, 
        REG_199 => \REG[200]\, REG_247 => \REG[248]\, REG_63 => 
        \REG[64]\, REG_424 => \REG[425]\, REG_64 => \REG[65]\, 
        REG_425 => \REG[426]\, REG_65 => \REG[66]\, REG_426 => 
        \REG[427]\, REG_66 => \REG[67]\, REG_427 => \REG[428]\, 
        REG_67 => \REG[68]\, REG_428 => \REG[429]\, REG_68 => 
        \REG[69]\, REG_429 => \REG[430]\, REG_69 => \REG[70]\, 
        REG_430 => \REG[431]\, REG_70 => \REG[71]\, REG_431 => 
        \REG[432]\, REG_71 => \REG[72]\, REG_432 => \REG[433]\, 
        REG_72 => \REG[73]\, REG_433 => \REG[434]\, REG_73 => 
        \REG[74]\, REG_434 => \REG[435]\, REG_74 => \REG[75]\, 
        REG_435 => \REG[436]\, REG_75 => \REG[76]\, REG_436 => 
        \REG[437]\, REG_76 => \REG[77]\, REG_437 => \REG[438]\, 
        REG_77 => \REG[78]\, REG_438 => \REG[439]\, REG_78 => 
        \REG[79]\, REG_439 => \REG[440]\, REG_4 => \REG[5]\, 
        REG_79 => \REG[80]\, TST_c_c(3) => \TST_c_c[3]\, TST_c_4
         => \TST_c[4]\, TST_c_0 => \TST_c[0]\, TST_c_5 => 
        \TST_c[5]\, TST_c_2 => \TST_c[2]\, TST_c_1 => \TST_c[1]\, 
        REG_i_0_116 => \REG_i_0[121]\, REG_i_0_0 => \REG_i_0[5]\, 
        REG_i_0_75 => \REG_i_0[80]\, REG_i_0_260 => 
        \REG_i_0[265]\, REG_i_0_261 => \REG_i_0[266]\, 
        REG_i_0_275 => \REG_i_0[280]\, REG_i_0_276 => 
        \REG_i_0[281]\, REG_i_0_277 => \REG_i_0[282]\, 
        REG_i_0_278 => \REG_i_0[283]\, REG_i_0_279 => 
        \REG_i_0[284]\, REG_i_0_280 => \REG_i_0[285]\, 
        REG_i_0_281 => \REG_i_0[286]\, REG_i_0_282 => 
        \REG_i_0[287]\, REG_i_0_283 => \REG_i_0[288]\, 
        REG_i_0_284 => \REG_i_0[289]\, REG_i_0_285 => 
        \REG_i_0[290]\, REG_i_0_286 => \REG_i_0[291]\, 
        REG_i_0_287 => \REG_i_0[292]\, REG_i_0_288 => 
        \REG_i_0[293]\, REG_i_0_289 => \REG_i_0[294]\, 
        REG_i_0_290 => \REG_i_0[295]\, REG_i_0_291 => 
        \REG_i_0[296]\, REG_i_0_393 => \REG_i_0[398]\, 
        REG_i_0_391 => \REG_i_0[396]\, REG_i_0_395 => 
        \REG_i_0[400]\, REG_i_0_388 => \REG_i_0[393]\, 
        REG_i_0_389 => \REG_i_0[394]\, REG_i_0_390 => 
        \REG_i_0[395]\, REG_i_0_392 => \REG_i_0[397]\, 
        REG_i_0_394 => \REG_i_0[399]\, REG_0(127) => \REG_0[127]\, 
        REG_0(126) => \REG_0[126]\, REG_0(125) => \REG_0[125]\, 
        REG_0(124) => \REG_0[124]\, HWRES_c_16 => HWRES_c_16, 
        HWRES_c_15 => HWRES_c_15, CLEAR_22 => CLEAR_22, CLEAR_21
         => CLEAR_21, CLEAR_25 => CLEAR_25, CLEAR_24 => CLEAR_24, 
        CLEAR_23 => CLEAR_23, CLEAR_27 => CLEAR_27, CLEAR_26 => 
        CLEAR_26, HWRES_c_18 => HWRES_c_18, HWRES_c_22 => 
        HWRES_c_22, CLEAR_28 => CLEAR_28, CLEAR => CLEAR, 
        HWRES_c_17 => HWRES_c_17, HWRES_c_21 => HWRES_c_21, 
        HWRES_c_12 => HWRES_c_12, HWRES_c_23 => HWRES_c_23, RAMRD
         => RAMRD, HWRES_c_19 => HWRES_c_19, OR_RACK => OR_RACK, 
        HWRES_c_14 => HWRES_c_14, OR_RREQ => OR_RREQ, HWRES_c_20
         => HWRES_c_20, EF => EF, CLEAR_20 => CLEAR_20, ASB_c => 
        ASB_c, un5_noe16ri_0_0 => un5_noe16ri_0_0, 
        un7_noe32ri_0_0 => un7_noe32ri_0_0, WRITEB_c => WRITEB_c, 
        nLBAS_c => nLBAS_c, LB_nOE => \I2.LB_nOE\, LWORDB_in => 
        LWORDB_in, MYBERR_c => MYBERR_c, IACKB_c => IACKB_c, 
        nLBRDY_c => nLBRDY_c, FWIMG2LOAD => FWIMG2LOAD, NLBLAST_c
         => NLBLAST_c, NLBRD_c => NLBRD_c, NLBCLR_c => NLBCLR_c, 
        EVREAD => EVREAD, NRDMEB => NRDMEB, DTEST_FIFO => 
        DTEST_FIFO, RUN_c => RUN_c, N_2052 => \I2.N_2052\, d_m7
         => \d_m7\, EV_RES_c => EV_RES_c, L0_c_c => L0_c_c, 
        L1A_c_c => L1A_c_c, L1R_c_c => L1R_c_c, L2A_c_c => 
        L2A_c_c, L2R_c_c => L2R_c_c, LOS_c_c => LOS_c_c, N_441
         => \I2.N_441\, SPULSE0_c_c => SPULSE0_c_c, SPULSE1_c_c
         => SPULSE1_c_c, SPULSE2_c_c => SPULSE2_c_c, DS1B_c => 
        DS1B_c, DS0B_c => DS0B_c, N_500 => \I2.N_500\, NDTKIN_c
         => NDTKIN_c, NOE16W_c => NOE16W_c, NOE32W_c => NOE32W_c, 
        NOEAD_c => NOEAD_c, NSELCLK_c => NSELCLK_c, NSELCLK_c_i_0
         => NSELCLK_c_i_0, CLEAR_0 => CLEAR_0, EVRDY_c => EVRDY_c, 
        HWRES_c_1 => HWRES_c_1, NOEAD_c_i_0 => NOEAD_c_i_0, 
        N_2613_0 => \I2.N_2613_0\, RUN_c_0 => RUN_c_0, HWRES_c_0
         => HWRES_c_0, NOEAD_c_0 => NOEAD_c_0, NOEAD_c_1 => 
        NOEAD_c_1, HWRES_c_22_0 => HWRES_c_22_0, ALICLK_c => 
        ALICLK_c, un7_noe32ri_0 => \I2.un7_noe32ri_0\, 
        un5_noe16ri_0 => \I2.un5_noe16ri_0\, WDOGTO => WDOGTO, 
        HWRES_c_0_6 => HWRES_c_0_6, HWRES_c_0_5 => HWRES_c_0_5, 
        HWRES_c_0_4 => HWRES_c_0_4, HWRES_c_0_3 => HWRES_c_0_3, 
        HWRES_c_23_0 => HWRES_c_23_0, HWRES_c_21_0 => 
        HWRES_c_21_0, HWRES_c_13_0 => HWRES_c_13_0, HWRES_c_0_0
         => HWRES_c_0_0, NOEAD_c_0_0 => NOEAD_c_0_0, HWRES_c_13
         => HWRES_c_13, CLK_c_c => CLK_c_c, RUN_c_0_0 => 
        RUN_c_0_0, HWRES_c_0_6_0 => HWRES_c_0_6_0);
    
    \AMB_pad[5]\ : IB33
      port map(PAD => AMB(5), Y => \AMB_c[5]\);
    
    \AE_PDL_pad[32]\ : OB33PH
      port map(PAD => AE_PDL(32), A => \AE_PDL_c[32]\);
    
    \LB_pad[2]\ : IOB33PH
      port map(PAD => LB(2), A => \I2.LB_i[2]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[2]\);
    
    L0_pad : IB33
      port map(PAD => L0, Y => L0_c_c);
    
    \SP_PDL_pad[34]\ : IOB33PH
      port map(PAD => SP_PDL(34), A => \I3.P0[34]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[34]\);
    
    NLBCS_pad : OB33PH
      port map(PAD => NLBCS, A => \GND\);
    
    \LBSP_pad[17]\ : IOB33PH
      port map(PAD => LBSP(17), A => \REG[362]\, EN => 
        \REG_i_0[282]\, Y => \LBSP_in[17]\);
    
    d_m7 : NOR2FT
      port map(A => d_N_7, B => \I2.N_2613_0\, Y => \d_m7\);
    
    \TST_pad[12]\ : OTB33PH
      port map(PAD => TST(12), A => \GND\, EN => \GND\);
    
    \SP_PDL_pad[36]\ : IOB33PH
      port map(PAD => SP_PDL(36), A => \I3.P0[36]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[36]\);
    
    I6 : CROM
      port map(CROMWDT(7) => \CROMWDT[7]\, CROMWDT(6) => 
        \CROMWDT[6]\, CROMWDT(5) => \CROMWDT[5]\, CROMWDT(4) => 
        \CROMWDT[4]\, CROMWDT(3) => \CROMWDT[3]\, CROMWDT(2) => 
        \CROMWDT[2]\, CROMWDT(1) => \CROMWDT[1]\, CROMWDT(0) => 
        \CROMWDT[0]\, RAMAD_VME(8) => \RAMAD_VME[8]\, 
        RAMAD_VME(7) => \RAMAD_VME[7]\, RAMAD_VME(6) => 
        \RAMAD_VME[6]\, RAMAD_VME(5) => \RAMAD_VME[5]\, 
        RAMAD_VME(4) => \RAMAD_VME[4]\, RAMAD_VME(3) => 
        \RAMAD_VME[3]\, RAMAD_VME(2) => \RAMAD_VME[2]\, 
        RAMAD_VME(1) => \RAMAD_VME[1]\, RAMAD_VME(0) => 
        \RAMAD_VME[0]\, CROMWAD(8) => \CROMWAD[8]\, CROMWAD(7)
         => \CROMWAD[7]\, CROMWAD(6) => \CROMWAD[6]\, CROMWAD(5)
         => \CROMWAD[5]\, CROMWAD(4) => \CROMWAD[4]\, CROMWAD(3)
         => \CROMWAD[3]\, CROMWAD(2) => \CROMWAD[2]\, CROMWAD(1)
         => \CROMWAD[1]\, CROMWAD(0) => \CROMWAD[0]\, RAMDT(7)
         => \RAMDT[7]\, RAMDT(6) => \RAMDT[6]\, RAMDT(5) => 
        \RAMDT[5]\, RAMDT(4) => \RAMDT[4]\, RAMDT(3) => 
        \RAMDT[3]\, RAMDT(2) => \RAMDT[2]\, RAMDT(1) => 
        \RAMDT[1]\, RAMDT(0) => \RAMDT[0]\, WRCROM => WRCROM, 
        RAMRD => RAMRD, CLK_c_c => CLK_c_c);
    
    I_9 : INV
      port map(A => \I5.sstate_0[2]\, Y => \I5.sstate_0_i_0[2]\);
    
    \VDB_pad_0[12]\ : BFR
      port map(A => \VDB_in[12]\, Y => \VDB_in_0[12]\);
    
    \LBSP_pad[11]\ : OB33PH
      port map(PAD => LBSP(11), A => SPULSE0_c_c);
    
    d_m4 : MUX2H
      port map(A => d_N_3, B => \I2.N_2052\, S => \I2.N_441\, Y
         => d_N_5);
    
    I0 : RESET_MOD
      port map(TICK_2_d0 => \TICK[2]\, TICK_1_d0 => \TICK[1]\, 
        TICK_0_d0 => \TICK[0]\, LBSP_c(2) => \LBSP_c[2]\, 
        PULSE(1) => \PULSE[1]\, LBSP_c_0(2) => \LBSP_c_0[2]\, 
        LBSP_c_1(2) => \LBSP_c_1[2]\, TST_c(15) => \TST_c[15]\, 
        TST_c(14) => \TST_c[14]\, TST_c(13) => \TST_c[13]\, 
        TICK_0_2 => \TICK_0[2]\, TICK_0_0 => \TICK_0[0]\, 
        TICK_1(0) => \TICK_1[0]\, TICK_2(0) => \TICK_2[0]\, 
        REG_464 => \REG[472]\, REG_463 => \REG[471]\, REG_462 => 
        \REG[470]\, REG_461 => \REG[469]\, REG_460 => \REG[468]\, 
        REG_459 => \REG[467]\, REG_458 => \REG[466]\, REG_456 => 
        \REG[464]\, REG_455 => \REG[463]\, REG_454 => \REG[462]\, 
        REG_453 => \REG[461]\, REG_451 => \REG[459]\, REG_457 => 
        \REG[465]\, REG_452 => \REG[460]\, REG_449 => \REG[457]\, 
        REG_450 => \REG[458]\, REG_0 => \REG[8]\, PON_LOAD_i => 
        PON_LOAD_i, EV_RES_c => EV_RES_c, RUN_c => RUN_c, 
        LOAD_RES => LOAD_RES, CLEAR => CLEAR, BNCRES_c => 
        BNCRES_c, EVRES_c => EVRES_c, WDOGTO => WDOGTO, HWRES_c
         => HWRES_c, HWRES_c_i_0 => HWRES_c_i_0, CLEAR_i_0 => 
        CLEAR_i_0, RUN_c_0 => RUN_c_0, ALICLK_c => ALICLK_c, 
        HWRES_c_0 => HWRES_c_0, HWRES_c_1 => HWRES_c_1, HWRES_c_2
         => HWRES_c_2, HWRES_c_3 => HWRES_c_3, HWRES_c_4 => 
        HWRES_c_4, HWRES_c_5 => HWRES_c_5, NPWON_c => NPWON_c, 
        HWRES_c_6 => HWRES_c_6, HWRES_c_7 => HWRES_c_7, HWRES_c_8
         => HWRES_c_8, HWRES_c_9 => HWRES_c_9, HWRES_c_10 => 
        HWRES_c_10, HWRES_c_11 => HWRES_c_11, HWRES_c_12 => 
        HWRES_c_12, HWRES_c_13 => HWRES_c_13, HWRES_c_14 => 
        HWRES_c_14, HWRES_c_15 => HWRES_c_15, HWRES_c_16 => 
        HWRES_c_16, HWRES_c_17 => HWRES_c_17, HWRES_c_18 => 
        HWRES_c_18, HWRES_c_19 => HWRES_c_19, HWRES_c_20 => 
        HWRES_c_20, HWRES_c_21 => HWRES_c_21, HWRES_c_22 => 
        HWRES_c_22, HWRES_c_23 => HWRES_c_23, HWRES_c_24 => 
        HWRES_c_24, HWRES_c_25 => HWRES_c_25, HWRES_c_26 => 
        HWRES_c_26, HWRES_c_27 => HWRES_c_27, HWRES_c_28 => 
        HWRES_c_28, HWRES_c_29 => HWRES_c_29, HWRES_c_30 => 
        HWRES_c_30, HWRES_c_31 => HWRES_c_31, HWRES_c_32 => 
        HWRES_c_32, HWRES_c_33 => HWRES_c_33, HWRES_c_34 => 
        HWRES_c_34, HWRES_c_35 => HWRES_c_35, HWRES_c_36 => 
        HWRES_c_36, CLEAR_0 => CLEAR_0, CLEAR_2 => CLEAR_2, 
        CLEAR_3 => CLEAR_3, CLEAR_4 => CLEAR_4, CLEAR_5 => 
        CLEAR_5, CLEAR_6 => CLEAR_6, CLEAR_7 => CLEAR_7, CLEAR_8
         => CLEAR_8, LOAD_RES_2 => LOAD_RES_2, CLEAR_9 => CLEAR_9, 
        CLEAR_10 => CLEAR_10, CLEAR_11 => CLEAR_11, CLEAR_12 => 
        CLEAR_12, CLEAR_13 => CLEAR_13, CLEAR_14 => CLEAR_14, 
        CLEAR_15 => CLEAR_15, CLEAR_16 => CLEAR_16, CLEAR_17 => 
        CLEAR_17, CLEAR_18 => CLEAR_18, LOAD_RES_1 => LOAD_RES_1, 
        CLEAR_19 => CLEAR_19, CLEAR_20 => CLEAR_20, CLEAR_21 => 
        CLEAR_21, CLEAR_22 => CLEAR_22, CLEAR_23 => CLEAR_23, 
        CLEAR_24 => CLEAR_24, CLEAR_25 => CLEAR_25, CLEAR_26 => 
        CLEAR_26, CLEAR_27 => CLEAR_27, LOAD_RES_0 => LOAD_RES_0, 
        CLEAR_28 => CLEAR_28, HWRES_c_36_0 => HWRES_c_36_0, 
        HWRES_c_32_0 => HWRES_c_32_0, NPWON_c_1 => NPWON_c_1, 
        HWRES_c_23_0 => HWRES_c_23_0, HWRES_c_22_0 => 
        HWRES_c_22_0, HWRES_c_21_0 => HWRES_c_21_0, HWRES_c_13_0
         => HWRES_c_13_0, HWRES_c_10_0 => HWRES_c_10_0, 
        HWRES_c_0_0 => HWRES_c_0_0, HWRES_c_0_2 => HWRES_c_0_2, 
        HWRES_c_0_3 => HWRES_c_0_3, HWRES_c_0_4 => HWRES_c_0_4, 
        HWRES_c_0_5 => HWRES_c_0_5, HWRES_c_0_6 => HWRES_c_0_6, 
        RUN_c_0_0 => RUN_c_0_0, NLBCLR_c => NLBCLR_c, SYSRESB_c
         => SYSRESB_c, CLK_c_c => CLK_c_c, NPWON_c_2 => NPWON_c_2, 
        HWRES_c_27_0 => HWRES_c_27_0, NPWON_c_3 => NPWON_c_3, 
        HWRES_c_7_0 => HWRES_c_7_0, NPWON_c_0 => NPWON_c_0, 
        HWRES_c_0_6_0 => HWRES_c_0_6_0);
    
    IACKOUTB_pad : OB33PH
      port map(PAD => IACKOUTB, A => \VCC\);
    
    I5 : SPI_INTERF
      port map(CROMWDT(7) => \CROMWDT[7]\, CROMWDT(6) => 
        \CROMWDT[6]\, CROMWDT(5) => \CROMWDT[5]\, CROMWDT(4) => 
        \CROMWDT[4]\, CROMWDT(3) => \CROMWDT[3]\, CROMWDT(2) => 
        \CROMWDT[2]\, CROMWDT(1) => \CROMWDT[1]\, CROMWDT(0) => 
        \CROMWDT[0]\, DACCFG_WDT(13) => \DACCFG_WDT[13]\, 
        DACCFG_WDT(12) => \DACCFG_WDT[12]\, DACCFG_WDT(11) => 
        \DACCFG_WDT[11]\, DACCFG_WDT(10) => \DACCFG_WDT[10]\, 
        DACCFG_WDT(9) => \DACCFG_WDT[9]\, DACCFG_WDT(8) => 
        \DACCFG_WDT[8]\, DACCFG_WDT(7) => \DACCFG_WDT[7]\, 
        DACCFG_WDT(6) => \DACCFG_WDT[6]\, DACCFG_WDT(5) => 
        \DACCFG_WDT[5]\, DACCFG_WDT(4) => \DACCFG_WDT[4]\, 
        TICK(1) => \TICK[1]\, FBOUT(7) => \FBOUT[7]\, FBOUT(6)
         => \FBOUT[6]\, FBOUT(5) => \FBOUT[5]\, FBOUT(4) => 
        \FBOUT[4]\, FBOUT(3) => \FBOUT[3]\, FBOUT(2) => 
        \FBOUT[2]\, FBOUT(1) => \FBOUT[1]\, FBOUT(0) => 
        \FBOUT[0]\, REG_i_0(80) => \REG_i_0[80]\, REG_400 => 
        \REG[480]\, REG_398 => \REG[478]\, REG_396 => \REG[476]\, 
        REG_393 => \REG[473]\, REG_0 => \REG[80]\, REG_1 => 
        \REG[81]\, REG_2 => \REG[82]\, REG_3 => \REG[83]\, REG_4
         => \REG[84]\, REG_5 => \REG[85]\, REG_6 => \REG[86]\, 
        REG_7 => \REG[87]\, REG_8 => \REG[88]\, REG_399 => 
        \REG[479]\, REG_395 => \REG[475]\, REG_397 => \REG[477]\, 
        REG_394 => \REG[474]\, CROMWAD(8) => \CROMWAD[8]\, 
        CROMWAD(7) => \CROMWAD[7]\, CROMWAD(6) => \CROMWAD[6]\, 
        CROMWAD(5) => \CROMWAD[5]\, CROMWAD(4) => \CROMWAD[4]\, 
        CROMWAD(3) => \CROMWAD[3]\, CROMWAD(2) => \CROMWAD[2]\, 
        CROMWAD(1) => \CROMWAD[1]\, CROMWAD(0) => \CROMWAD[0]\, 
        sstate_0_2 => \I5.sstate_0[2]\, PULSE_6 => \PULSE[6]\, 
        PULSE_0 => \PULSE[0]\, PULSE_10 => \PULSE[10]\, 
        sstate_0_i_0(2) => \I5.sstate_0_i_0[2]\, HWRES_c_30 => 
        HWRES_c_30, HWRES_c_23_0 => HWRES_c_23_0, HWRES_c_28 => 
        HWRES_c_28, HWRES_c_31 => HWRES_c_31, HWRES_c_24 => 
        HWRES_c_24, HWRES_c_25 => HWRES_c_25, DACCFG_nWR => 
        DACCFG_nWR, PDLCFG_nWR => PDLCFG_nWR, HWRES_c_32 => 
        HWRES_c_32, WRCROM => WRCROM, HWRES_c_26 => HWRES_c_26, 
        HWRES_c_27 => HWRES_c_27, NCYC_RELOAD_in => 
        NCYC_RELOAD_in, HWRES_c_29 => HWRES_c_29, un1_drive_spi
         => un1_drive_spi, F_SO_c => F_SO_c, LOAD_RES => LOAD_RES, 
        DRIVE_RELOAD => \I5.DRIVE_RELOAD\, ISCK => \I5.ISCK\, 
        FWIMG2LOAD => FWIMG2LOAD, ISI => \I5.ISI\, FCS_c => FCS_c, 
        PON_LOAD_i => PON_LOAD_i, HWRES_c_32_0 => HWRES_c_32_0, 
        LOAD_RES_0 => LOAD_RES_0, LOAD_RES_1 => LOAD_RES_1, 
        LOAD_RES_2 => LOAD_RES_2, CLK_c_c => CLK_c_c, 
        HWRES_c_27_0 => HWRES_c_27_0, LOAD_RES_3 => LOAD_RES_3);
    
    \SP_PDL_pad[14]\ : IOB33PH
      port map(PAD => SP_PDL(14), A => \I3.P0[14]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[14]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \AE_PDL_pad[40]\ : OB33PH
      port map(PAD => AE_PDL(40), A => \AE_PDL_c[40]\);
    
    \AE_PDL_pad[21]\ : OB33PH
      port map(PAD => AE_PDL(21), A => \AE_PDL_c[21]\);
    
    \TST_pad[14]\ : OB33PH
      port map(PAD => TST(14), A => \TST_c[14]\);
    
    \SP_PDL_pad[16]\ : IOB33PH
      port map(PAD => SP_PDL(16), A => \I3.P0[16]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[16]\);
    
    \LB_pad[31]\ : IOB33PH
      port map(PAD => LB(31), A => \I2.LB_i[31]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[31]\);
    
    \LBSP_pad[2]\ : OB33PH
      port map(PAD => LBSP(2), A => \LBSP_c[2]\);
    
    SPULSE0_pad : IB33
      port map(PAD => SPULSE0, Y => SPULSE0_c_c);
    
    \TST_pad[1]\ : OB33PH
      port map(PAD => TST(1), A => \TST_c[1]\);
    
    \VDB_pad[4]\ : IOB33PH
      port map(PAD => VDB(4), A => \I2.VDBm[4]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[4]\);
    
    \SP_PDL_pad[29]\ : IOB33PH
      port map(PAD => SP_PDL(29), A => \I3.P0[29]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[29]\);
    
    SDA0_pad : IOB33PH
      port map(PAD => SDA0, A => \I1.SDAout_del2\, EN => 
        un1_sdaa_0_a3, Y => SDA0_in);
    
    \LBSP_pad[16]\ : IOB33PH
      port map(PAD => LBSP(16), A => \REG[361]\, EN => 
        \REG_i_0[281]\, Y => \LBSP_in[16]\);
    
    \VDB_pad[11]\ : IOB33PH
      port map(PAD => VDB(11), A => \VDBm_i_m2[11]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[11]\);
    
    \SYNC_pad[7]\ : OB33PH
      port map(PAD => SYNC(7), A => \SYNC_c[7]\);
    
    \SP_PDL_pad[41]\ : IOB33PH
      port map(PAD => SP_PDL(41), A => \I3.P0[41]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[41]\);
    
    \AE_PDL_pad[7]\ : OB33PH
      port map(PAD => AE_PDL(7), A => \AE_PDL_c[7]\);
    
    \LBSP_pad[13]\ : OB33PH
      port map(PAD => LBSP(13), A => SPULSE2_c_c);
    
    \LBSP_pad[0]\ : IOB33PH
      port map(PAD => LBSP(0), A => \REG[345]\, EN => 
        \REG_i_0[265]\, Y => \LBSP_in[0]\);
    
    I10 : ROC32
      port map(DPR(31) => \DPR[31]\, DPR(30) => \DPR[30]\, 
        DPR(29) => \DPR[29]\, DPR(28) => \DPR[28]\, DPR(27) => 
        \DPR[27]\, DPR(26) => \DPR[26]\, DPR(25) => \DPR[25]\, 
        DPR(24) => \DPR[24]\, DPR(23) => \DPR[23]\, DPR(22) => 
        \DPR[22]\, DPR(21) => \DPR[21]\, DPR(20) => \DPR[20]\, 
        DPR(19) => \DPR[19]\, DPR(18) => \DPR[18]\, DPR(17) => 
        \DPR[17]\, DPR(16) => \DPR[16]\, DPR(15) => \DPR[15]\, 
        DPR(14) => \DPR[14]\, DPR(13) => \DPR[13]\, DPR(12) => 
        \DPR[12]\, DPR(11) => \DPR[11]\, DPR(10) => \DPR[10]\, 
        DPR(9) => \DPR[9]\, DPR(8) => \DPR[8]\, DPR(7) => 
        \DPR[7]\, DPR(6) => \DPR[6]\, DPR(5) => \DPR[5]\, DPR(4)
         => \DPR[4]\, DPR(3) => \DPR[3]\, DPR(2) => \DPR[2]\, 
        DPR(1) => \DPR[1]\, DPR(0) => \DPR[0]\, un2_evread_0 => 
        \I10.un2_evread[14]\, CHANNEL(2) => \CHANNEL[2]\, 
        CHANNEL(1) => \CHANNEL[1]\, CHANNEL(0) => \CHANNEL[0]\, 
        CHIP_ADDR(2) => \CHIP_ADDR[2]\, CHIP_ADDR(1) => 
        \CHIP_ADDR[1]\, CHIP_ADDR(0) => \CHIP_ADDR[0]\, 
        I2C_RDATA(9) => \I2C_RDATA[9]\, I2C_RDATA(8) => 
        \I2C_RDATA[8]\, I2C_RDATA(7) => \I2C_RDATA[7]\, 
        I2C_RDATA(6) => \I2C_RDATA[6]\, I2C_RDATA(5) => 
        \I2C_RDATA[5]\, I2C_RDATA(4) => \I2C_RDATA[4]\, 
        I2C_RDATA(3) => \I2C_RDATA[3]\, I2C_RDATA(2) => 
        \I2C_RDATA[2]\, I2C_RDATA(1) => \I2C_RDATA[1]\, 
        I2C_RDATA(0) => \I2C_RDATA[0]\, OR_RDATA(9) => 
        \OR_RDATA[9]\, OR_RDATA(8) => \OR_RDATA[8]\, OR_RDATA(7)
         => \OR_RDATA[7]\, OR_RDATA(6) => \OR_RDATA[6]\, 
        OR_RDATA(5) => \OR_RDATA[5]\, OR_RDATA(4) => 
        \OR_RDATA[4]\, OR_RDATA(3) => \OR_RDATA[3]\, OR_RDATA(2)
         => \OR_RDATA[2]\, OR_RDATA(1) => \OR_RDATA[1]\, 
        OR_RDATA(0) => \OR_RDATA[0]\, PDL_RDATA(7) => 
        \PDL_RDATA[7]\, PDL_RDATA(6) => \PDL_RDATA[6]\, 
        PDL_RDATA(5) => \PDL_RDATA[5]\, PDL_RDATA(4) => 
        \PDL_RDATA[4]\, PDL_RDATA(3) => \PDL_RDATA[3]\, 
        PDL_RDATA(2) => \PDL_RDATA[2]\, PDL_RDATA(1) => 
        \PDL_RDATA[1]\, PDL_RDATA(0) => \PDL_RDATA[0]\, GA_c(3)
         => \GA_c[3]\, GA_c(2) => \GA_c[2]\, GA_c(1) => \GA_c[1]\, 
        GA_c(0) => \GA_c[0]\, OR_RADDR(5) => \OR_RADDR[5]\, 
        OR_RADDR(4) => \OR_RADDR[4]\, OR_RADDR(3) => 
        \OR_RADDR[3]\, OR_RADDR(2) => \OR_RADDR[2]\, OR_RADDR(1)
         => \OR_RADDR[1]\, OR_RADDR(0) => \OR_RADDR[0]\, 
        PDL_RADDR(5) => \PDL_RADDR[5]\, PDL_RADDR(4) => 
        \PDL_RADDR[4]\, PDL_RADDR(3) => \PDL_RADDR[3]\, 
        PDL_RADDR(2) => \PDL_RADDR[2]\, PDL_RADDR(1) => 
        \PDL_RADDR[1]\, PDL_RADDR(0) => \PDL_RADDR[0]\, LBSP_c(2)
         => \LBSP_c[2]\, LBSP_c_1(2) => \LBSP_c_1[2]\, 
        LBSP_c_0(2) => \LBSP_c_0[2]\, PULSE(3) => \PULSE[3]\, 
        PULSE(2) => \PULSE[2]\, REG_i_0(5) => \REG_i_0[5]\, 
        REG_c(23) => \REG_c[23]\, REG_c(22) => \REG_c[22]\, 
        REG_c(21) => \REG_c[21]\, REG_330 => \REG[335]\, REG_329
         => \REG[334]\, REG_328 => \REG[333]\, REG_408 => 
        \REG[413]\, REG_410 => \REG[415]\, REG_432 => \REG[437]\, 
        REG_415 => \REG[420]\, REG_406 => \REG[411]\, REG_418 => 
        \REG[423]\, REG_421 => \REG[426]\, REG_430 => \REG[435]\, 
        REG_433 => \REG[438]\, REG_424 => \REG[429]\, REG_427 => 
        \REG[432]\, REG_416 => \REG[421]\, REG_419 => \REG[424]\, 
        REG_412 => \REG[417]\, REG_413 => \REG[418]\, REG_428 => 
        \REG[433]\, REG_431 => \REG[436]\, REG_422 => \REG[427]\, 
        REG_425 => \REG[430]\, REG_414 => \REG[419]\, REG_417 => 
        \REG[422]\, REG_409 => \REG[414]\, REG_411 => \REG[416]\, 
        REG_426 => \REG[431]\, REG_429 => \REG[434]\, REG_420 => 
        \REG[425]\, REG_423 => \REG[428]\, REG_407 => \REG[412]\, 
        REG_434 => \REG[439]\, REG_435 => \REG[440]\, REG_404 => 
        \REG[409]\, REG_405 => \REG[410]\, REG_43 => \REG[48]\, 
        REG_44 => \REG[49]\, REG_45 => \REG[50]\, REG_46 => 
        \REG[51]\, REG_47 => \REG[52]\, REG_48 => \REG[53]\, 
        REG_49 => \REG[54]\, REG_50 => \REG[55]\, REG_51 => 
        \REG[56]\, REG_52 => \REG[57]\, REG_53 => \REG[58]\, 
        REG_54 => \REG[59]\, REG_55 => \REG[60]\, REG_56 => 
        \REG[61]\, REG_57 => \REG[62]\, REG_58 => \REG[63]\, 
        REG_59 => \REG[64]\, REG_60 => \REG[65]\, REG_61 => 
        \REG[66]\, REG_62 => \REG[67]\, REG_63 => \REG[68]\, 
        REG_64 => \REG[69]\, REG_65 => \REG[70]\, REG_66 => 
        \REG[71]\, REG_67 => \REG[72]\, REG_68 => \REG[73]\, 
        REG_69 => \REG[74]\, REG_70 => \REG[75]\, REG_71 => 
        \REG[76]\, REG_72 => \REG[77]\, REG_73 => \REG[78]\, 
        REG_74 => \REG[79]\, REG_41 => \REG[46]\, REG_42 => 
        \REG[47]\, REG_0 => \REG[5]\, REG_15 => \REG[20]\, REG_27
         => \REG[32]\, REG_28 => \REG[33]\, REG_30 => \REG[35]\, 
        REG_29 => \REG[34]\, REG_39 => \REG[44]\, REG_37 => 
        \REG[42]\, REG_36 => \REG[41]\, REG_34 => \REG[39]\, 
        REG_33 => \REG[38]\, REG_38 => \REG[43]\, REG_35 => 
        \REG[40]\, REG_40 => \REG[45]\, REG_31 => \REG[36]\, 
        REG_32 => \REG[37]\, EF => EF, FF_c => \REG[17]\, NRDMEB
         => NRDMEB, CLEAR_i_0 => CLEAR_i_0, CLEAR_14 => CLEAR_14, 
        CLEAR_13 => CLEAR_13, CLEAR_4 => CLEAR_4, CLEAR_3 => 
        CLEAR_3, CLEAR_2 => CLEAR_2, CLEAR_8 => CLEAR_8, CLEAR_7
         => CLEAR_7, CLEAR_6 => CLEAR_6, CLEAR_11 => CLEAR_11, 
        CLEAR_10 => CLEAR_10, CLEAR_19 => CLEAR_19, CLEAR_9 => 
        CLEAR_9, CLEAR_18 => CLEAR_18, CLEAR_12 => CLEAR_12, 
        CLEAR_15 => CLEAR_15, CLEAR_20 => CLEAR_20, CLEAR_5 => 
        CLEAR_5, PDL_RACK => PDL_RACK, CLEAR_17 => CLEAR_17, 
        OR_RACK => OR_RACK, CLEAR_16 => CLEAR_16, L2R_c_c => 
        L2R_c_c, L2A_c_c => L2A_c_c, HWRES_c_12 => HWRES_c_12, 
        L1A_c_c => L1A_c_c, ALICLK_c => ALICLK_c, HWRES_c_11 => 
        HWRES_c_11, DTEST_FIFO => DTEST_FIFO, I2C_CHAIN => 
        I2C_CHAIN, PDL_RREQ => PDL_RREQ, I2C_RREQ => I2C_RREQ, 
        EVRDY_c => EVRDY_c, OR_RREQ => OR_RREQ, I2C_RACK => 
        I2C_RACK, EVNT_TRG => \I10.EVNT_TRG\, EVREAD => EVREAD, 
        CLK_c_c => CLK_c_c, CLEAR_0 => CLEAR_0, I_8 => \I_8\, 
        I_16 => \I_16\);
    
    \SYNC_pad[6]\ : OB33PH
      port map(PAD => SYNC(6), A => \SYNC_c[6]\);
    
    I1 : I2C_INTERF
      port map(PULSE(7) => \PULSE[7]\, I2C_RDATA(9) => 
        \I2C_RDATA[9]\, I2C_RDATA(8) => \I2C_RDATA[8]\, 
        I2C_RDATA(7) => \I2C_RDATA[7]\, I2C_RDATA(6) => 
        \I2C_RDATA[6]\, I2C_RDATA(5) => \I2C_RDATA[5]\, 
        I2C_RDATA(4) => \I2C_RDATA[4]\, I2C_RDATA(3) => 
        \I2C_RDATA[3]\, I2C_RDATA(2) => \I2C_RDATA[2]\, 
        I2C_RDATA(1) => \I2C_RDATA[1]\, I2C_RDATA(0) => 
        \I2C_RDATA[0]\, CHIP_ADDR(2) => \CHIP_ADDR[2]\, 
        CHIP_ADDR(1) => \CHIP_ADDR[1]\, CHIP_ADDR(0) => 
        \CHIP_ADDR[0]\, CHANNEL(2) => \CHANNEL[2]\, CHANNEL(1)
         => \CHANNEL[1]\, CHANNEL(0) => \CHANNEL[0]\, TICK(0) => 
        \TICK[0]\, TICK_2(0) => \TICK_2[0]\, REG_107 => 
        \REG[113]\, REG_108 => \REG[114]\, REG_109 => \REG[115]\, 
        REG_110 => \REG[116]\, REG_111 => \REG[117]\, REG_112 => 
        \REG[118]\, REG_113 => \REG[119]\, REG_114 => \REG[120]\, 
        REG_0 => \REG[6]\, REG_84 => \REG[90]\, REG_85 => 
        \REG[91]\, REG_91 => \REG[97]\, REG_92 => \REG[98]\, 
        REG_99 => \REG[105]\, REG_93 => \REG[99]\, REG_94 => 
        \REG[100]\, REG_95 => \REG[101]\, REG_96 => \REG[102]\, 
        REG_97 => \REG[103]\, REG_98 => \REG[104]\, REG_83 => 
        \REG[89]\, REG_100 => \REG[106]\, TICK_1(0) => 
        \TICK_1[0]\, TICK_0(0) => \TICK_0[0]\, HWRES_c_4 => 
        HWRES_c_4, HWRES_c_7 => HWRES_c_7, HWRES_c_11 => 
        HWRES_c_11, HWRES_c_10 => HWRES_c_10, HWRES_c_5 => 
        HWRES_c_5, HWRES_c_3 => HWRES_c_3, HWRES_c_6 => HWRES_c_6, 
        I2C_RACK => I2C_RACK, SDAout_del2 => \I1.SDAout_del2\, 
        HWRES_c_9 => HWRES_c_9, HWRES_c_8 => HWRES_c_8, 
        un1_sdaa_0_a3 => un1_sdaa_0_a3, RUN_c_0_0 => RUN_c_0_0, 
        RUN_c_0 => RUN_c_0, I2C_CHAIN => I2C_CHAIN, I2C_RREQ => 
        I2C_RREQ, SDA1_in => SDA1_in, SDA0_in => SDA0_in, 
        un1_sdab_i => un1_sdab_i, SCLB_i_a3 => SCLB_i_a3, 
        SCLA_i_a3 => SCLA_i_a3, HWRES_c_10_0 => HWRES_c_10_0, 
        CLK_c_c => CLK_c_c, HWRES_c_7_0 => HWRES_c_7_0);
    
    \VAD_pad[3]\ : IOB33PH
      port map(PAD => VAD(3), A => \I2.VADm[3]\, EN => NOEAD_c, Y
         => \VAD_in[3]\);
    
    I7 : ctrl
      port map(TST_c_c(3) => \TST_c_c[3]\, PULSE(2) => \PULSE[2]\, 
        TICK_0(2) => \TICK_0[2]\, REG_15 => \REG[456]\, REG_0 => 
        \REG[441]\, REG_1 => \REG[442]\, REG_2 => \REG[443]\, 
        REG_3 => \REG[444]\, REG_4 => \REG[445]\, REG_5 => 
        \REG[446]\, TICK(2) => \TICK[2]\, nLBRDY_c => nLBRDY_c, 
        EVNT_TRG => \I10.EVNT_TRG\, HWRES_c_32_0 => HWRES_c_32_0, 
        RUN_c => RUN_c, HWRES_c_34 => HWRES_c_34, CLK_c_c => 
        CLK_c_c, HWRES_c_33 => HWRES_c_33, N_18 => N_18, N_20 => 
        N_20, N_22 => N_22, N_24 => N_24, N_26 => N_26, N_28 => 
        N_28);
    
    \LBSP_pad[29]\ : IOB33PH
      port map(PAD => LBSP(29), A => \REG[374]\, EN => 
        \REG_i_0[294]\, Y => \LBSP_in[29]\);
    
    \LBSP_pad[4]\ : OB33PH
      port map(PAD => LBSP(4), A => L0_c_c);
    
    \AE_PDL_pad[8]\ : OB33PH
      port map(PAD => AE_PDL(8), A => \AE_PDL_c[8]\);
    
    L1R_pad : IB33
      port map(PAD => L1R, Y => L1R_c_c);
    
    ALICLK_pad : GL33
      port map(PAD => ALICLK, GL => ALICLK_c);
    
    \VAD_pad[21]\ : OTB33PH
      port map(PAD => VAD(21), A => \I2.VADm[21]\, EN => 
        NOEAD_c_1);
    
    \SYNC_pad[11]\ : OB33PH
      port map(PAD => SYNC(11), A => \SYNC_c[11]\);
    
    \VAD_pad[24]\ : OTB33PH
      port map(PAD => VAD(24), A => \I2.VADm[24]\, EN => 
        NOEAD_c_1);
    
    \VDB_pad[6]\ : IOB33PH
      port map(PAD => VDB(6), A => \I2.VDBm[6]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[6]\);
    
    \VAD_pad[23]\ : OTB33PH
      port map(PAD => VAD(23), A => \I2.VADm[23]\, EN => 
        NOEAD_c_1);
    
    \P_PDL_pad[4]\ : OB33PH
      port map(PAD => P_PDL(4), A => \P_PDL_c[4]\);
    
    \AE_PDL_pad[24]\ : OB33PH
      port map(PAD => AE_PDL(24), A => \AE_PDL_c[24]\);
    
    \VDB_pad_0[4]\ : BFR
      port map(A => \VDB_in[4]\, Y => \VDB_in_0[4]\);
    
    NOE64R_pad : OB33PH
      port map(PAD => NOE64R, A => NOEAD_c_i_0);
    
    \AE_PDL_pad[25]\ : OB33PH
      port map(PAD => AE_PDL(25), A => \AE_PDL_c[25]\);
    
    \VAD_pad[7]\ : IOB33PH
      port map(PAD => VAD(7), A => \I2.VADm[7]\, EN => NOEAD_c, Y
         => \VAD_in[7]\);
    
    L2R_pad : IB33
      port map(PAD => L2R, Y => L2R_c_c);
    
    \SYNC_pad[8]\ : OB33PH
      port map(PAD => SYNC(8), A => \SYNC_c[8]\);
    
    \VDB_pad[23]\ : IOB33PH
      port map(PAD => VDB(23), A => \I2.VDBm[23]\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[23]\);
    
    \SP_PDL_pad[43]\ : IOB33PH
      port map(PAD => SP_PDL(43), A => \I3.P0[43]\, EN => 
        MD_PDL_c, Y => \SP_PDL_in[43]\);
    
    \LED_pad[1]\ : OB33PH
      port map(PAD => LED(1), A => N_20);
    
    \LB_pad[3]\ : IOB33PH
      port map(PAD => LB(3), A => \I2.LB_i[3]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[3]\);
    
    \GA_pad[2]\ : IB33
      port map(PAD => GA(2), Y => \GA_c[2]\);
    
    \AE_PDL_pad[11]\ : OB33PH
      port map(PAD => AE_PDL(11), A => \AE_PDL_c[11]\);
    
    \P_PDL_pad[2]\ : OB33PH
      port map(PAD => P_PDL(2), A => \P_PDL_c[2]\);
    
    \VDB_pad[24]\ : IOB33PH
      port map(PAD => VDB(24), A => \I2.VDBm[24]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[24]\);
    
    \AE_PDL_pad[28]\ : OB33PH
      port map(PAD => AE_PDL(28), A => \AE_PDL_c[28]\);
    
    \AE_PDL_pad[22]\ : OB33PH
      port map(PAD => AE_PDL(22), A => \AE_PDL_c[22]\);
    
    ADLTC_pad : OB33PH
      port map(PAD => ADLTC, A => \GND\);
    
    \VAD_pad[11]\ : IOB33PH
      port map(PAD => VAD(11), A => \I2.VADm[11]\, EN => 
        NOEAD_c_0, Y => \VAD_in[11]\);
    
    \VDB_pad[22]\ : IOB33PH
      port map(PAD => VDB(22), A => \I2.VDBm[22]\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[22]\);
    
    \VAD_pad[27]\ : OTB33PH
      port map(PAD => VAD(27), A => \I2.VADm[27]\, EN => 
        NOEAD_c_1);
    
    \VAD_pad[14]\ : IOB33PH
      port map(PAD => VAD(14), A => \I2.VADm[14]\, EN => 
        NOEAD_c_0_0, Y => \VAD_in[14]\);
    
    \SP_PDL_pad[0]\ : IOB33PH
      port map(PAD => SP_PDL(0), A => \I3.P0[0]\, EN => 
        MD_PDL_c_0, Y => \SP_PDL_in[0]\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \SP_PDL_pad[4]\ : IOB33PH
      port map(PAD => SP_PDL(4), A => \I3.P0[4]\, EN => MD_PDL_c, 
        Y => \SP_PDL_in[4]\);
    
    \VAD_pad[13]\ : IOB33PH
      port map(PAD => VAD(13), A => \I2.VADm[13]\, EN => 
        NOEAD_c_0_0, Y => \VAD_in[13]\);
    
    NPWON_pad_1 : BFR
      port map(A => NPWON_c, Y => NPWON_c_1);
    
    \SP_PDL_pad[30]\ : IOB33PH
      port map(PAD => SP_PDL(30), A => \I3.P0[30]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[30]\);
    
    \LBSP_pad[31]\ : IOB33PH
      port map(PAD => LBSP(31), A => \REG[376]\, EN => 
        \REG_i_0[296]\, Y => \LBSP_in[31]\);
    
    \VDB_pad[16]\ : IOB33PH
      port map(PAD => VDB(16), A => \I2.VDBm[16]\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[16]\);
    
    \SP_PDL_pad[32]\ : IOB33PH
      port map(PAD => SP_PDL(32), A => \I3.P0[32]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[32]\);
    
    \VAD_pad[31]\ : IOB33PH
      port map(PAD => VAD(31), A => \I2.VADm[31]\, EN => NOEAD_c, 
        Y => \VAD_in[31]\);
    
    I8 : DAC_INTERF
      port map(TICK_0(2) => \TICK_0[2]\, SYNC_c(15) => 
        \SYNC_c[15]\, SYNC_c(14) => \SYNC_c[14]\, SYNC_c(13) => 
        \SYNC_c[13]\, SYNC_c(12) => \SYNC_c[12]\, SYNC_c(11) => 
        \SYNC_c[11]\, SYNC_c(10) => \SYNC_c[10]\, SYNC_c(9) => 
        \SYNC_c[9]\, SYNC_c(8) => \SYNC_c[8]\, SYNC_c(7) => 
        \SYNC_c[7]\, SYNC_c(6) => \SYNC_c[6]\, SYNC_c(5) => 
        \SYNC_c[5]\, SYNC_c(4) => \SYNC_c[4]\, SYNC_c(3) => 
        \SYNC_c[3]\, SYNC_c(2) => \SYNC_c[2]\, SYNC_c(1) => 
        \SYNC_c[1]\, SYNC_c(0) => \SYNC_c[0]\, DACCFG_DT(15) => 
        \DACCFG_DT[15]\, DACCFG_DT(14) => \DACCFG_DT[14]\, 
        DACCFG_DT(13) => \DACCFG_DT[13]\, DACCFG_DT(12) => 
        \DACCFG_DT[12]\, DACCFG_DT(11) => \DACCFG_DT[11]\, 
        DACCFG_DT(10) => \DACCFG_DT[10]\, DACCFG_DT(9) => 
        \DACCFG_DT[9]\, DACCFG_DT(8) => \DACCFG_DT[8]\, 
        DACCFG_DT(7) => \DACCFG_DT[7]\, DACCFG_DT(6) => 
        \DACCFG_DT[6]\, DACCFG_DT(5) => \DACCFG_DT[5]\, 
        DACCFG_DT(4) => \DACCFG_DT[4]\, DACCFG_DT(3) => 
        \DACCFG_DT[3]\, DACCFG_DT(2) => \DACCFG_DT[2]\, 
        DACCFG_DT(1) => \DACCFG_DT[1]\, DACCFG_DT(0) => 
        \DACCFG_DT[0]\, REG(264) => \REG[264]\, REG(263) => 
        \REG[263]\, REG(262) => \REG[262]\, REG(261) => 
        \REG[261]\, REG(260) => \REG[260]\, REG(259) => 
        \REG[259]\, REG(258) => \REG[258]\, REG(257) => 
        \REG[257]\, REG(256) => \REG[256]\, REG(255) => 
        \REG[255]\, REG(254) => \REG[254]\, REG(253) => 
        \REG[253]\, REG(252) => \REG[252]\, REG(251) => 
        \REG[251]\, REG(250) => \REG[250]\, REG(249) => 
        \REG[249]\, REG(248) => \REG[248]\, REG(247) => 
        \REG[247]\, REG(246) => \REG[246]\, REG(245) => 
        \REG[245]\, REG(244) => \REG[244]\, REG(243) => 
        \REG[243]\, REG(242) => \REG[242]\, REG(241) => 
        \REG[241]\, REG(240) => \REG[240]\, REG(239) => 
        \REG[239]\, REG(238) => \REG[238]\, REG(237) => 
        \REG[237]\, REG(236) => \REG[236]\, REG(235) => 
        \REG[235]\, REG(234) => \REG[234]\, REG(233) => 
        \REG[233]\, PULSE(9) => \PULSE[9]\, DACCFG_RAD(3) => 
        \DACCFG_RAD[3]\, DACCFG_RAD(2) => \DACCFG_RAD[2]\, 
        DACCFG_RAD(1) => \DACCFG_RAD[1]\, DACCFG_RAD(0) => 
        \DACCFG_RAD[0]\, HWRES_c_36 => HWRES_c_36, HWRES_c_34 => 
        HWRES_c_34, HWRES_c_35 => HWRES_c_35, RUN_c_0 => RUN_c_0, 
        DACCFG_nRD => DACCFG_nRD, SCLK_DAC_c => SCLK_DAC_c, 
        SDIN_DAC_c => SDIN_DAC_c, HWRES_c_0 => HWRES_c_0, 
        HWRES_c_3 => HWRES_c_3, HWRES_c_0_6_0 => HWRES_c_0_6_0, 
        HWRES_c_2 => HWRES_c_2, HWRES_c_1 => HWRES_c_1, 
        HWRES_c_36_0 => HWRES_c_36_0, CLK_c_c => CLK_c_c, HWRES_c
         => HWRES_c);
    
    \SP_PDL_pad[21]\ : IOB33PH
      port map(PAD => SP_PDL(21), A => \I3.P0[21]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[21]\);
    
    \LBSP_pad[12]\ : OB33PH
      port map(PAD => LBSP(12), A => SPULSE1_c_c);
    
    PSM_RES_pad : OB33PH
      port map(PAD => PSM_RES, A => \GND\);
    
    \SP_PDL_pad[10]\ : IOB33PH
      port map(PAD => SP_PDL(10), A => \I3.P0[10]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[10]\);
    
    \AE_PDL_pad[36]\ : OB33PH
      port map(PAD => AE_PDL(36), A => \AE_PDL_c[36]\);
    
    \AE_PDL_pad[33]\ : OB33PH
      port map(PAD => AE_PDL(33), A => \AE_PDL_c[33]\);
    
    \LB_pad[8]\ : IOB33PH
      port map(PAD => LB(8), A => \I2.LB_i[8]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[8]\);
    
    \SYNC_pad[9]\ : OB33PH
      port map(PAD => SYNC(9), A => \SYNC_c[9]\);
    
    \SP_PDL_pad[12]\ : IOB33PH
      port map(PAD => SP_PDL(12), A => \I3.P0[12]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[12]\);
    
    \AE_PDL_pad[14]\ : OB33PH
      port map(PAD => AE_PDL(14), A => \AE_PDL_c[14]\);
    
    \SYNC_pad[14]\ : OB33PH
      port map(PAD => SYNC(14), A => \SYNC_c[14]\);
    
    \SP_PDL_pad[45]\ : IOB33PH
      port map(PAD => SP_PDL(45), A => \I3.P0[45]\, EN => 
        MD_PDL_c, Y => \SP_PDL_in[45]\);
    
    \AE_PDL_pad[15]\ : OB33PH
      port map(PAD => AE_PDL(15), A => \AE_PDL_c[15]\);
    
    \VAD_pad[17]\ : OTB33PH
      port map(PAD => VAD(17), A => \I2.VADm[17]\, EN => 
        NOEAD_c_1);
    
    \SP_PDL_pad[9]\ : IOB33PH
      port map(PAD => SP_PDL(9), A => \I3.P0[9]\, EN => MD_PDL_c, 
        Y => \SP_PDL_in[9]\);
    
    \SYNC_pad[12]\ : OB33PH
      port map(PAD => SYNC(12), A => \SYNC_c[12]\);
    
    \LBSP_pad[6]\ : OB33PH
      port map(PAD => LBSP(6), A => L1R_c_c);
    
    INTR1_pad : OB33PH
      port map(PAD => INTR1, A => \VCC\);
    
    \VDB_pad[15]\ : IOB33PH
      port map(PAD => VDB(15), A => \I2.VDBm[15]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[15]\);
    
    \TST_pad[10]\ : OTB33PH
      port map(PAD => TST(10), A => \GND\, EN => \GND\);
    
    \VDB_pad[3]\ : IOB33PH
      port map(PAD => VDB(3), A => \I2.VDBm[3]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[3]\);
    
    \P_PDL_pad[6]\ : OB33PH
      port map(PAD => P_PDL(6), A => \P_PDL_c[6]\);
    
    \AE_PDL_pad[18]\ : OB33PH
      port map(PAD => AE_PDL(18), A => \AE_PDL_c[18]\);
    
    \AE_PDL_pad[12]\ : OB33PH
      port map(PAD => AE_PDL(12), A => \AE_PDL_c[12]\);
    
    \VAD_pad[25]\ : OTB33PH
      port map(PAD => VAD(25), A => \I2.VADm[25]\, EN => 
        NOEAD_c_1);
    
    \SP_PDL_pad[23]\ : IOB33PH
      port map(PAD => SP_PDL(23), A => \I3.P0[23]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[23]\);
    
    \LBSP_pad[3]\ : OB33PH
      port map(PAD => LBSP(3), A => EV_RES_c);
    
    \LBSP_pad[10]\ : OB33PH
      port map(PAD => LBSP(10), A => LOS_c_c);
    
    SPULSE1_pad : IB33
      port map(PAD => SPULSE1, Y => SPULSE1_c_c);
    
    \AE_PDL_pad[41]\ : OB33PH
      port map(PAD => AE_PDL(41), A => \AE_PDL_c[41]\);
    
    \LBSP_pad[1]\ : IOB33PH
      port map(PAD => LBSP(1), A => \REG[346]\, EN => 
        \REG_i_0[266]\, Y => \LBSP_in[1]\);
    
    \LBSP_pad[14]\ : OB33PH
      port map(PAD => LBSP(14), A => \REG_c[0]\);
    
    NSELCLK_pad : OB33PH
      port map(PAD => NSELCLK, A => NSELCLK_c);
    
    \SYNC_pad[2]\ : OB33PH
      port map(PAD => SYNC(2), A => \SYNC_c[2]\);
    
    RSELC0_pad : OTB33PH
      port map(PAD => RSELC0, A => \REG[380]\, EN => 
        \REG_i_0[396]\);
    
    \VDB_pad[19]\ : IOB33PH
      port map(PAD => VDB(19), A => \I2.VDBm[19]\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[19]\);
    
    \LED_pad[5]\ : OB33PH
      port map(PAD => LED(5), A => N_28);
    
    \TST_pad[3]\ : OB33PH
      port map(PAD => TST(3), A => \TST_c_c[3]\);
    
    \DIR_CTTM_pad[3]\ : OB33PH
      port map(PAD => DIR_CTTM(3), A => \VCC\);
    
    \LBSP_pad[28]\ : IOB33PH
      port map(PAD => LBSP(28), A => \REG[373]\, EN => 
        \REG_i_0[293]\, Y => \LBSP_in[28]\);
    
    I_16 : INV
      port map(A => EVREAD, Y => \I_16\);
    
    \TST_pad[0]\ : OB33PH
      port map(PAD => TST(0), A => \TST_c[0]\);
    
    NLBRD_pad : OB33PH
      port map(PAD => NLBRD, A => NLBRD_c);
    
    \VAD_pad[15]\ : IOB33PH
      port map(PAD => VAD(15), A => \I2.VADm[15]\, EN => 
        NOEAD_c_0_0, Y => \VAD_in[15]\);
    
    \SP_PDL_pad[28]\ : IOB33PH
      port map(PAD => SP_PDL(28), A => \I3.P0[28]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[28]\);
    
    \AE_PDL_pad[37]\ : OB33PH
      port map(PAD => AE_PDL(37), A => \AE_PDL_c[37]\);
    
    \TST_pad[5]\ : OB33PH
      port map(PAD => TST(5), A => \TST_c[5]\);
    
    SCL1_pad : OB33PH
      port map(PAD => SCL1, A => SCLB_i_a3);
    
    \VDB_pad[7]\ : IOB33PH
      port map(PAD => VDB(7), A => \I2.VDBm[7]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[7]\);
    
    \SP_PDL_pad[37]\ : IOB33PH
      port map(PAD => SP_PDL(37), A => \I3.P0[37]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[37]\);
    
    \SP_PDL_pad[25]\ : IOB33PH
      port map(PAD => SP_PDL(25), A => \I3.P0[25]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[25]\);
    
    \LBSP_pad[25]\ : IOB33PH
      port map(PAD => LBSP(25), A => \REG[370]\, EN => 
        \REG_i_0[290]\, Y => \LBSP_in[25]\);
    
    \VAD_pad[29]\ : IOB33PH
      port map(PAD => VAD(29), A => \I2.VADm[29]\, EN => NOEAD_c, 
        Y => \VAD_in[29]\);
    
    \VDB_pad_0[6]\ : BFR
      port map(A => \VDB_in[6]\, Y => \VDB_in_0[6]\);
    
    \LED_pad[4]\ : OB33PH
      port map(PAD => LED(4), A => N_26);
    
    F_SCK_pad : OTB33PH
      port map(PAD => F_SCK, A => \I5.ISCK\, EN => un1_drive_spi);
    
    \AE_PDL_pad[44]\ : OB33PH
      port map(PAD => AE_PDL(44), A => \AE_PDL_c[44]\);
    
    \AE_PDL_pad[1]\ : OB33PH
      port map(PAD => AE_PDL(1), A => \AE_PDL_c[1]\);
    
    \VDB_pad_0[3]\ : BFR
      port map(A => \VDB_in[3]\, Y => \VDB_in_0[3]\);
    
    \LED_pad[0]\ : OB33PH
      port map(PAD => LED(0), A => N_18);
    
    \AE_PDL_pad[45]\ : OB33PH
      port map(PAD => AE_PDL(45), A => \AE_PDL_c[45]\);
    
    \VAD_pad[28]\ : IOB33PH
      port map(PAD => VAD(28), A => \I2.VADm[28]\, EN => NOEAD_c, 
        Y => \VAD_in[28]\);
    
    NPWON_pad_2 : BFR
      port map(A => NPWON_c, Y => NPWON_c_2);
    
    \DIR_CTTM_pad[5]\ : OB33PH
      port map(PAD => DIR_CTTM(5), A => \VCC\);
    
    \SP_PDL_pad[17]\ : IOB33PH
      port map(PAD => SP_PDL(17), A => \I3.P0[17]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[17]\);
    
    \AE_PDL_pad[26]\ : OB33PH
      port map(PAD => AE_PDL(26), A => \AE_PDL_c[26]\);
    
    \AE_PDL_pad[23]\ : OB33PH
      port map(PAD => AE_PDL(23), A => \AE_PDL_c[23]\);
    
    IACKB_pad : IB33
      port map(PAD => IACKB, Y => IACKB_c);
    
    \TST_pad[8]\ : OTB33PH
      port map(PAD => TST(8), A => \GND\, EN => \GND\);
    
    LOS_pad : IB33
      port map(PAD => LOS, Y => LOS_c_c);
    
    \AE_PDL_pad[42]\ : OB33PH
      port map(PAD => AE_PDL(42), A => \AE_PDL_c[42]\);
    
    \VDB_pad[30]\ : IOB33PH
      port map(PAD => VDB(30), A => \I2.VDBm[30]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[30]\);
    
    LTM_DRDY_pad : OB33PH
      port map(PAD => LTM_DRDY, A => EVRDY_c);
    
    \LB_pad[9]\ : IOB33PH
      port map(PAD => LB(9), A => \I2.LB_i[9]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[9]\);
    
    NPWON_pad_3 : BFR
      port map(A => NPWON_c, Y => NPWON_c_3);
    
    \VAD_pad[5]\ : IOB33PH
      port map(PAD => VAD(5), A => \I2.VADm[5]\, EN => NOEAD_c, Y
         => \VAD_in[5]\);
    
    \VAD_pad[19]\ : OTB33PH
      port map(PAD => VAD(19), A => \I2.VADm[19]\, EN => 
        NOEAD_c_1);
    
    \LBSP_pad[8]\ : OB33PH
      port map(PAD => LBSP(8), A => L2R_c_c);
    
    \SP_PDL_pad[39]\ : IOB33PH
      port map(PAD => SP_PDL(39), A => \I3.P0[39]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[39]\);
    
    \VAD_pad[4]\ : IOB33PH
      port map(PAD => VAD(4), A => \I2.VADm[4]\, EN => NOEAD_c, Y
         => \VAD_in[4]\);
    
    \VAD_pad[2]\ : IOB33PH
      port map(PAD => VAD(2), A => \I2.VADm[2]\, EN => NOEAD_c, Y
         => \VAD_in[2]\);
    
    \VAD_pad[18]\ : OTB33PH
      port map(PAD => VAD(18), A => \I2.VADm[18]\, EN => 
        NOEAD_c_1);
    
    \LBSP_pad[30]\ : IOB33PH
      port map(PAD => LBSP(30), A => \REG[375]\, EN => 
        \REG_i_0[295]\, Y => \LBSP_in[30]\);
    
    PSM_SP3_pad : IB33
      port map(PAD => PSM_SP3, Y => \REG_c[21]\);
    
    nLBAS_pad : OB33PH
      port map(PAD => nLBAS, A => nLBAS_c);
    
    RSELC1_pad : OTB33PH
      port map(PAD => RSELC1, A => \REG[379]\, EN => 
        \REG_i_0[395]\);
    
    \LB_pad[7]\ : IOB33PH
      port map(PAD => LB(7), A => \I2.LB_i[7]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[7]\);
    
    \VAD_pad[9]\ : IOB33PH
      port map(PAD => VAD(9), A => \I2.VADm[9]\, EN => NOEAD_c, Y
         => \VAD_in[9]\);
    
    \SP_PDL_pad[8]\ : IOB33PH
      port map(PAD => SP_PDL(8), A => \I3.P0[8]\, EN => MD_PDL_c, 
        Y => \SP_PDL_in[8]\);
    
    SCLK_DAC_pad : OB33PH
      port map(PAD => SCLK_DAC, A => SCLK_DAC_c);
    
    NLBRES_pad : OB33PH
      port map(PAD => NLBRES, A => HWRES_c_i_0);
    
    MYBERR_pad : OB33PH
      port map(PAD => MYBERR, A => MYBERR_c);
    
    \VDB_pad_0[9]\ : BFR
      port map(A => \VDB_in[9]\, Y => \VDB_in_0[9]\);
    
    \VAD_pad[8]\ : IOB33PH
      port map(PAD => VAD(8), A => \I2.VADm[8]\, EN => NOEAD_c, Y
         => \VAD_in[8]\);
    
    \TST_pad[15]\ : OB33PH
      port map(PAD => TST(15), A => \TST_c[15]\);
    
    \SP_PDL_pad[19]\ : IOB33PH
      port map(PAD => SP_PDL(19), A => \I3.P0[19]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[19]\);
    
    NOE16W_pad : OB33PH
      port map(PAD => NOE16W, A => NOE16W_c);
    
    I_8 : INV
      port map(A => \I10.un2_evread[14]\, Y => \I_8\);
    
    \TST_pad[13]\ : OB33PH
      port map(PAD => TST(13), A => \TST_c[13]\);
    
    \LB_pad[6]\ : IOB33PH
      port map(PAD => LB(6), A => \I2.LB_i[6]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[6]\);
    
    \VDB_pad_0[10]\ : BFR
      port map(A => \VDB_in[10]\, Y => \VDB_in_0[10]\);
    
    \LBSP_pad[19]\ : IOB33PH
      port map(PAD => LBSP(19), A => \REG[364]\, EN => 
        \REG_i_0[284]\, Y => \LBSP_in[19]\);
    
    DS1B_pad : IB33
      port map(PAD => DS1B, Y => DS1B_c);
    
    \AE_PDL_pad[16]\ : OB33PH
      port map(PAD => AE_PDL(16), A => \AE_PDL_c[16]\);
    
    \AE_PDL_pad[13]\ : OB33PH
      port map(PAD => AE_PDL(13), A => \AE_PDL_c[13]\);
    
    \VDB_pad[31]\ : IOB33PH
      port map(PAD => VDB(31), A => \I2.VDBm[31]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[31]\);
    
    \VDB_pad[13]\ : IOB33PH
      port map(PAD => VDB(13), A => \I2.VDBm[13]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[13]\);
    
    NOE32W_pad : OB33PH
      port map(PAD => NOE32W, A => NOE32W_c);
    
    \AE_PDL_pad[4]\ : OB33PH
      port map(PAD => AE_PDL(4), A => \AE_PDL_c[4]\);
    
    \SP_PDL_pad[44]\ : IOB33PH
      port map(PAD => SP_PDL(44), A => \I3.P0[44]\, EN => 
        MD_PDL_c, Y => \SP_PDL_in[44]\);
    
    NPWON_pad_0 : BFR
      port map(A => NPWON_c, Y => NPWON_c_0);
    
    \DIR_CTTM_pad[6]\ : OB33PH
      port map(PAD => DIR_CTTM(6), A => \VCC\);
    
    \TST_pad_i[7]\ : INV
      port map(A => \I2.un7_noe32ri_0\, Y => \I2.un7_noe32ri_i_0\);
    
    \SP_PDL_pad[3]\ : IOB33PH
      port map(PAD => SP_PDL(3), A => \I3.P0[3]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[3]\);
    
    NOE32R_pad : OB33PH
      port map(PAD => NOE32R, A => \I2.un7_noe32ri_i_0\);
    
    \AE_PDL_pad[27]\ : OB33PH
      port map(PAD => AE_PDL(27), A => \AE_PDL_c[27]\);
    
    \VDB_pad[14]\ : IOB33PH
      port map(PAD => VDB(14), A => \I2.VDBm[14]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[14]\);
    
    SDIN_DAC_pad : OB33PH
      port map(PAD => SDIN_DAC, A => SDIN_DAC_c);
    
    \LB_pad_i_0[31]\ : INV
      port map(A => \I2.LB_nOE\, Y => \I2.LB_nOE_i_0_0\);
    
    \SP_PDL_pad[46]\ : IOB33PH
      port map(PAD => SP_PDL(46), A => \I3.P0[46]\, EN => 
        MD_PDL_c, Y => \SP_PDL_in[46]\);
    
    NLBWAIT_pad : OB33PH
      port map(PAD => NLBWAIT, A => \VCC\);
    
    LTM_BUSY_pad : OB33PH
      port map(PAD => LTM_BUSY, A => \REG[17]\);
    
    \TST_pad[6]\ : OB33PH
      port map(PAD => TST(6), A => \I2.un5_noe16ri_i_0\);
    
    \VDB_pad[27]\ : IOB33PH
      port map(PAD => VDB(27), A => \I2.VDBm[27]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[27]\);
    
    \VDB_pad[12]\ : IOB33PH
      port map(PAD => VDB(12), A => \I2.VDBm[12]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[12]\);
    
    ASB_pad : GL33
      port map(PAD => ASB, GL => ASB_c);
    
    \VAD_pad[20]\ : OTB33PH
      port map(PAD => VAD(20), A => \I2.VADm[20]\, EN => 
        NOEAD_c_1);
    
    SDA1_pad : IOB33PH
      port map(PAD => SDA1, A => \I1.SDAout_del2\, EN => 
        un1_sdab_i, Y => SDA1_in);
    
    \VAD_pad[1]\ : IOB33PH
      port map(PAD => VAD(1), A => \I2.VADm[1]\, EN => NOEAD_c_1, 
        Y => \VAD_in[1]\);
    
    \SYNC_pad[1]\ : OB33PH
      port map(PAD => SYNC(1), A => \SYNC_c[1]\);
    
    FCS_pad : OB33PH
      port map(PAD => FCS, A => FCS_c);
    
    RSELA0_pad : OTB33PH
      port map(PAD => RSELA0, A => \REG[384]\, EN => 
        \REG_i_0[400]\);
    
    \LB_pad[5]\ : IOB33PH
      port map(PAD => LB(5), A => \I2.LB_i[5]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[5]\);
    
    \LB_pad[12]\ : IOB33PH
      port map(PAD => LB(12), A => \I2.LB_i[12]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[12]\);
    
    \AE_PDL_pad[3]\ : OB33PH
      port map(PAD => AE_PDL(3), A => \AE_PDL_c[3]\);
    
    \DIR_CTTM_pad[7]\ : OB33PH
      port map(PAD => DIR_CTTM(7), A => \VCC\);
    
    \VDB_pad[28]\ : IOB33PH
      port map(PAD => VDB(28), A => \I2.VDBm[28]\, EN => 
        un7_noe32ri_0_0, Y => \VDB_in[28]\);
    
    PSM_SP4_pad : IB33
      port map(PAD => PSM_SP4, Y => \REG_c[22]\);
    
    \AMB_pad[3]\ : IB33
      port map(PAD => AMB(3), Y => \AMB_c[3]\);
    
    \SP_PDL_pad[31]\ : IOB33PH
      port map(PAD => SP_PDL(31), A => \I3.P0[31]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[31]\);
    
    \SYNC_pad[15]\ : OB33PH
      port map(PAD => SYNC(15), A => \SYNC_c[15]\);
    
    L1A_pad : IB33
      port map(PAD => L1A, Y => L1A_c_c);
    
    \VDB_pad[0]\ : IOB33PH
      port map(PAD => VDB(0), A => \I2.VDBm[0]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[0]\);
    
    F_SO_pad : IB33
      port map(PAD => F_SO, Y => F_SO_c);
    
    \SP_PDL_pad[1]\ : IOB33PH
      port map(PAD => SP_PDL(1), A => \I3.P0[1]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[1]\);
    
    \LB_pad[22]\ : IOB33PH
      port map(PAD => LB(22), A => \I2.LB_i[22]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[22]\);
    
    L2A_pad : IB33
      port map(PAD => L2A, Y => L2A_c_c);
    
    \VAD_pad[10]\ : IOB33PH
      port map(PAD => VAD(10), A => \I2.VADm[10]\, EN => 
        NOEAD_c_0, Y => \VAD_in[10]\);
    
    \LB_pad_i[31]\ : INV
      port map(A => \I2.LB_nOE\, Y => \I2.LB_nOE_i_0\);
    
    \DIR_CTTM_pad[1]\ : OB33PH
      port map(PAD => DIR_CTTM(1), A => \VCC\);
    
    \SP_PDL_pad[11]\ : IOB33PH
      port map(PAD => SP_PDL(11), A => \I3.P0[11]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[11]\);
    
    \LB_pad_i_1[31]\ : INV
      port map(A => \I2.LB_nOE\, Y => \I2.LB_nOE_i_0_1\);
    
    \LBSP_pad[27]\ : IOB33PH
      port map(PAD => LBSP(27), A => \REG[372]\, EN => 
        \REG_i_0[292]\, Y => \LBSP_in[27]\);
    
    \VDB_pad_0[13]\ : BFR
      port map(A => \VDB_in[13]\, Y => \VDB_in_0[13]\);
    
    \AE_PDL_pad[17]\ : OB33PH
      port map(PAD => AE_PDL(17), A => \AE_PDL_c[17]\);
    
    \SYNC_pad[10]\ : OB33PH
      port map(PAD => SYNC(10), A => \SYNC_c[10]\);
    
    \SYNC_pad[0]\ : OB33PH
      port map(PAD => SYNC(0), A => \SYNC_c[0]\);
    
    \VAD_pad[6]\ : IOB33PH
      port map(PAD => VAD(6), A => \I2.VADm[6]\, EN => NOEAD_c, Y
         => \VAD_in[6]\);
    
    \VDB_pad[20]\ : IOB33PH
      port map(PAD => VDB(20), A => \I2.VDBm[20]\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[20]\);
    
    \LBSP_pad[21]\ : IOB33PH
      port map(PAD => LBSP(21), A => \REG[366]\, EN => 
        \REG_i_0[286]\, Y => \LBSP_in[21]\);
    
    \TST_pad[7]\ : OB33PH
      port map(PAD => TST(7), A => \I2.un7_noe32ri_i_0\);
    
    SI_PDL_pad : OB33PH
      port map(PAD => SI_PDL, A => SI_PDL_c);
    
    SELCLK_pad : OB33PH
      port map(PAD => SELCLK, A => NSELCLK_c_i_0);
    
    I14 : DACCFG
      port map(DACCFG_WDT(13) => \DACCFG_WDT[13]\, DACCFG_WDT(12)
         => \DACCFG_WDT[12]\, DACCFG_WDT(11) => \DACCFG_WDT[11]\, 
        DACCFG_WDT(10) => \DACCFG_WDT[10]\, DACCFG_WDT(9) => 
        \DACCFG_WDT[9]\, DACCFG_WDT(8) => \DACCFG_WDT[8]\, 
        DACCFG_WDT(7) => \DACCFG_WDT[7]\, DACCFG_WDT(6) => 
        \DACCFG_WDT[6]\, DACCFG_WDT(5) => \DACCFG_WDT[5]\, 
        DACCFG_WDT(4) => \DACCFG_WDT[4]\, DACCFG_RAD(3) => 
        \DACCFG_RAD[3]\, DACCFG_RAD(2) => \DACCFG_RAD[2]\, 
        DACCFG_RAD(1) => \DACCFG_RAD[1]\, DACCFG_RAD(0) => 
        \DACCFG_RAD[0]\, DACCFG_DT(15) => \DACCFG_DT[15]\, 
        DACCFG_DT(14) => \DACCFG_DT[14]\, DACCFG_DT(13) => 
        \DACCFG_DT[13]\, DACCFG_DT(12) => \DACCFG_DT[12]\, 
        DACCFG_DT(11) => \DACCFG_DT[11]\, DACCFG_DT(10) => 
        \DACCFG_DT[10]\, DACCFG_DT(9) => \DACCFG_DT[9]\, 
        DACCFG_DT(8) => \DACCFG_DT[8]\, DACCFG_DT(7) => 
        \DACCFG_DT[7]\, DACCFG_DT(6) => \DACCFG_DT[6]\, 
        DACCFG_DT(5) => \DACCFG_DT[5]\, DACCFG_DT(4) => 
        \DACCFG_DT[4]\, DACCFG_DT(3) => \DACCFG_DT[3]\, 
        DACCFG_DT(2) => \DACCFG_DT[2]\, DACCFG_DT(1) => 
        \DACCFG_DT[1]\, DACCFG_DT(0) => \DACCFG_DT[0]\, 
        CROMWAD(4) => \CROMWAD[4]\, CROMWAD(3) => \CROMWAD[3]\, 
        CROMWAD(2) => \CROMWAD[2]\, CROMWAD(1) => \CROMWAD[1]\, 
        DACCFG_nRD => DACCFG_nRD, DACCFG_nWR => DACCFG_nWR, 
        CLK_c_c => CLK_c_c);
    
    \VAD_pad[30]\ : IOB33PH
      port map(PAD => VAD(30), A => \I2.VADm[30]\, EN => NOEAD_c, 
        Y => \VAD_in[30]\);
    
    \SP_PDL_pad[24]\ : IOB33PH
      port map(PAD => SP_PDL(24), A => \I3.P0[24]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[24]\);
    
    \LED_pad[3]\ : OB33PH
      port map(PAD => LED(3), A => N_24);
    
    \AE_PDL_pad[46]\ : OB33PH
      port map(PAD => AE_PDL(46), A => \AE_PDL_c[46]\);
    
    \AE_PDL_pad[43]\ : OB33PH
      port map(PAD => AE_PDL(43), A => \AE_PDL_c[43]\);
    
    \AE_PDL_pad[30]\ : OB33PH
      port map(PAD => AE_PDL(30), A => \AE_PDL_c[30]\);
    
    \VAD_pad[26]\ : OTB33PH
      port map(PAD => VAD(26), A => \I2.VADm[26]\, EN => 
        NOEAD_c_1);
    
    \AMB_pad[4]\ : IB33
      port map(PAD => AMB(4), Y => \AMB_c[4]\);
    
    \SP_PDL_pad[33]\ : IOB33PH
      port map(PAD => SP_PDL(33), A => \I3.P0[33]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[33]\);
    
    \SP_PDL_pad[26]\ : IOB33PH
      port map(PAD => SP_PDL(26), A => \I3.P0[26]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[26]\);
    
    \DIR_CTTM_pad[4]\ : OB33PH
      port map(PAD => DIR_CTTM(4), A => \VCC\);
    
    \SP_PDL_pad[2]\ : IOB33PH
      port map(PAD => SP_PDL(2), A => \I3.P0[2]\, EN => 
        MD_PDL_c_2, Y => \SP_PDL_in[2]\);
    
    \VDB_pad[5]\ : IOB33PH
      port map(PAD => VDB(5), A => \I2.VDBm[5]\, EN => 
        un5_noe16ri_0_0, Y => \VDB_in[5]\);
    
    \TST_pad[11]\ : OTB33PH
      port map(PAD => TST(11), A => \GND\, EN => \GND\);
    
    NDTKIN_pad : OB33PH
      port map(PAD => NDTKIN, A => NDTKIN_c);
    
    \VDB_pad[1]\ : IOB33PH
      port map(PAD => VDB(1), A => \I2.VDBm[1]\, EN => 
        \I2.un5_noe16ri_0\, Y => \VDB_in[1]\);
    
    \VAD_pad[22]\ : OTB33PH
      port map(PAD => VAD(22), A => \I2.VADm[22]\, EN => 
        NOEAD_c_1);
    
    \P_PDL_pad[3]\ : OB33PH
      port map(PAD => P_PDL(3), A => \P_PDL_c[3]\);
    
    \AE_PDL_pad[39]\ : OB33PH
      port map(PAD => AE_PDL(39), A => \AE_PDL_c[39]\);
    
    \LBSP_pad[9]\ : OB33PH
      port map(PAD => LBSP(9), A => RUN_c);
    
    \LBSP_pad[26]\ : IOB33PH
      port map(PAD => LBSP(26), A => \REG[371]\, EN => 
        \REG_i_0[291]\, Y => \LBSP_in[26]\);
    
    \VDB_pad_0[5]\ : BFR
      port map(A => \VDB_in[5]\, Y => \VDB_in_0[5]\);
    
    \DIR_CTTM_pad[0]\ : OB33PH
      port map(PAD => DIR_CTTM(0), A => \VCC\);
    
    \SP_PDL_pad[13]\ : IOB33PH
      port map(PAD => SP_PDL(13), A => \I3.P0[13]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[13]\);
    
    \LED_pad[2]\ : OB33PH
      port map(PAD => LED(2), A => N_22);
    
    \LB_pad[17]\ : IOB33PH
      port map(PAD => LB(17), A => \I2.LB_i[17]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[17]\);
    
    \LBSP_pad[23]\ : IOB33PH
      port map(PAD => LBSP(23), A => \REG[368]\, EN => 
        \REG_i_0[288]\, Y => \LBSP_in[23]\);
    
    NOEAD_pad : OB33PH
      port map(PAD => NOEAD, A => NOEAD_c_0);
    
    \SP_PDL_pad[40]\ : IOB33PH
      port map(PAD => SP_PDL(40), A => \I3.P0[40]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[40]\);
    
    \LB_pad[1]\ : IOB33PH
      port map(PAD => LB(1), A => \I2.LB_i[1]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[1]\);
    
    \SP_PDL_pad[42]\ : IOB33PH
      port map(PAD => SP_PDL(42), A => \I3.P0[42]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[42]\);
    
    RSELA1_pad : OTB33PH
      port map(PAD => RSELA1, A => \REG[383]\, EN => 
        \REG_i_0[399]\);
    
    \SP_PDL_pad[38]\ : IOB33PH
      port map(PAD => SP_PDL(38), A => \I3.P0[38]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[38]\);
    
    \VAD_pad[16]\ : OTB33PH
      port map(PAD => VAD(16), A => \I2.VADm[16]\, EN => 
        NOEAD_c_0_0);
    
    \P_PDL_pad[7]\ : OB33PH
      port map(PAD => P_PDL(7), A => \P_PDL_c[7]\);
    
    \AMB_pad[1]\ : IB33
      port map(PAD => AMB(1), Y => \AMB_c[1]\);
    
    \LBSP_pad[18]\ : IOB33PH
      port map(PAD => LBSP(18), A => \REG[363]\, EN => 
        \REG_i_0[283]\, Y => \LBSP_in[18]\);
    
    \VDB_pad[21]\ : IOB33PH
      port map(PAD => VDB(21), A => \I2.N_500\, EN => 
        \I2.un7_noe32ri_0\, Y => \VDB_in[21]\);
    
    \SYNC_pad[4]\ : OB33PH
      port map(PAD => SYNC(4), A => \SYNC_c[4]\);
    
    SPULSE2_pad : IB33
      port map(PAD => SPULSE2, Y => SPULSE2_c_c);
    
    \AE_PDL_pad[2]\ : OB33PH
      port map(PAD => AE_PDL(2), A => \AE_PDL_c[2]\);
    
    \VAD_pad[12]\ : IOB33PH
      port map(PAD => VAD(12), A => \I2.VADm[12]\, EN => 
        NOEAD_c_0_0, Y => \VAD_in[12]\);
    
    \SP_PDL_pad[35]\ : IOB33PH
      port map(PAD => SP_PDL(35), A => \I3.P0[35]\, EN => 
        MD_PDL_c_3, Y => \SP_PDL_in[35]\);
    
    \VDB_pad_0[1]\ : BFR
      port map(A => \VDB_in[1]\, Y => \VDB_in_0[1]\);
    
    \LB_pad[27]\ : IOB33PH
      port map(PAD => LB(27), A => \I2.LB_i[27]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[27]\);
    
    \LB_pad[13]\ : IOB33PH
      port map(PAD => LB(13), A => \I2.LB_i[13]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[13]\);
    
    \TST_pad[2]\ : OB33PH
      port map(PAD => TST(2), A => \TST_c[2]\);
    
    \SP_PDL_pad[18]\ : IOB33PH
      port map(PAD => SP_PDL(18), A => \I3.P0[18]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[18]\);
    
    RSELB0_pad : OTB33PH
      port map(PAD => RSELB0, A => \REG[382]\, EN => 
        \REG_i_0[398]\);
    
    \SP_PDL_pad[7]\ : IOB33PH
      port map(PAD => SP_PDL(7), A => \I3.P0[7]\, EN => MD_PDL_c, 
        Y => \SP_PDL_in[7]\);
    
    d_m6 : MUX2H
      port map(A => d_N_5, B => \REG[473]\, S => \I2.REGMAP[35]\, 
        Y => d_N_7);
    
    \P_PDL_pad[5]\ : OB33PH
      port map(PAD => P_PDL(5), A => \P_PDL_c[5]\);
    
    \AE_PDL_pad[47]\ : OB33PH
      port map(PAD => AE_PDL(47), A => \AE_PDL_c[47]\);
    
    \LBSP_pad[15]\ : IOB33PH
      port map(PAD => LBSP(15), A => \REG[360]\, EN => 
        \REG_i_0[280]\, Y => \LBSP_in[15]\);
    
    \AE_PDL_pad[6]\ : OB33PH
      port map(PAD => AE_PDL(6), A => \AE_PDL_c[6]\);
    
    \SYNC_pad[3]\ : OB33PH
      port map(PAD => SYNC(3), A => \SYNC_c[3]\);
    
    \VDB_pad_0[0]\ : BFR
      port map(A => \VDB_in[0]\, Y => \VDB_in_0[0]\);
    
    \SP_PDL_pad[15]\ : IOB33PH
      port map(PAD => SP_PDL(15), A => \I3.P0[15]\, EN => 
        MD_PDL_c_1, Y => \SP_PDL_in[15]\);
    
    \LB_pad[10]\ : IOB33PH
      port map(PAD => LB(10), A => \I2.LB_i[10]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[10]\);
    
    \LB_pad[23]\ : IOB33PH
      port map(PAD => LB(23), A => \I2.LB_i[23]\, EN => 
        \I2.LB_nOE_i_0_1\, Y => \LB_in[23]\);
    
    SCLK_PDL_pad : OB33PH
      port map(PAD => SCLK_PDL, A => SCLK_PDL_c);
    
    \TST_pad[4]\ : OB33PH
      port map(PAD => TST(4), A => \TST_c[4]\);
    
    \LB_pad[4]\ : IOB33PH
      port map(PAD => LB(4), A => \I2.LB_i[4]\, EN => 
        \I2.LB_nOE_i_0\, Y => \LB_in[4]\);
    
    \LB_pad[18]\ : IOB33PH
      port map(PAD => LB(18), A => \I2.LB_i[18]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[18]\);
    
    \SP_PDL_pad[5]\ : IOB33PH
      port map(PAD => SP_PDL(5), A => \I3.P0[5]\, EN => MD_PDL_c, 
        Y => \SP_PDL_in[5]\);
    
    \LB_pad[19]\ : IOB33PH
      port map(PAD => LB(19), A => \I2.LB_i[19]\, EN => 
        \I2.LB_nOE_i_0_0\, Y => \LB_in[19]\);
    

end DEF_ARCH; 
