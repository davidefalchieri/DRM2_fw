-- Version: 8.3 8.3.0.22

library ieee;
use ieee.std_logic_1164.all;
library APA;
use APA.all;

entity V1390trm is

    port( AMB          : in    std_logic_vector(5 downto 0);
          ASB          : in    std_logic;
          BERRVME      : in    std_logic;
          BNC_RESIN    : in    std_logic;
          CHAINA_ERR   : in    std_logic;
          CHAINB_ERR   : in    std_logic;
          CLK          : in    std_logic;
          COM_SER      : in    std_logic;
          DPR          : in    std_logic_vector(31 downto 0);
          DPR_P        : in    std_logic;
          DS0B         : in    std_logic;
          DS1B         : in    std_logic;
          EF           : in    std_logic;
          EV_RESIN     : in    std_logic;
          F_SO         : in    std_logic;
          GA           : in    std_logic_vector(4 downto 0);
          IACKB        : in    std_logic;
          IACKINB      : in    std_logic;
          INT_ERRA     : in    std_logic;
          INT_ERRB     : in    std_logic;
          L0           : in    std_logic;
          L1A          : in    std_logic;
          L1R          : in    std_logic;
          L2A          : in    std_logic;
          L2R          : in    std_logic;
          MROK         : in    std_logic;
          MSERCLK      : in    std_logic;
          MTDIA        : in    std_logic;
          MWOK         : in    std_logic;
          NPWON        : in    std_logic;
          PAE          : in    std_logic;
          PAF          : in    std_logic;
          SYSRESB      : in    std_logic;
          TDCDA        : in    std_logic_vector(31 downto 0);
          TDCDB        : in    std_logic_vector(31 downto 0);
          TDCDRYA      : in    std_logic;
          TDCDRYB      : in    std_logic;
          TOKOUTA      : in    std_logic;
          TOKOUTA_BP   : in    std_logic;
          TOKOUTB      : in    std_logic;
          TOKOUTB_BP   : in    std_logic;
          WRITEB       : in    std_logic;
          ff           : in    std_logic;
          ADE          : out   std_logic_vector(15 downto 0);
          ADLTC        : out   std_logic;
          ADO          : out   std_logic_vector(15 downto 0);
          BNC_RES      : out   std_logic;
          CHAINA_EN244 : out   std_logic;
          CHAINB_EN244 : out   std_logic;
          EV_RES       : out   std_logic;
          FCS          : out   std_logic;
          FID          : out   std_logic_vector(31 downto 0);
          FID_P        : out   std_logic;
          F_SCK        : out   std_logic;
          F_SI         : out   std_logic;
          IACKOUTB     : out   std_logic;
          INTR1        : out   std_logic;
          INTR2        : out   std_logic;
          LED_G        : out   std_logic;
          LED_R        : out   std_logic;
          MTDCRESA     : out   std_logic;
          MTDCRESB     : out   std_logic;
          MYBERR       : out   std_logic;
          NDTKIN       : out   std_logic;
          NLD          : out   std_logic;
          NMRSFIF      : out   std_logic;
          NOE16R       : out   std_logic;
          NOE16W       : out   std_logic;
          NOE32R       : out   std_logic;
          NOE32W       : out   std_logic;
          NOE64R       : out   std_logic;
          NOEAD        : out   std_logic;
          NOEDTK       : out   std_logic;
          NOELUT       : out   std_logic;
          NOEMIC       : out   std_logic;
          NOESRAME     : out   std_logic;
          NOESRAMO     : out   std_logic;
          NPRSFIF      : out   std_logic;
          NRDMEB       : out   std_logic;
          NWEN         : out   std_logic;
          NWRLUT       : out   std_logic;
          NWRSRAME     : out   std_logic;
          NWRSRAMO     : out   std_logic;
          NWRSRAM_TST  : out   std_logic;
          RAMAD        : out   std_logic_vector(17 downto 0);
          RMIC         : out   std_logic;
          SCLA         : out   std_logic;
          SCLB         : out   std_logic;
          STBMIC       : out   std_logic;
          TDCGDA       : out   std_logic;
          TDCGDB       : out   std_logic;
          TDCTRG       : out   std_logic;
          TDC_RESA     : out   std_logic;
          TDC_RESB     : out   std_logic;
          TOKINA       : out   std_logic;
          TOKINB       : out   std_logic;
          TRM_BUSY     : out   std_logic;
          TRM_DRDY     : out   std_logic;
          WMIC         : out   std_logic;
          SP0          : out   std_logic;
          SP1          : out   std_logic;
          SP2          : out   std_logic;
          SP3          : out   std_logic;
          SP4          : out   std_logic;
          SP5          : out   std_logic;
          DTE          : inout std_logic_vector(31 downto 0) := (others => 'Z');
          DTO          : inout std_logic_vector(31 downto 0) := (others => 'Z');
          LWORDB       : inout std_logic := 'Z';
          RAMDT        : inout std_logic_vector(13 downto 0) := (others => 'Z');
          SDAA         : inout std_logic := 'Z';
          SDAB         : inout std_logic := 'Z';
          VAD          : inout std_logic_vector(31 downto 1) := (others => 'Z');
          VDB          : inout std_logic_vector(31 downto 0) := (others => 'Z')
        );

end V1390trm;

architecture DEF_ARCH of V1390trm is 

  component MUX2L
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component BFR
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MUX2H
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IB33
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFF
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component LD
    port( EN : in    std_logic := 'U';
          D  : in    std_logic := 'U';
          Q  : out   std_logic
        );
  end component;

  component OB33PH
    port( PAD : out   std_logic;
          A   : in    std_logic := 'U'
        );
  end component;

  component NAND3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FFT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOB33PH
    port( PAD : inout   std_logic;
          A   : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component OAI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2FT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI21FTT
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GL33
    port( PAD : in    std_logic := 'U';
          GL  : out   std_logic
        );
  end component;

  component RAM256x9SST
    generic (MEMORYFILE:string := "");

    port( DO8    : out   std_logic;
          DO7    : out   std_logic;
          DO6    : out   std_logic;
          DO5    : out   std_logic;
          DO4    : out   std_logic;
          DO3    : out   std_logic;
          DO2    : out   std_logic;
          DO1    : out   std_logic;
          DO0    : out   std_logic;
          WPE    : out   std_logic;
          RPE    : out   std_logic;
          DOS    : out   std_logic;
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          DI8    : in    std_logic := 'U';
          DI7    : in    std_logic := 'U';
          DI6    : in    std_logic := 'U';
          DI5    : in    std_logic := 'U';
          DI4    : in    std_logic := 'U';
          DI3    : in    std_logic := 'U';
          DI2    : in    std_logic := 'U';
          DI1    : in    std_logic := 'U';
          DI0    : in    std_logic := 'U';
          WRB    : in    std_logic := 'U';
          RDB    : in    std_logic := 'U';
          WBLKB  : in    std_logic := 'U';
          RBLKB  : in    std_logic := 'U';
          PARODD : in    std_logic := 'U';
          WCLKS  : in    std_logic := 'U';
          RCLKS  : in    std_logic := 'U';
          DIS    : in    std_logic := 'U'
        );
  end component;

  component PLLCORE
    port( SDOUT    : out   std_logic;
          SCLK     : in    std_logic := 'U';
          SDIN     : in    std_logic := 'U';
          SSHIFT   : in    std_logic := 'U';
          SUPDATE  : in    std_logic := 'U';
          GLB      : out   std_logic;
          CLK      : in    std_logic := 'U';
          GLA      : out   std_logic;
          CLKA     : in    std_logic := 'U';
          LOCK     : out   std_logic;
          MODE     : in    std_logic := 'U';
          FBDIV5   : in    std_logic := 'U';
          EXTFB    : in    std_logic := 'U';
          FBSEL0   : in    std_logic := 'U';
          FBSEL1   : in    std_logic := 'U';
          FINDIV0  : in    std_logic := 'U';
          FINDIV1  : in    std_logic := 'U';
          FINDIV2  : in    std_logic := 'U';
          FINDIV3  : in    std_logic := 'U';
          FINDIV4  : in    std_logic := 'U';
          FBDIV0   : in    std_logic := 'U';
          FBDIV1   : in    std_logic := 'U';
          FBDIV2   : in    std_logic := 'U';
          FBDIV3   : in    std_logic := 'U';
          FBDIV4   : in    std_logic := 'U';
          STATBSEL : in    std_logic := 'U';
          DLYB0    : in    std_logic := 'U';
          DLYB1    : in    std_logic := 'U';
          OBDIV0   : in    std_logic := 'U';
          OBDIV1   : in    std_logic := 'U';
          STATASEL : in    std_logic := 'U';
          DLYA0    : in    std_logic := 'U';
          DLYA1    : in    std_logic := 'U';
          OADIV0   : in    std_logic := 'U';
          OADIV1   : in    std_logic := 'U';
          OAMUX0   : in    std_logic := 'U';
          OAMUX1   : in    std_logic := 'U';
          OBMUX0   : in    std_logic := 'U';
          OBMUX1   : in    std_logic := 'U';
          OBMUX2   : in    std_logic := 'U';
          FBDLY0   : in    std_logic := 'U';
          FBDLY1   : in    std_logic := 'U';
          FBDLY2   : in    std_logic := 'U';
          FBDLY3   : in    std_logic := 'U';
          XDLYSEL  : in    std_logic := 'U'
        );
  end component;

  component AOI21TTF
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFFLC
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OTB33PH
    port( PAD : out   std_logic;
          A   : in    std_logic := 'U';
          EN  : in    std_logic := 'U'
        );
  end component;

  component PWR
    port( Y : out   std_logic
        );
  end component;

  component RAM256x9SA
    generic (MEMORYFILE:string := "");

    port( DO8    : out   std_logic;
          DO7    : out   std_logic;
          DO6    : out   std_logic;
          DO5    : out   std_logic;
          DO4    : out   std_logic;
          DO3    : out   std_logic;
          DO2    : out   std_logic;
          DO1    : out   std_logic;
          DO0    : out   std_logic;
          WPE    : out   std_logic;
          RPE    : out   std_logic;
          DOS    : out   std_logic;
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          DI8    : in    std_logic := 'U';
          DI7    : in    std_logic := 'U';
          DI6    : in    std_logic := 'U';
          DI5    : in    std_logic := 'U';
          DI4    : in    std_logic := 'U';
          DI3    : in    std_logic := 'U';
          DI2    : in    std_logic := 'U';
          DI1    : in    std_logic := 'U';
          DI0    : in    std_logic := 'U';
          WRB    : in    std_logic := 'U';
          RDB    : in    std_logic := 'U';
          WBLKB  : in    std_logic := 'U';
          RBLKB  : in    std_logic := 'U';
          PARODD : in    std_logic := 'U';
          WCLKS  : in    std_logic := 'U';
          DIS    : in    std_logic := 'U'
        );
  end component;

  component DFFLB
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFFLS
    port( CLK : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          SET : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFFCI
    port( CLK  : in    std_logic := 'U';
          D    : in    std_logic := 'U';
          CLR  : in    std_logic := 'U';
          QBAR : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal PULSEl1r, PULSEl2r, PULSEl3r, PULSEl4r, PULSEl5r, 
        PULSEl6r, PULSEl7r, PULSEl8r, PULSEl9r, TICKl0r, 
        CLEAR_STAT, FLUSH, END_FLUSH, LSRAM_FL_RD, END_TDC, 
        LEAD_FLAGl0r, LEAD_FLAGl1r, LEAD_FLAGl2r, LEAD_FLAGl3r, 
        LEAD_FLAGl4r, LEAD_FLAGl5r, LEAD_FLAGl6r, LEAD_FLAGl7r, 
        COM_SERS, LOAD_RES, PLL_LOCK, HWCLEAR, BNC_RES_E, EVREAD, 
        DTEST_FIFO, RAMAD_VMEl0r, RAMAD_VMEl1r, RAMAD_VMEl2r, 
        RAMAD_VMEl3r, RAMAD_VMEl4r, RAMAD_VMEl5r, RAMAD_VMEl6r, 
        RAMAD_VMEl7r, RAMAD_VMEl8r, RAMAD_VMEl9r, RAMAD_VMEl10r, 
        RAMAD_VMEl11r, RAMAD_VMEl12r, RAMAD_VMEl13r, 
        RAMAD_VMEl14r, RAMAD_VMEl15r, RAMAD_VMEl16r, 
        RAMAD_VMEl17r, REGl26r, REGl27r, REGl32r, REGl33r, 
        REGl34r, REGl35r, REGl36r, REGl37r, REGl38r, REGl39r, 
        REGl40r, REGl41r, REGl43r, REGl44r, REGl45r, REGl46r, 
        REGl47r, REGl48r, REGl49r, REGl50r, REGl51r, REGl52r, 
        REGl53r, REGl54r, REGl55r, REGl56r, REGl57r, REGl58r, 
        REGl59r, REGl60r, REGl61r, REGl62r, REGl63r, REGl64r, 
        REGl65r, REGl66r, REGl67r, REGl68r, REGl69r, REGl70r, 
        REGl71r, REGl72r, REGl73r, REGl74r, REGl75r, REGl76r, 
        REGl77r, REGl78r, REGl79r, REGl80r, REGl81r, REGl82r, 
        REGl83r, REGl84r, REGl85r, REGl86r, REGl87r, REGl88r, 
        REGl89r, REGl90r, REGl101r, REGl102r, REGl103r, REGl109r, 
        REGl110r, REGl111r, REGl112r, REGl113r, REGl114r, 
        REGl115r, REGl116r, REGl117r, REGl118r, REGl125r, 
        REGl126r, REGl127r, REGl128r, REGl129r, REGl130r, 
        REGl131r, REGl132r, REGl406r, REGl407r, REGl408r, 
        REGl409r, REGl410r, REGl411r, REGl412r, REGl413r, 
        REGl414r, REGl415r, REGl416r, REGl417r, REGl418r, 
        REGl419r, REGl420r, REGl421r, REGl422r, REGl423r, 
        REGl424r, REGl425r, REGl426r, REGl427r, REGl428r, 
        REGl429r, REGl430r, REGl431r, REGl434r, REGl435r, 
        REGl436r, REGl437r, REGl438r, REGl439r, REGl440r, 
        REGl441r, REGl442r, REGl443r, REGl444r, REGl445r, 
        REGl446r, REGl447r, \I3.REG1l3r_net_1\, 
        \I3.REG2l3r_net_1\, \I3.VADml0r\, \I3.VADml1r\, 
        \I3.VADml2r\, \I3.VADml3r\, \I3.VADml4r\, \I3.VADml5r\, 
        \I3.VADml6r\, \I3.VADml7r\, \I3.VADml8r\, \I3.VADml9r\, 
        \I3.VADml10r\, \I3.VADml11r\, \I3.VADml12r\, 
        \I3.VADml13r\, \I3.VADml14r\, \I3.VADml15r\, 
        \I3.VADml16r\, \I3.VADml17r\, \I3.VADml18r\, 
        \I3.VADml19r\, \I3.VADml20r\, \I3.VADml21r\, 
        \I3.VADml22r\, \I3.VADml23r\, \I3.VADml24r\, 
        \I3.VADml25r\, \I3.VADml26r\, \I3.VADml27r\, 
        \I3.VADml28r\, \I3.VADml29r\, \I3.VADml30r\, 
        \I3.VADml31r\, \I3.REG3l3r_net_1\, \I3.VDBml0r_net_1\, 
        \I3.VDBml1r_net_1\, \I3.VDBml2r_net_1\, 
        \I3.VDBml3r_net_1\, \I3.VDBml4r_net_1\, 
        \I3.VDBml6r_net_1\, \I3.VDBml8r_net_1\, 
        \I3.VDBml9r_net_1\, \I3.VDBml10r_net_1\, 
        \I3.VDBml11r_net_1\, \I3.VDBml12r_net_1\, 
        \I3.VDBml13r_net_1\, \I3.VDBml14r_net_1\, 
        \I3.VDBml15r_net_1\, \I3.VDBml16r_net_1\, 
        \I3.VDBml17r_net_1\, \I3.VDBml18r_net_1\, 
        \I3.VDBml19r_net_1\, \I3.VDBml20r_net_1\, 
        \I3.VDBml21r_net_1\, \I3.VDBml22r_net_1\, 
        \I3.VDBml23r_net_1\, \I3.VDBml24r_net_1\, 
        \I3.VDBml25r_net_1\, \I3.VDBml26r_net_1\, 
        \I3.VDBml27r_net_1\, \I3.VDBml28r_net_1\, 
        \I3.VDBml29r_net_1\, \I3.VDBml30r_net_1\, 
        \I3.VDBml31r_net_1\, \I3.N_11\, VDBm_i_i_m2l5r, 
        LED_R_i_a3, \I1.RAMDT_SPI_e_net_1\, 
        \I1.RAMDT_SPI_1l0r_net_1\, \I1.RAMDT_SPI_1l1r_net_1\, 
        \I1.RAMDT_SPI_1l2r_net_1\, \I1.RAMDT_SPI_1l3r_net_1\, 
        \I1.RAMDT_SPI_1l4r_net_1\, \I1.RAMDT_SPI_1l5r_net_1\, 
        \I1.RAMDT_SPI_1l6r_net_1\, \I2.DTE_cll31r\, 
        \I2.DTO_cl_32l31r\, \I2.DTO_cll31r\, \I2.DTE_cl_32l31r\, 
        \I2.DTE_1l0r_net_1\, \I2.DTE_1l1r_net_1\, 
        \I2.DTE_1l2r_net_1\, \I2.DTE_1l3r_net_1\, 
        \I2.DTE_1l5r_net_1\, \I2.DTE_1l29r_net_1\, 
        \I2.DTE_1l30r_net_1\, \I2.DTE_1l31r_net_1\, 
        \I2.CHAINA_EN244_i\, un1_sdaa_0_a2, un1_sdab_0_a2, 
        \I5.SDAout_net_1\, \I5.N_106\, \I5.N_107\, AMB_cl0r, 
        AMB_cl1r, AMB_cl2r, AMB_cl3r, AMB_cl4r, ASB_c, 
        BNC_RESIN_c, CHAINA_ERR_c, CHAINB_ERR_c, CLK_c, COM_SER_c, 
        DPR_cl0r, DPR_cl1r, DPR_cl2r, DPR_cl3r, DPR_cl4r, 
        DPR_cl5r, DPR_cl6r, DPR_cl7r, DPR_cl8r, DPR_cl9r, 
        DPR_cl10r, DPR_cl11r, DPR_cl12r, DPR_cl13r, DPR_cl14r, 
        DPR_cl15r, DPR_cl16r, DPR_cl17r, DPR_cl18r, DPR_cl19r, 
        DPR_cl20r, DPR_cl21r, DPR_cl22r, DPR_cl23r, DPR_cl24r, 
        DPR_cl25r, DPR_cl26r, DPR_cl27r, DPR_cl28r, DPR_cl29r, 
        DPR_cl30r, DPR_cl31r, DS0B_c, DS1B_c, EF_c, EV_RESIN_c, 
        F_SO_c, GA_cl0r, GA_cl1r, GA_cl2r, GA_cl3r, IACKB_c, 
        INT_ERRA_c, INT_ERRB_c, L1A_c, L2A_c, L2R_c, MROK_c, 
        MSERCLK_c, MTDIA_c, MWOK_c, NPWON_c, PAF_c, SYSRESB_c, 
        TDCDA_cl0r, TDCDA_cl1r, TDCDA_cl2r, TDCDA_cl3r, 
        TDCDA_cl4r, TDCDA_cl5r, TDCDA_cl6r, TDCDA_cl7r, 
        TDCDA_cl8r, TDCDA_cl9r, TDCDA_cl10r, TDCDA_cl11r, 
        TDCDA_cl12r, TDCDA_cl13r, TDCDA_cl14r, TDCDA_cl15r, 
        TDCDA_cl16r, TDCDA_cl17r, TDCDA_cl18r, TDCDA_cl19r, 
        TDCDA_cl20r, TDCDA_cl21r, TDCDA_cl22r, TDCDA_cl23r, 
        TDCDA_cl24r, TDCDA_cl25r, TDCDA_cl26r, TDCDA_cl27r, 
        TDCDA_cl28r, TDCDA_cl29r, TDCDA_cl30r, TDCDA_cl31r, 
        TDCDB_cl0r, TDCDB_cl1r, TDCDB_cl2r, TDCDB_cl3r, 
        TDCDB_cl4r, TDCDB_cl5r, TDCDB_cl6r, TDCDB_cl7r, 
        TDCDB_cl8r, TDCDB_cl9r, TDCDB_cl10r, TDCDB_cl11r, 
        TDCDB_cl12r, TDCDB_cl13r, TDCDB_cl14r, TDCDB_cl15r, 
        TDCDB_cl16r, TDCDB_cl17r, TDCDB_cl18r, TDCDB_cl19r, 
        TDCDB_cl20r, TDCDB_cl21r, TDCDB_cl22r, TDCDB_cl23r, 
        TDCDB_cl24r, TDCDB_cl25r, TDCDB_cl26r, TDCDB_cl27r, 
        TDCDB_cl28r, TDCDB_cl29r, TDCDB_cl30r, TDCDB_cl31r, 
        TDCDRYA_c, TDCDRYB_c, TOKOUTA_c, TOKOUTA_BP_c, TOKOUTB_c, 
        TOKOUTB_BP_c, WRITEB_c, ADE_cl0r, ADE_cl1r, ADE_cl2r, 
        ADE_cl3r, ADE_cl4r, ADE_cl5r, ADE_cl6r, ADE_cl7r, 
        ADE_cl8r, ADE_cl9r, ADE_cl10r, ADE_cl11r, ADE_cl12r, 
        ADE_cl13r, ADE_cl14r, ADE_cl15r, ADO_cl0r, ADO_cl1r, 
        ADO_cl2r, ADO_cl3r, ADO_cl4r, ADO_cl5r, ADO_cl6r, 
        ADO_cl7r, ADO_cl8r, ADO_cl9r, ADO_cl10r, ADO_cl11r, 
        ADO_cl12r, ADO_cl13r, ADO_cl14r, ADO_cl15r, BNC_RES_c, 
        EV_RES_c, FID_cl0r, FID_cl1r, FID_cl2r, FID_cl3r, 
        FID_cl4r, FID_cl5r, FID_cl6r, FID_cl7r, FID_cl8r, 
        FID_cl9r, FID_cl10r, FID_cl11r, FID_cl12r, FID_cl13r, 
        FID_cl14r, FID_cl15r, FID_cl16r, FID_cl17r, FID_cl18r, 
        FID_cl19r, FID_cl20r, FID_cl21r, FID_cl22r, FID_cl23r, 
        FID_cl24r, FID_cl25r, FID_cl26r, FID_cl27r, FID_cl28r, 
        FID_cl29r, FID_cl30r, FID_cl31r, F_SI_c, \VCC\, LED_G_c, 
        MTDCRESA_c, MTDCRESB_c, MYBERR_c, NDTKIN_c, NLD_c, 
        NOE16R_c, NOE32R_c, NOEDTK_c, NOELUT_c, NOEMIC_c, 
        NOESRAME_c, NOESRAMO_c, NMRSFIF_c_c, NRDMEB_c, NWEN_c, 
        NWRLUT_c, NWRSRAME_c, NWRSRAMO_c, NWRSRAM_TST_c, 
        RAMAD_cl0r, RAMAD_cl1r, RAMAD_cl2r, RAMAD_cl3r, 
        RAMAD_cl4r, RAMAD_cl5r, RAMAD_cl6r, RAMAD_cl7r, 
        RAMAD_cl8r, RAMAD_cl9r, RAMAD_cl10r, RAMAD_cl11r, 
        RAMAD_cl12r, RAMAD_cl13r, RAMAD_cl14r, RAMAD_cl15r, 
        RAMAD_cl16r, RAMAD_cl17r, RMIC_c, STBMIC_c, TDCGDA_c, 
        TDCGDB_c, TDCTRG_c, TDC_RES_c_c, TOKINA_c, TOKINB_c, 
        TRM_BUSY_c, EVRDY_c, WMIC_c, DTE_inl0r, DTE_inl1r, 
        DTE_inl2r, DTE_inl3r, DTE_inl4r, DTE_inl5r, DTE_inl6r, 
        DTE_inl7r, DTE_inl8r, DTE_inl9r, DTE_inl10r, DTE_inl11r, 
        DTE_inl12r, DTE_inl13r, DTE_inl14r, DTE_inl15r, 
        DTE_inl16r, DTE_inl17r, DTE_inl18r, DTE_inl19r, 
        DTE_inl20r, DTE_inl21r, DTE_inl22r, DTE_inl23r, 
        DTE_inl24r, DTE_inl25r, DTE_inl26r, DTE_inl27r, 
        DTE_inl28r, DTE_inl29r, DTE_inl30r, DTE_inl31r, DTO_inl0r, 
        DTO_inl1r, DTO_inl2r, DTO_inl3r, DTO_inl4r, DTO_inl5r, 
        DTO_inl6r, DTO_inl7r, DTO_inl8r, DTO_inl9r, DTO_inl10r, 
        DTO_inl11r, DTO_inl12r, DTO_inl13r, DTO_inl14r, 
        DTO_inl15r, DTO_inl16r, DTO_inl17r, DTO_inl18r, 
        DTO_inl19r, DTO_inl20r, DTO_inl21r, DTO_inl22r, 
        DTO_inl23r, DTO_inl24r, DTO_inl25r, DTO_inl26r, 
        DTO_inl27r, DTO_inl28r, DTO_inl29r, DTO_inl30r, 
        DTO_inl31r, LWORDB_in, RAMDT_inl0r, RAMDT_inl1r, 
        RAMDT_inl2r, RAMDT_inl3r, RAMDT_inl4r, RAMDT_inl5r, 
        RAMDT_inl6r, RAMDT_inl7r, RAMDT_inl8r, RAMDT_inl9r, 
        RAMDT_inl10r, RAMDT_inl11r, RAMDT_inl12r, RAMDT_inl13r, 
        SDAA_in, SDAB_in, \GND\, VAD_inl1r, VAD_inl2r, VAD_inl3r, 
        VAD_inl4r, VAD_inl5r, VAD_inl6r, VAD_inl7r, VAD_inl8r, 
        VAD_inl9r, VAD_inl10r, VAD_inl11r, VAD_inl12r, VAD_inl13r, 
        VAD_inl14r, VAD_inl15r, VAD_inl28r, VAD_inl29r, 
        VAD_inl30r, VAD_inl31r, VDB_inl0r, VDB_inl1r, VDB_inl2r, 
        VDB_inl3r, VDB_inl4r, VDB_inl5r, VDB_inl6r, VDB_inl7r, 
        VDB_inl8r, VDB_inl9r, VDB_inl10r, VDB_inl11r, VDB_inl12r, 
        VDB_inl13r, VDB_inl14r, VDB_inl15r, VDB_inl16r, 
        VDB_inl17r, VDB_inl18r, VDB_inl19r, VDB_inl20r, 
        VDB_inl21r, VDB_inl22r, VDB_inl23r, VDB_inl24r, 
        VDB_inl25r, VDB_inl26r, VDB_inl27r, VDB_inl28r, 
        VDB_inl29r, VDB_inl30r, VDB_inl31r, NPWON_c_i_0, 
        REG_i_0_il42r, PAF_c_i_0, NOE32R_c_i_0, AMB_c_i_0_il5r, 
        \I2.N_4239_i_0_1\, \I2.N_4178_i_0_1\, \I1.RAMDT_SPI_E_0\, 
        \I3.un1_vdb_0\, LOAD_RES_1, TICKL0R_2, TICKL0R_3, 
        \I5.SENS_ADDR_1_sqmuxa_1_0_net_1\, \I5.sstate1l13r_net_1\, 
        \I5.sstate1_ns_el0r\, \I5.AIR_CHAIN_net_1\, 
        \I5.sstate2l0r_net_1\, \I5.COMMANDl0r_net_1\, 
        \I5.sstate1l11r_net_1\, \I5.REG_1_sqmuxa_0_net_1\, 
        \I5.DWACT_ADD_CI_0_g_array_1l0r\, 
        \I5.DWACT_ADD_CI_0_TMPl0r\, \I5.SENS_ADDRl1r_net_1\, 
        \I5.SCL_net_1\, \I5.CHAIN_SELECT_net_1\, 
        \I5.sstate1l12r_net_1\, \I5.sstate1l6r_net_1\, 
        \I5.sstate1l7r_net_1\, \I5.sstate1l1r_net_1\, 
        \I5.sstate2se_2_i_net_1\, \I5.sstate2l2r_net_1\, 
        \I5.sstate2l1r_net_1\, \I5.sstate2se_3_i_net_1\, 
        \I5.sstate2_ns_el2r\, \I5.sstate2_ns_el1r\, 
        \I5.sstate2l4r_net_1\, \I5.sstate2l3r_net_1\, 
        \I5.sstate2_ns_el0r\, \I5.sstate2_5_sqmuxa\, 
        \I5.sstate1l0r_net_1\, \I5.sstate1l5r_net_1\, 
        \I5.sstate1_ns_el8r\, \I5.N_130\, \I5.sstate1l8r_net_1\, 
        \I5.sstate1_ns_el5r\, \I5.sstate1_ns_el1r\, \I5.N_64\, 
        \I5.COMMANDl1r_net_1\, \I5.COMMANDl2r_net_1\, 
        \I5.PULSE_FL_net_1\, \I5.BITCNT_86_net_1\, \I5.BITCNT_c0\, 
        \I5.N_50\, \I5.BITCNTe\, \I5.N_94\, \I5.N_144\, 
        \I5.BITCNT_85_net_1\, \I5.BITCNTl1r_net_1\, \I5.N_52\, 
        \I5.BITCNT_84_net_1\, \I5.BITCNTl2r_net_1\, \I5.N_75\, 
        \I5.N_71\, \I5.SDAnoe_83_net_1\, \I5.SDAnoe_net_1\, 
        \I5.SDAnoe_8\, \I5.SDAout_82_net_1\, \I5.SDAout_12\, 
        \I5.N_150\, \I5.COMMANDl15r_net_1\, \I5.SBYTEl7r_net_1\, 
        \I5.TEMPDATA_81_net_1\, \I5.TEMPDATAl7r_net_1\, 
        \I5.N_443\, \I5.TEMPDATA_80_net_1\, 
        \I5.TEMPDATAl6r_net_1\, \I5.TEMPDATA_79_net_1\, 
        \I5.TEMPDATAl5r_net_1\, \I5.TEMPDATA_78_net_1\, 
        \I5.TEMPDATAl4r_net_1\, \I5.TEMPDATA_77_net_1\, 
        \I5.TEMPDATAl3r_net_1\, \I5.TEMPDATA_76_net_1\, 
        \I5.TEMPDATAl2r_net_1\, \I5.TEMPDATA_75_net_1\, 
        \I5.TEMPDATAl1r_net_1\, \I5.TEMPDATA_74_net_1\, 
        \I5.TEMPDATAl0r_net_1\, \I5.TEMP_ACK_73_net_1\, 
        \I5.TEMP_ACK_net_1\, \I5.SBYTE_72_net_1\, \I5.SBYTE_9l7r\, 
        \I5.N_406\, \I5.SBYTEl6r_net_1\, \I5.SBYTE_71_net_1\, 
        \I5.N_26\, \I5.COMMANDl14r_net_1\, \I5.SBYTEl5r_net_1\, 
        \I5.SBYTE_70_net_1\, \I5.N_24\, \I5.COMMANDl13r_net_1\, 
        \I5.SBYTEl4r_net_1\, \I5.SBYTE_69_net_1\, \I5.N_22\, 
        \I5.COMMANDl12r_net_1\, \I5.SBYTEl3r_net_1\, 
        \I5.SBYTE_68_net_1\, \I5.N_20\, \I5.COMMANDl11r_net_1\, 
        \I5.SBYTEl2r_net_1\, \I5.SBYTE_67_net_1\, \I5.N_18\, 
        \I5.COMMANDl10r_net_1\, \I5.SBYTEl1r_net_1\, 
        \I5.SBYTE_66_net_1\, \I5.N_16\, \I5.COMMANDl9r_net_1\, 
        \I5.SBYTEl0r_net_1\, \I5.SBYTE_65_net_1\, \I5.SBYTE_9l0r\, 
        \I5.COMMANDl8r_net_1\, \I5.N_101\, 
        \I5.AIR_PULSE_64_net_1\, \I5.AIR_PULSE_net_1\, 
        \I5.AIR_PULSE_3_net_1\, \I5.N_459\, 
        \I5.un1_sstate2_3_0_net_1\, \I5.AIR_START_net_1\, 
        \I5.SCL_63_net_1\, \I5.N_484\, \I5.N_82\, 
        \I5.AIR_WDATA_62_net_1\, \I5.AIR_WDATAl15r_net_1\, 
        \I5.N_461\, \I5.AIR_WDATA_61_net_1\, 
        \I5.AIR_WDATAl11r_net_1\, \I5.SENS_ADDRl2r_net_1\, 
        \I5.AIR_WDATA_60_net_1\, \I5.AIR_WDATAl10r_net_1\, 
        \I5.AIR_WDATA_59_net_1\, \I5.AIR_WDATAl9r_net_1\, 
        \I5.SENS_ADDRl0r_net_1\, \I5.AIR_WDATA_58_net_1\, 
        \I5.AIR_WDATAl8r_net_1\, \I5.AIR_WDATA_57_net_1\, 
        \I5.AIR_WDATAl2r_net_1\, \I5.AIR_WDATA_56_net_1\, 
        \I5.AIR_WDATAl1r_net_1\, \I5.AIR_WDATA_55_net_1\, 
        \I5.AIR_WDATAl0r_net_1\, \I5.REG_1_54_net_1\, 
        \I5.PULSE_FL_53_net_1\, \I5.COMMAND_52_net_1\, 
        \I5.COMMAND_51_net_1\, \I5.COMMAND_50_net_1\, 
        \I5.COMMAND_49_net_1\, \I5.COMMAND_48_net_1\, 
        \I5.SSTATE1L13R_4\, \I5.COMMAND_47_net_1\, 
        \I5.COMMAND_46_net_1\, \I5.COMMAND_45_net_1\, 
        \I5.REG_1_44_net_1\, \I5.REG_1_43_net_1\, 
        \I5.REG_1_42_net_1\, \I5.REG_1_41_net_1\, 
        \I5.REG_1_40_net_1\, \I5.REG_1_39_net_1\, 
        \I5.REG_1_38_net_1\, \I5.REG_1_37_net_1\, 
        \I5.REG_1_36_net_1\, \I5.REG_1_35_net_1\, 
        \I5.REG_1_34_net_1\, \I5.REG_1_33_net_1\, 
        \I5.REG_1_32_net_1\, \I5.REG_1_31_net_1\, 
        \I5.REG_1_30_net_1\, \I5.REG_1_29_net_1\, 
        \I5.REG_1_28_net_1\, \I5.REG_1_27_net_1\, 
        \I5.REG_1_26_net_1\, \I5.REG_1_25_net_1\, 
        \I5.REG_1_24_net_1\, \I5.REG_1_23_net_1\, 
        \I5.REG_1_22_net_1\, \I5.REG_1_21_net_1\, 
        \I5.REG_1_20_net_1\, \I5.REG_1_19_net_1\, 
        \I5.REG_1_18_net_1\, \I5.REG_1_17_net_1\, 
        \I5.AIR_CHAIN_15_net_1\, \I5.COMMAND_14_net_1\, 
        \I5.COMMAND_13_net_1\, \I5.COMMAND_12_net_1\, 
        \I5.CHAIN_SELECT_11_net_1\, \I5.DATA_12_ivl1r_net_1\, 
        \I5.SDAin_m_1_net_1\, \I5.SENS_ADDR_6l2r_net_1\, 
        \I5.SENS_ADDR_1_sqmuxa_net_1\, \I5.I_14\, 
        \I5.SENS_ADDR_6l0r_net_1\, 
        \I5.DWACT_ADD_CI_0_partial_suml0r\, \I5.I_13\, 
        \I4.STATE1l1r_net_1\, \I4.END_FLUSH_2_net_1\, 
        \I4.STATE1_nsl2r\, \I4.FLUSH_0_sqmuxa_net_1\, 
        \I4.STATE1_nsl1r_net_1\, \I4.STATE1_nsl0r_net_1\, 
        \I4.STATE1l2r_net_1\, \I4.STATE1l0r_net_1\, 
        \I4.LSRAM_FL_RD_4_net_1\, \I4.FLUSH_3_net_1\, 
        \I4.un1_FLUSH_1_sqmuxa_1_net_1\, \I0.un12_clear_i\, 
        \I0.CLEAR_STATi_4_net_1\, \I0.un4_hwresi_i\, 
        \I0.CLEARF1_net_1\, \I0.CLEAR_net_1\, \I0.CLEAR_i_0\, 
        \I0.REG_1_3_net_1\, \I0.TDC_RESi_1_net_1\, 
        \I0.COM_SERF1_net_1\, \I0.CLEARF2_i\, 
        \I0.BNC_RESF1_net_1\, \I0.EV_RESF1_net_1\, 
        \I0.BNC_RESF3_net_1\, \I2.GIROT_452\, \I2.GIROT_net_1\, 
        \I2.N_3760\, \I2.N_3794\, \I2.un9_tdctrgi_i_0\, 
        \I2.TRGCNT_n4\, \I2.N_3764\, \I2.TRGCNT_n4_0\, 
        \I2.TRGCNTl4r_net_1\, \I2.TRGCNT_i_0_il3r\, 
        \I2.TRGCNT_n3\, \I2.N_3763\, \I2.TRGCNT_n3_0\, 
        \I2.N_3796\, \I2.TRGCNTl2r_net_1\, \I2.TRGCNT_n2\, 
        \I2.N_3762\, \I2.TRGCNT_n2_0\, \I2.TRGCNT_i_0_il1r\, 
        \I2.TRGCNT_n1\, \I2.N_3761\, \I2.TRGCNT_n1_0\, 
        \I2.TRGCNTl0r_net_1\, \I2.STATE1l17r_net_1\, 
        \I2.LSRAM_RADDRi_501\, \I2.PIPE4_DTl23r_net_1\, 
        \I2.LSRAM_RADDRil2r_net_1\, \I2.N_4642\, 
        \I2.LSRAM_RADDRi_500\, \I2.PIPE4_DTl22r_net_1\, 
        \I2.LSRAM_RADDRil1r_net_1\, \I2.LSRAM_RADDRi_499\, 
        \I2.PIPE4_DTl21r_net_1\, \I2.LSRAM_RADDRil0r_net_1\, 
        \I2.N_4524\, \I2.TRAIL_MIS6_491\, \I2.N_4643\, 
        \I2.TRAIL_MIS6_net_1\, \I2.PIPE4_DTl30r_net_1\, 
        \I2.NWPIPE4_net_1\, \I2.NWPIPE5_net_1\, 
        \I2.PIPE4_DTl31r_net_1\, \I2.BITCNT_940\, \I2.BITCNT_c0\, 
        \I2.BITCNT_n0\, \I2.BITCNTe\, \I2.BITCNT_939\, 
        \I2.BITCNTl1r_net_1\, \I2.N_4322\, \I2.BITCNT_938\, 
        \I2.BITCNTl2r_net_1\, \I2.N_4323\, \I2.BITCNT_937\, 
        \I2.BITCNTl3r_net_1\, \I2.N_4324\, \I2.BITCNT_936\, 
        \I2.BITCNT_i_0_il4r\, \I2.N_4325\, 
        \I2.ERR_WORDS_RDY_0_sqmuxa\, \I2.BITCNT_935\, 
        \I2.BITCNTl5r_net_1\, \I2.N_4326\, \I2.FID_436\, 
        \I2.FID_7l20r\, \I2.FID_435\, \I2.FID_7l19r\, 
        \I2.FID_434\, \I2.FID_7l18r\, \I2.FID_433\, 
        \I2.FID_7l17r\, \I2.FID_432\, \I2.FID_7l16r\, 
        \I2.FID_431\, \I2.FID_7l15r\, \I2.FID_430\, 
        \I2.FID_7l14r\, \I2.FID_429\, \I2.FID_7l13r\, 
        \I2.FID_428\, \I2.FID_7l12r\, \I2.FID_427\, 
        \I2.FID_7l11r\, \I2.FID_426\, \I2.FID_7l10r\, 
        \I2.STATE3l7r_net_1\, \I2.FID_447\, \I2.FID_7l31r\, 
        \I2.FID_446\, \I2.FID_7l30r\, \I2.FID_445\, 
        \I2.FID_7l29r\, \I2.FID_444\, \I2.FID_7l28r\, 
        \I2.FID_443\, \I2.FID_7l27r\, \I2.FID_442\, 
        \I2.FID_7l26r\, \I2.FID_441\, \I2.FID_7l25r\, 
        \I2.FID_440\, \I2.FID_7l24r\, \I2.FID_439\, 
        \I2.FID_7l23r\, \I2.FID_438\, \I2.FID_7l22r\, 
        \I2.FID_437\, \I2.FID_7l21r\, \I2.N_2796_i_0\, 
        \I2.STATE2_nsl3r\, \I2.N_176_i\, \I2.PIPE7_DTl30r_net_1\, 
        \I2.PIPE7_DTl31r_net_1\, \I2.PIPE7_DT_i_0l33r\, 
        \I2.NWPIPE8_i_0_i_0_0\, \I2.CLK_tdc\, 
        \I2.STATE1_nsl6r_net_1\, \I2.NWPIPE3_net_1\, 
        \I2.NWPIPE6_net_1\, \I2.PIPE6_DTl24r_net_1\, 
        \I2.PIPE6_DTl25r_net_1\, \I2.PIPE6_DTl26r_net_1\, 
        \I2.PIPE6_DTl27r_net_1\, \I2.NWPIPE9_0_net_1\, 
        \I2.PIPE5_DT_698_net_1\, \I2.STATE2_nsl1r\, 
        \I2.STATE2_nsl2r\, \I2.STATE3_nsl10r_net_1\, 
        \I2.STATE3_ns_il11r_net_1\, \I2.STATE3_nsl6r_net_1\, 
        \I2.L2SERV_919_net_1\, \I2.N_154\, \I2.STATE1l2r_net_1\, 
        \I2.STATE1_ns_0l5r\, \I2.N_3287_i_0\, \I2.N_3888\, 
        \I2.CHAINB_EN244_c_0\, \I2.N_3279_0\, \I2.N_3280\, 
        \I2.STATE1l14r_net_1\, \I2.STATE1l4r_net_1\, 
        \I2.DTE_cl_0_sqmuxa_2_0\, 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_net_1\, 
        \I2.N_4241_1\, \I2.N_2870\, \I2.N_4282\, \I2.N_2868_1\, 
        \I2.N_237\, \I2.N_4641\, \I2.DTO_cl_0_sqmuxa_0\, 
        \I2.NWPIPE2_net_1\, \I2.N_2864_0\, \I2.N_4680_0\, 
        \I2.N_3965_0\, \I2.ROFFSET_0_sqmuxa_1\, \I2.N_12254_i\, 
        \I2.STATE3_nsl13r\, \I2.FIFO_END_EVNT_net_1\, 
        \I2.PIPE1_DT_42_3_0l28r\, \I2.N_12169_i\, 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\, 
        \I2.PIPE1_DT_42_0l27r_net_1\, \I2.TDCGDA1_net_1\, 
        \I2.END_CHAINA1_1_sqmuxa_3\, \I2.NWPIPE1_4_sqmuxa_1_0\, 
        \I2.FIRST_TDC_1_sqmuxa_net_1\, \I2.N_3798\, 
        \I2.PIPE1_DT_2_sqmuxa_1_1_net_1\, \I2.TDCGDB1_net_1\, 
        \I2.N_3879\, \I2.TDCDASl31r_net_1\, \I2.TDCDBSl31r_net_1\, 
        \I2.TDCDBSl29r_net_1\, \I2.N_3283\, \I2.N_4283_i_0\, 
        \I2.TEMPF_net_1\, \I2.N_2867_1\, 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, \I2.LEAD_FLAG6_0_sqmuxa\, 
        \I2.un1_NWPIPE5_1_i\, \I2.SUB9_0_sqmuxa_0\, 
        \I2.NWPIPE8_I_0_I_0_0_5\, \I2.PIPE8_DTl30r_net_1\, 
        \I2.N_4273\, \I2.CRC32_1_sqmuxa_0\, \I2.N_2838_i_0\, 
        \I2.SUB8_1_sqmuxa_0\, \I2.N_4482_0\, \I2.L2RF3_i\, 
        \I2.L2RF2_net_1\, \I2.DTE_0_sqmuxa_i_0_N_3_1\, 
        \I2.NWPIPE8_I_0_I_0_0_6\, \I2.WOFFSETl0r_net_1\, 
        \I2.N_4707_i_0\, \I2.TRGARRl1r_net_1\, 
        \I2.TRGARRl2r_net_1\, \I2.TRGSERVl2r_net_1\, \I2.N_45\, 
        \I2.BNC_IDl1r_net_1\, \I2.BNC_IDl0r_net_1\, \I2.N_37\, 
        \I2.BNC_IDl3r_net_1\, \I2.DWACT_FINC_El0r\, \I2.N_14\, 
        \I2.BNC_IDl8r_net_1\, \I2.DWACT_FINC_El4r\, \I2.N_50\, 
        \I2.N_42\, \I2.DWACT_FINC_E_0l0r\, \I2.N_19\, 
        \I2.DWACT_FINC_E_0l4r\, \I2.N_4\, \I2.PIPE6_DTl33r_net_1\, 
        \I2.L1AF2_net_1\, \I2.STATE4_ns_il2r_net_1\, 
        \I2.STATE4l2r_net_1\, \I2.N_3376_1\, \I2.STATE4l1r_net_1\, 
        \I2.STATE3l9r_net_1\, \I2.un12_clear_stat_i\, 
        \I2.TOKENTOB_RES_net_1\, \I2.un6_clear_stat_i\, 
        \I2.TOKENTOA_RES_net_1\, \I2.OFFSETl0r_net_1\, 
        \I2.STATEe_i_0l0r_net_1\, \I2.STATEe_illegalpipe2_net_1\, 
        \I2.N_3234_i_0\, \I2.N_3234\, \I2.N_4284\, 
        \I2.STATE2_ns_i_0_1_il0r\, \I2.STATE2l0r_net_1\, 
        \I2.STATE2l2r_net_1\, \I2.un8_hwres_i\, \I2.N_3206_i_0\, 
        \I2.N_3272\, \I2.N_3316\, \I2.N_3275\, 
        \I2.STATE1l10r_net_1\, \I2.N_3214_i_0\, \I2.N_3347_1\, 
        \I2.STATE1l5r_net_1\, \I2.N_4628_i_0\, \I2.N_4627_i_0\, 
        \I2.N_4625_i_0\, \I2.N_4620_i_0\, \I2.N_4618_i_0\, 
        \I2.N_4617_i_0\, \I2.N_4616_i_0\, \I2.N_4614_i_0\, 
        \I2.N_4611_i_0\, \I2.N_4608_i_0\, \I2.N_4607_i_0\, 
        \I2.N_4606_i_0\, \I2.N_3875_i_0\, \I2.N_3887\, 
        \I2.N_3208_i_0\, \I2.END_CHAINA1_net_1\, \I2.N_3288\, 
        \I2.STATE5_ns_il1r\, \I2.N_4338_1\, \I2.STATE5l3r_net_1\, 
        \I2.un9_clear_stat_i\, \I2.CHAINA_ERRS_net_1\, 
        \I2.un15_clear_stat_i\, \I2.CHAINB_ERRS_net_1\, 
        \I2.N_4180_i_0\, \I2.un1_DTO_cl_1_sqmuxa_2\, 
        \I2.N_4612_i_0\, \I2.N_4619_i_0\, \I2.N_4609_i_0\, 
        \I2.N_4626_i_0\, \I2.N_4615_i_0\, \I2.N_4623_i_0\, 
        \I2.N_4610_i_0\, \I2.N_4622_i_0\, \I2.N_4605_i_0\, 
        \I2.N_4621_i_0\, \I2.N_4613_i_0\, \I2.N_4624_i_0\, 
        \I2.STATE1_ns_il5r_net_1\, \I2.un3_hwres_i\, 
        \I2.STATE3_ns_il7r_net_1\, \I2.FIFO_FULL_net_1\, 
        \I2.SRAM_FULL_net_1\, \I2.CLK_sram\, \I2.WROi_net_1\, 
        \I2.WREi_net_1\, \I2.ERR_WORDS_RDY_net_1\, 
        \I2.STATE1l1r_net_1\, \I2.STATE4_ns_a3_il0r_net_1\, 
        \I2.TOKOUTBS_3_i_net_1\, \I2.TOKOUTAS_3_i_net_1\, 
        \I2.DTO_cl_64_il31r_net_1\, \I2.un1_DTO_cl_0_sqmuxa\, 
        \I2.STATEe_nsl2r\, \I2.STATEe_ns_il1r_net_1\, 
        \I2.STATEe_ns_i_0_il1r\, \I2.INT_ERRS_net_1\, 
        \I2.STATEe_nsl4r_net_1\, \I2.N_3510\, 
        \I2.STATEe_nsl3r_net_1\, \I2.STATEel4r_net_1\, 
        \I2.STATEe_nsl0r_net_1\, \I2.N_3453\, \I2.STATEe_ipl0r\, 
        \I2.N_3450\, \I2.STATEe_ipl1r\, \I2.STATEe_ipl2r\, 
        \I2.STATEe_ipl3r\, \I2.MSERCLKS_net_1\, 
        \I2.STATE5_ns_i_0l0r_net_1\, \I2.STATE5l0r_net_1\, 
        \I2.STATE5_ns_i_0_1_il0r\, \I2.N_4332\, \I2.STATE5_nsl3r\, 
        \I2.W_ERR_WORDS_net_1\, \I2.STATE4_ns_i_0l1r_net_1\, 
        \I2.N_4481\, \I2.N_4464\, \I2.L1AF3_i_0\, 
        \I2.STATE1_nsl7r\, \I2.STATE1_ns_1l7r\, 
        \I2.STATE1_ns_o2_0l0r_net_1\, \I2.N_3358\, 
        \I2.STATE1_ns_il14r_net_1\, \I2.END_CHAINB1_net_1\, 
        \I2.N_158\, \I2.STATE1_ns_il4r_net_1\, \I2.STATE1_nsl11r\, 
        \I2.un1_STATE1_27\, \I2.N_3889\, \I2.un1_STATE1_28\, 
        \I2.STATE1_1_sqmuxa_3\, \I2.STATE3l1r_net_1\, \I2.N_3015\, 
        \I2.N_3012\, \I2.STOP_RDSRAM_453_i_net_1\, \I2.N_145\, 
        \I2.STOP_RDSRAM_net_1\, \I2.STATE3_nsl12r_net_1\, 
        \I2.STATE3_nsl8r_net_1\, \I2.STATE3l5r_net_1\, 
        \I2.STATE3_il8r\, \I2.STATE3l6r_net_1\, 
        \I2.EVNT_NUM_963_net_1\, \I2.EVNT_NUM_n0_net_1\, 
        \I2.EVNT_NUMl0r_net_1\, \I2.N_3770\, \I2.N_1211\, 
        \I2.EVNT_NUM_962_net_1\, \I2.EVNT_NUM_n1_net_1\, 
        \I2.EVNT_NUMl1r_net_1\, \I2.N_1213\, 
        \I2.EVNT_NUM_961_net_1\, \I2.EVNT_NUM_n2_net_1\, 
        \I2.EVNT_NUMl2r_net_1\, \I2.EVNT_NUM_960_net_1\, 
        \I2.EVNT_NUM_n3_net_1\, \I2.EVNT_NUMl3r_net_1\, 
        \I2.EVNT_NUM_959_net_1\, \I2.EVNT_NUM_n4_net_1\, 
        \I2.EVNT_NUMl4r_net_1\, \I2.EVNT_NUM_958_net_1\, 
        \I2.EVNT_NUM_n5_net_1\, \I2.EVNT_NUMl5r_net_1\, 
        \I2.EVNT_NUM_957_net_1\, \I2.EVNT_NUM_n6_net_1\, 
        \I2.EVNT_NUMl6r_net_1\, \I2.EVNT_NUM_956_net_1\, 
        \I2.EVNT_NUM_n7_net_1\, \I2.EVNT_NUMl7r_net_1\, 
        \I2.EVNT_NUM_955_net_1\, \I2.EVNT_NUM_n8_net_1\, 
        \I2.EVNT_NUMl8r_net_1\, \I2.EVNT_NUM_954_net_1\, 
        \I2.EVNT_NUM_n9_net_1\, \I2.EVNT_NUMl9r_net_1\, 
        \I2.EVNT_NUM_953_net_1\, \I2.EVNT_NUM_n10_net_1\, 
        \I2.EVNT_NUMl10r_net_1\, \I2.EVNT_NUM_952_net_1\, 
        \I2.EVNT_NUM_n11_net_1\, \I2.EVNT_NUMl11r_net_1\, 
        \I2.N_1232\, \I2.N_1233\, \I2.FCNT_947_net_1\, 
        \I2.N_1236\, \I2.FCNT_c0\, \I2.N_3267\, 
        \I2.FCNT_946_net_1\, \I2.FCNT_n1_net_1\, 
        \I2.FCNTl1r_net_1\, \I2.N_1237\, \I2.un1_STATE1_22\, 
        \I2.FCNT_945_net_1\, \I2.FCNT_n2_i\, \I2.FCNTl2r_net_1\, 
        \I2.STATE1l13r_net_1\, \I2.FCNT_n2_tz_i\, \I2.FCNT_c1\, 
        \I2.L2ARR_944_net_1\, \I2.L2ARRl0r_net_1\, 
        \I2.L2ARR_943_net_1\, \I2.L2ARRl1r_net_1\, 
        \I2.L2ARR_942_net_1\, \I2.L2ARRl2r_net_1\, 
        \I2.L2ARR_941_net_1\, \I2.L2ARRl3r_net_1\, 
        \I2.G_EVNT_NUM_934_net_1\, \I2.G_EVNT_NUM_n0\, 
        \I2.N_3769\, \I2.G_EVNT_NUM_933_net_1\, \I2.N_4637\, 
        \I2.G_EVNT_NUMl1r_net_1\, \I2.G_EVNT_NUM_932_net_1\, 
        \I2.N_4342\, \I2.G_EVNT_NUMl2r_net_1\, 
        \I2.G_EVNT_NUM_931_net_1\, \I2.N_4343\, 
        \I2.G_EVNT_NUMl3r_net_1\, \I2.G_EVNT_NUM_930_net_1\, 
        \I2.N_4344\, \I2.G_EVNT_NUMl4r_net_1\, 
        \I2.G_EVNT_NUM_929_net_1\, \I2.N_4345\, 
        \I2.G_EVNT_NUMl5r_net_1\, \I2.G_EVNT_NUM_928_net_1\, 
        \I2.N_4638\, \I2.G_EVNT_NUMl6r_net_1\, 
        \I2.G_EVNT_NUM_927_net_1\, \I2.N_4639\, 
        \I2.G_EVNT_NUMl7r_net_1\, \I2.G_EVNT_NUM_926_net_1\, 
        \I2.N_4640\, \I2.G_EVNT_NUMl8r_net_1\, 
        \I2.G_EVNT_NUM_925_net_1\, \I2.G_EVNT_NUM_n9\, 
        \I2.G_EVNT_NUMl9r_net_1\, \I2.G_EVNT_NUM_924_net_1\, 
        \I2.G_EVNT_NUM_n10\, \I2.G_EVNT_NUMl10r_net_1\, 
        \I2.G_EVNT_NUM_n10_0_a2_0_0_i\, \I2.N_285_1\, 
        \I2.G_EVNT_NUM_923_net_1\, \I2.G_EVNT_NUM_n11\, 
        \I2.G_EVNT_NUMl11r_net_1\, \I2.N_287\, 
        \I2.L2SERV_922_net_1\, \I2.L2SERVe\, \I2.RPAGEl12r\, 
        \I2.L2SERV_921_net_1\, \I2.RPAGEl13r\, 
        \I2.L2SERV_920_net_1\, \I2.RPAGEl14r\, 
        \I2.EVNT_REJ_2_sqmuxa_net_1\, \I2.ROFFSET_918_net_1\, 
        \I2.ROFFSETl0r_net_1\, \I2.ROFFSET_n0_net_1\, \I2.N_1355\, 
        \I2.ROFFSET_917_net_1\, \I2.ROFFSETl1r_net_1\, 
        \I2.ROFFSET_n1_net_1\, \I2.N_1357\, 
        \I2.ROFFSET_916_net_1\, \I2.ROFFSETl2r_net_1\, 
        \I2.ROFFSET_n2_net_1\, \I2.ROFFSET_915_net_1\, 
        \I2.ROFFSETl3r_net_1\, \I2.ROFFSET_n3_net_1\, 
        \I2.ROFFSET_914_net_1\, \I2.ROFFSETl4r_net_1\, 
        \I2.ROFFSET_n4_net_1\, \I2.ROFFSET_913_net_1\, 
        \I2.ROFFSETl5r_net_1\, \I2.ROFFSET_n5_net_1\, 
        \I2.ROFFSET_912_net_1\, \I2.ROFFSETl6r_net_1\, 
        \I2.ROFFSET_n6_net_1\, \I2.ROFFSET_911_net_1\, 
        \I2.ROFFSETl7r_net_1\, \I2.ROFFSET_n7_net_1\, 
        \I2.ROFFSET_910_net_1\, \I2.ROFFSETl8r_net_1\, 
        \I2.ROFFSET_n8_net_1\, \I2.ROFFSET_909_net_1\, 
        \I2.ROFFSETl9r_net_1\, \I2.ROFFSET_n9_net_1\, 
        \I2.ROFFSET_908_net_1\, \I2.ROFFSETl10r_net_1\, 
        \I2.ROFFSET_n10_net_1\, \I2.ROFFSET_907_net_1\, 
        \I2.ROFFSETl11r_net_1\, \I2.ROFFSET_n11_net_1\, 
        \I2.ROFFSET_906_net_1\, \I2.ROFFSETl12r_net_1\, 
        \I2.ROFFSET_n12_net_1\, \I2.N_1378\, \I2.N_1379\, 
        \I2.DTO_16_1l31r\, \I2.DTO_9l31r\, \I2.DT_SRAMl31r_net_1\, 
        \I2.DT_TEMPl31r_net_1\, \I2.DTO_16_1_ivl30r_net_1\, 
        \I2.DT_SRAMl30r_net_1\, \I2.DTO_16_1_iv_1l30r_net_1\, 
        \I2.DTO_9_ivl30r_net_1\, \I2.DT_TEMPl30r_net_1\, 
        \I2.DTO_16_1l29r\, \I2.N_4159\, \I2.DT_SRAMl29r_net_1\, 
        \I2.DT_TEMPl29r_net_1\, \I2.DTO_16_1_ivl28r_net_1\, 
        \I2.DT_SRAM_i_m_0l28r_net_1\, 
        \I2.DTO_16_1_iv_0l28r_net_1\, \I2.DT_TEMPl28r_net_1\, 
        \I2.DT_SRAMl28r_net_1\, \I2.DT_TEMPl27r_net_1\, 
        \I2.N_4671\, \I2.N_457\, \I2.N_197\, \I2.N_4647\, 
        \I2.DT_TEMPl26r_net_1\, \I2.DT_SRAMl26r_net_1\, 
        \I2.DT_TEMPl25r_net_1\, \I2.DT_SRAMl25r_net_1\, 
        \I2.DTO_9l24r\, \I2.N_4194\, \I2.DT_TEMPl24r_net_1\, 
        \I2.DTO_9l23r\, \I2.DT_SRAMl23r_net_1\, 
        \I2.DT_TEMPl23r_net_1\, \I2.DTO_9l22r\, 
        \I2.DT_SRAMl22r_net_1\, \I2.DT_TEMPl22r_net_1\, 
        \I2.DT_TEMPl21r_net_1\, \I2.DT_SRAMl21r_net_1\, 
        \I2.DTO_9l20r\, \I2.DT_SRAMl20r_net_1\, 
        \I2.DT_TEMPl20r_net_1\, \I2.N_196\, 
        \I2.DT_TEMPl19r_net_1\, \I2.DT_SRAMl19r_net_1\, 
        \I2.N_202_i\, \I2.DTO_16_1_iv_0_a2_4_18_N_12_i\, 
        \I2.DTO_16_1_iv_0_a2_4_18_N_14_i\, 
        \I2.DTO_16_1_iv_0_a2_4_18_m7_0_0_i\, 
        \I2.DT_TEMPl18r_net_1\, \I2.ENDF_net_1\, 
        \I2.END_EVNT2_net_1\, \I2.DTO_16_1_iv_0_a2_4_18_N_11\, 
        \I2.END_EVNT5_net_1\, \I2.END_EVNT10_net_1\, 
        \I2.DT_TEMPl17r_net_1\, \I2.N_188\, 
        \I2.DT_TEMPl16r_net_1\, \I2.DT_SRAMl16r_net_1\, 
        \I2.DTO_9l15r\, \I2.DT_SRAMl15r_net_1\, 
        \I2.DT_TEMPl15r_net_1\, \I2.DTO_9l14r\, 
        \I2.DT_SRAMl14r_net_1\, \I2.DT_TEMPl14r_net_1\, 
        \I2.N_4048\, \I2.DT_TEMPl13r_net_1\, 
        \I2.DT_SRAMl12r_net_1\, \I2.N_3966\, 
        \I2.DT_TEMPl12r_net_1\, \I2.DTO_9l11r\, 
        \I2.DT_SRAMl11r_net_1\, \I2.DT_TEMPl11r_net_1\, 
        \I2.DT_TEMPl10r_net_1\, \I2.DT_SRAMl10r_net_1\, 
        \I2.DT_TEMPl9r_net_1\, \I2.N_4047\, \I2.N_223\, 
        \I2.DT_SRAMl8r_net_1\, \I2.N_3967\, \I2.DT_TEMPl8r_net_1\, 
        \I2.DTO_9l7r\, \I2.DT_SRAMl7r_net_1\, 
        \I2.DT_TEMPl7r_net_1\, \I2.DT_TEMPl6r_net_1\, 
        \I2.DT_SRAMl6r_net_1\, \I2.N_4030\, \I2.DTO_16_1l5r\, 
        \I2.DT_SRAMl5r_net_1\, \I2.DT_TEMPl5r_net_1\, 
        \I2.DTO_9l5r\, \I2.DT_TEMPl4r_net_1\, 
        \I2.DT_SRAMl4r_net_1\, \I2.DTO_16_1_ivl3r_net_1\, 
        \I2.DT_SRAMl3r_net_1\, \I2.DTO_16_1_iv_1l3r_net_1\, 
        \I2.DTO_9_ivl3r_net_1\, \I2.DT_TEMPl3r_net_1\, 
        \I2.DTO_16_1_ivl2r\, \I2.N_4193\, 
        \I2.DTO_16_1_iv_0_1l2r_net_1\, \I2.DTO_9_ivl2r\, 
        \I2.DT_TEMPl2r_net_1\, \I2.DTO_16_1_ivl1r_net_1\, 
        \I2.DT_SRAMl1r_net_1\, \I2.DTO_16_1_iv_1l1r_net_1\, 
        \I2.DTO_9_ivl1r_net_1\, \I2.DT_TEMPl1r_net_1\, 
        \I2.DTO_16_1_ivl0r\, \I2.DT_SRAMl0r_net_1\, 
        \I2.DTO_16_1_iv_0_0_1l0r_net_1\, \I2.DTO_9_ivl0r\, 
        \I2.DT_TEMPl0r_net_1\, \I2.STATE2l5r_net_1\, 
        \I2.PIPE2_DTl18r_net_1\, \I2.N_4038\, 
        \I2.DTO_cl_63_871_net_1\, \I2.N_2836\, 
        \I2.DTE_cl_63_870_net_1\, \I2.N_2822\, 
        \I2.DTE_1_869_net_1\, \I2.DTE_21_1l31r\, 
        \I2.DTE_1_868_net_1\, \I2.DTE_21_1_0_ivl30r_net_1\, 
        \I2.DTE_21_1_0_iv_1l30r_net_1\, 
        \I2.DT_SRAM_i_ml30r_net_1\, \I2.DTE_1_867_net_1\, 
        \I2.DTE_21_1l29r\, \I2.L_LUT_net_1\, \I2.CRC32l11r_net_1\, 
        \I2.CRC32l23r_net_1\, \I2.CRC32l10r_net_1\, 
        \I2.CRC32l22r_net_1\, \I2.CRC32l21r_net_1\, 
        \I2.CRC32l8r_net_1\, \I2.CRC32l20r_net_1\, 
        \I2.CRC32l31r_net_1\, \I2.CRC32l19r_net_1\, 
        \I2.CRC32l7r_net_1\, \I2.CRC32l30r_net_1\, 
        \I2.CRC32l18r_net_1\, \I2.CRC32l6r_net_1\, 
        \I2.CRC32l29r_net_1\, \I2.CRC32l17r_net_1\, 
        \I2.CRC32l5r_net_1\, \I2.CRC32l28r_net_1\, 
        \I2.CRC32l16r_net_1\, \I2.CRC32l4r_net_1\, 
        \I2.CRC32l27r_net_1\, \I2.CRC32l15r_net_1\, 
        \I2.CRC32l26r_net_1\, \I2.CRC32l14r_net_1\, 
        \I2.CRC32l2r_net_1\, \I2.DTE_1_845_net_1\, 
        \I2.DTE_21_1l5r\, \I2.N_4266\, \I2.DT_TEMP_7l5r_net_1\, 
        \I2.CRC32l25r_net_1\, \I2.CRC32l13r_net_1\, 
        \I2.CRC32l24r_net_1\, \I2.CRC32l12r_net_1\, 
        \I2.CRC32l0r_net_1\, \I2.DTE_1_843_net_1\, 
        \I2.DTE_21_1_iv_i_0l3r\, \I2.DTE_21_1_iv_2_il3r\, 
        \I2.DTE_1_842_net_1\, \I2.DTE_21_1_iv_i_0l2r\, 
        \I2.DTE_21_1_iv_2_il2r\, \I2.DTE_1_841_net_1\, 
        \I2.DTE_21_1_iv_i_0l1r\, \I2.DTE_21_1_iv_2_il1r\, 
        \I2.DTE_1_840_net_1\, \I2.DTE_21_1_iv_i_0l0r\, 
        \I2.DTE_21_1_iv_2_il0r\, 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_N_20_i\, 
        \I2.NWPIPE10_net_1\, \I2.I_73\, \I2.N_4262\, \I2.I_66\, 
        \I2.I_56\, \I2.I_52\, \I2.I_45\, \I2.I_38\, \I2.I_31\, 
        \I2.I_24\, \I2.I_20\, \I2.I_13_1\, \I2.I_9_0\, \I2.I_5_0\, 
        \I2.WOFFSET_13l0r\, \I2.CRC32_826_net_1\, \I2.N_3948\, 
        \I2.N_244_i_i_0\, \I2.N_232_i_i\, \I2.CRC32_825_net_1\, 
        \I2.N_3947\, \I2.N_245_i_i_0\, \I2.N_231_i_i\, 
        \I2.CRC32_824_net_1\, \I2.N_3946\, \I2.N_18_i_0_i_0\, 
        \I2.N_4157_i_i\, \I2.CRC32_823_net_1\, \I2.N_3945\, 
        \I2.N_19_i_0_i_0\, \I2.N_4156_i_i\, \I2.CRC32_822_net_1\, 
        \I2.N_3944\, \I2.N_246_i_i_0\, \I2.N_230_i_i\, 
        \I2.CRC32_821_net_1\, \I2.N_3943\, \I2.N_127_i_0_i_0\, 
        \I2.N_4271_i_i\, \I2.CRC32_820_net_1\, \I2.N_3942\, 
        \I2.N_42_i_0_i_0\, \I2.N_4349_i_i\, \I2.CRC32_819_net_1\, 
        \I2.N_3941\, \I2.N_128_i_0_i_0\, \I2.N_4270_i_i\, 
        \I2.CRC32_818_net_1\, \I2.N_3940\, \I2.N_129_i_0_i_0\, 
        \I2.N_4269_i_i\, \I2.CRC32_817_net_1\, \I2.N_3939\, 
        \I2.N_130_i_0_i_0\, \I2.N_4268_i_i\, \I2.CRC32_816_net_1\, 
        \I2.N_3938\, \I2.N_58_i_0_i_0\, \I2.N_4039_i_i\, 
        \I2.CRC32_815_net_1\, \I2.N_3937\, \I2.N_111_i_i_0\, 
        \I2.N_3962_i_i\, \I2.CRC32_814_net_1\, \I2.N_3936\, 
        \I2.N_247_i_i_0\, \I2.N_229_i_i\, \I2.CRC32_813_net_1\, 
        \I2.N_3935\, \I2.N_52_i_0_i_0\, \I2.N_4096_i_i\, 
        \I2.CRC32_812_net_1\, \I2.N_3934\, \I2.N_252_i_i_0\, 
        \I2.N_224_i_i\, \I2.CRC32_811_net_1\, \I2.N_3933\, 
        \I2.N_112_i_i_0\, \I2.N_3961_i_i\, \I2.CRC32_810_net_1\, 
        \I2.N_3932\, \I2.N_113_i_i_0\, \I2.N_3960_i_i\, 
        \I2.CRC32_809_net_1\, \I2.N_3931\, \I2.N_4026_i_0\, 
        \I2.N_3959_i_i\, \I2.CRC32_808_net_1\, \I2.N_3930\, 
        \I2.N_115_i_i_0\, \I2.N_3958_i_i\, \I2.CRC32_807_net_1\, 
        \I2.N_3929\, \I2.N_116_i_i_0\, \I2.N_3957_i_i\, 
        \I2.CRC32_806_net_1\, \I2.N_3928\, \I2.N_248_i_i_0\, 
        \I2.N_228_i_i\, \I2.CRC32_805_net_1\, \I2.N_3927\, 
        \I2.N_249_i_i_0\, \I2.N_227_i_i\, \I2.CRC32l9r_net_1\, 
        \I2.N_3926\, \I2.N_56_i_0\, \I2.CRC32_803_net_1\, 
        \I2.N_3925\, \I2.N_117_i_i_0\, \I2.N_3956_i_i\, 
        \I2.CRC32_802_net_1\, \I2.N_3924\, \I2.N_250_i_i_0\, 
        \I2.N_226_i_i\, \I2.CRC32_801_net_1\, \I2.N_3923\, 
        \I2.N_251_i_i_0\, \I2.N_225_i_i\, \I2.CRC32_800_net_1\, 
        \I2.N_3922\, \I2.N_131_i_0_i_0\, \I2.N_4267_i_i\, 
        \I2.CRC32_799_net_1\, \I2.N_3921\, \I2.N_118_i_i_0\, 
        \I2.N_3955_i_i\, \I2.CRC32l3r_net_1\, \I2.N_3920\, 
        \I2.CRC32_2l3r_net_1\, \I2.CRC32_797_net_1\, \I2.N_3919\, 
        \I2.N_73_i_0_i_0\, \I2.N_4187_i_i\, \I2.CRC32l1r_net_1\, 
        \I2.N_3918\, \I2.N_999\, \I2.CRC32_2_il1r\, 
        \I2.CRC32_795_net_1\, \I2.N_3917\, \I2.N_4184\, 
        \I2.N_4027_i_0\, \I2.N_3954_i_i\, \I2.WREi_794_net_1\, 
        \I2.N_4203\, \I2.WREi_8_i_i_a2_1_net_1\, 
        \I2.WROi_793_net_1\, \I2.WROi_10\, \I2.DT_TEMP_792_net_1\, 
        \I2.DT_TEMP_7l31r_net_1\, \I2.PIPE2_DTl31r_net_1\, 
        \I2.N_899\, \I2.PIPE5_DTl31r_net_1\, 
        \I2.PIPE10_DTl31r_net_1\, \I2.DT_TEMP_791_net_1\, 
        \I2.DT_TEMP_7l30r_net_1\, \I2.PIPE2_DTl30r_net_1\, 
        \I2.N_898\, \I2.PIPE5_DTl30r_net_1\, 
        \I2.PIPE10_DTl30r_net_1\, \I2.DT_TEMP_790_net_1\, 
        \I2.DT_TEMP_7l29r_net_1\, \I2.PIPE2_DTl29r_net_1\, 
        \I2.N_897\, \I2.PIPE5_DTl29r_net_1\, 
        \I2.PIPE10_DTl29r_net_1\, \I2.DT_TEMP_789_net_1\, 
        \I2.DT_TEMP_7l28r_net_1\, \I2.PIPE2_DTl28r_net_1\, 
        \I2.N_896\, \I2.PIPE5_DTl28r_net_1\, 
        \I2.PIPE10_DTl28r_net_1\, \I2.DT_TEMP_788_net_1\, 
        \I2.DT_TEMP_7l27r_net_1\, \I2.PIPE2_DTl27r_net_1\, 
        \I2.DT_SRAM_0_il27r_net_1\, \I2.PIPE10_DTl27r_net_1\, 
        \I2.PIPE5_DTl27r_net_1\, \I2.DT_TEMP_787_net_1\, 
        \I2.DT_TEMP_7l26r_net_1\, \I2.PIPE2_DTl26r_net_1\, 
        \I2.N_894\, \I2.PIPE5_DTl26r_net_1\, 
        \I2.PIPE10_DTl26r_net_1\, \I2.DT_TEMP_786_net_1\, 
        \I2.DT_TEMP_7l25r_net_1\, \I2.PIPE2_DTl25r_net_1\, 
        \I2.N_893\, \I2.PIPE5_DTl25r_net_1\, 
        \I2.PIPE10_DTl25r_net_1\, \I2.DT_TEMP_785_net_1\, 
        \I2.DT_TEMP_7l24r_net_1\, \I2.PIPE2_DTl24r_net_1\, 
        \I2.N_4192\, \I2.PIPE5_DTl24r_net_1\, 
        \I2.PIPE10_DTl24r_net_1\, \I2.DT_TEMP_784_net_1\, 
        \I2.DT_TEMP_7l23r_net_1\, \I2.PIPE2_DTl23r_net_1\, 
        \I2.N_891\, \I2.PIPE5_DTl23r_net_1\, 
        \I2.PIPE10_DTl23r_net_1\, \I2.DT_TEMP_783_net_1\, 
        \I2.DT_TEMP_7l22r_net_1\, \I2.PIPE2_DTl22r_net_1\, 
        \I2.N_890\, \I2.PIPE10_DTl22r_net_1\, 
        \I2.DT_TEMP_782_net_1\, \I2.DT_TEMP_7l21r_net_1\, 
        \I2.PIPE2_DTl21r_net_1\, \I2.N_889\, 
        \I2.PIPE5_DTl21r_net_1\, \I2.PIPE10_DTl21r_net_1\, 
        \I2.DT_TEMP_781_net_1\, \I2.DT_TEMP_7l20r_net_1\, 
        \I2.PIPE2_DTl20r_net_1\, \I2.N_888\, 
        \I2.PIPE5_DTl20r_net_1\, \I2.PIPE10_DTl20r_net_1\, 
        \I2.DT_TEMP_780_net_1\, \I2.DT_TEMP_7l19r_net_1\, 
        \I2.PIPE2_DTl19r_net_1\, \I2.N_887\, 
        \I2.PIPE5_DTl19r_net_1\, \I2.PIPE10_DTl19r_net_1\, 
        \I2.DT_TEMP_779_net_1\, \I2.DT_TEMP_7l18r_net_1\, 
        \I2.PIPE5_DTl18r_net_1\, \I2.PIPE10_DTl18r_net_1\, 
        \I2.DT_TEMP_778_net_1\, \I2.DT_TEMP_7l17r_net_1\, 
        \I2.PIPE2_DTl17r_net_1\, \I2.N_4645\, 
        \I2.PIPE5_DTl17r_net_1\, \I2.PIPE10_DTl17r_net_1\, 
        \I2.DT_TEMP_777_net_1\, \I2.DT_TEMP_7l16r_net_1\, 
        \I2.PIPE2_DTl16r_net_1\, \I2.N_884\, 
        \I2.PIPE5_DTl16r_net_1\, \I2.PIPE10_DTl16r_net_1\, 
        \I2.DT_TEMP_776_net_1\, \I2.DT_TEMP_7l15r_net_1\, 
        \I2.PIPE2_DTl15r_net_1\, \I2.N_883\, 
        \I2.PIPE5_DTl15r_net_1\, \I2.PIPE10_DTl15r_net_1\, 
        \I2.DT_TEMP_775_net_1\, \I2.DT_TEMP_7l14r_net_1\, 
        \I2.PIPE2_DTl14r_net_1\, \I2.N_882\, 
        \I2.PIPE5_DTl14r_net_1\, \I2.PIPE10_DTl14r_net_1\, 
        \I2.DT_TEMP_774_net_1\, \I2.DT_TEMP_7l13r_net_1\, 
        \I2.PIPE2_DTl13r_net_1\, \I2.N_4046\, 
        \I2.PIPE5_DTl13r_net_1\, \I2.PIPE10_DTl13r_net_1\, 
        \I2.DT_TEMP_773_net_1\, \I2.DT_TEMP_7l12r_net_1\, 
        \I2.PIPE2_DTl12r_net_1\, \I2.N_880\, 
        \I2.PIPE5_DTl12r_net_1\, \I2.PIPE10_DTl12r_net_1\, 
        \I2.DT_TEMP_772_net_1\, \I2.DT_TEMP_7l11r_net_1\, 
        \I2.PIPE2_DTl11r_net_1\, \I2.N_879\, 
        \I2.PIPE5_DTl11r_net_1\, \I2.PIPE10_DTl11r_net_1\, 
        \I2.DT_TEMP_771_net_1\, \I2.DT_TEMP_7l10r_net_1\, 
        \I2.PIPE2_DTl10r_net_1\, \I2.N_878\, 
        \I2.PIPE5_DTl10r_net_1\, \I2.PIPE10_DTl10r_net_1\, 
        \I2.DT_TEMP_770_net_1\, \I2.DT_TEMP_7l9r_net_1\, 
        \I2.PIPE2_DTl9r_net_1\, \I2.N_4045\, 
        \I2.PIPE5_DTl9r_net_1\, \I2.PIPE10_DTl9r_net_1\, 
        \I2.DT_TEMP_769_net_1\, \I2.DT_TEMP_7l8r_net_1\, 
        \I2.PIPE2_DTl8r_net_1\, \I2.N_876\, 
        \I2.PIPE5_DTl8r_net_1\, \I2.PIPE10_DTl8r_net_1\, 
        \I2.DT_TEMP_768_net_1\, \I2.DT_TEMP_7l7r_net_1\, 
        \I2.PIPE2_DTl7r_net_1\, \I2.N_875\, 
        \I2.PIPE5_DTl7r_net_1\, \I2.PIPE10_DTl7r_net_1\, 
        \I2.DT_TEMP_767_net_1\, \I2.DT_TEMP_7l6r_net_1\, 
        \I2.PIPE2_DTl6r_net_1\, \I2.N_874\, 
        \I2.PIPE5_DTl6r_net_1\, \I2.PIPE10_DTl6r_net_1\, 
        \I2.DT_TEMP_766_net_1\, \I2.PIPE2_DTl5r_net_1\, 
        \I2.N_873\, \I2.PIPE5_DTl5r_net_1\, 
        \I2.PIPE10_DTl5r_net_1\, \I2.DT_TEMP_765_net_1\, 
        \I2.DT_TEMP_7l4r_net_1\, \I2.PIPE2_DTl4r_net_1\, 
        \I2.N_872\, \I2.PIPE5_DTl4r_net_1\, 
        \I2.PIPE10_DTl4r_net_1\, \I2.DT_TEMP_764_net_1\, 
        \I2.DT_TEMP_7l3r_net_1\, \I2.PIPE2_DTl3r_net_1\, 
        \I2.N_871\, \I2.PIPE5_DTl3r_net_1\, 
        \I2.PIPE10_DTl3r_net_1\, \I2.DT_TEMP_763_net_1\, 
        \I2.DT_TEMP_7l2r_net_1\, \I2.PIPE2_DTl2r_net_1\, 
        \I2.N_4191\, \I2.PIPE5_DTl2r_net_1\, 
        \I2.PIPE10_DTl2r_net_1\, \I2.DT_TEMP_762_net_1\, 
        \I2.DT_TEMP_7l1r_net_1\, \I2.PIPE2_DTl1r_net_1\, 
        \I2.N_869\, \I2.PIPE5_DTl1r_net_1\, 
        \I2.PIPE10_DTl1r_net_1\, \I2.DT_TEMP_761_net_1\, 
        \I2.DT_TEMP_7l0r_net_1\, \I2.PIPE2_DTl0r_net_1\, 
        \I2.N_868\, \I2.PIPE5_DTl0r_net_1\, 
        \I2.PIPE10_DTl0r_net_1\, \I2.TEMPF_760_net_1\, 
        \I2.N_2849\, \I2.INC_EVNT_NUM_net_1\, 
        \I2.PIPE1_DT_758_net_1\, \I2.PIPE1_DT_42l31r\, 
        \I2.PIPE1_DTl31r_net_1\, \I2.PIPE1_DT_757_net_1\, 
        \I2.PIPE1_DT_42l30r\, \I2.PIPE1_DTl30r_net_1\, 
        \I2.TDCDASl28r_net_1\, \I2.TDCDBSl28r_net_1\, 
        \I2.PIPE1_DT_756_net_1\, \I2.PIPE1_DT_42l29r\, 
        \I2.PIPE1_DTl29r_net_1\, \I2.N_3254\, 
        \I2.PIPE1_DT_755_net_1\, \I2.PIPE1_DT_42l28r\, 
        \I2.PIPE1_DTl28r_net_1\, \I2.PIPE1_DT_754_net_1\, 
        \I2.PIPE1_DT_42_1_iv_i_0l27r\, \I2.PIPE1_DTl27r_net_1\, 
        \I2.PIPE1_DT_42_1_iv_2_il27r\, \I2.TDCDBSl27r_net_1\, 
        \I2.TDCDASl27r_net_1\, \I2.PIPE1_DT_753_net_1\, 
        \I2.PIPE1_DT_42_1_iv_i_0l26r\, \I2.PIPE1_DTl26r_net_1\, 
        \I2.PIPE1_DT_42_1_iv_2_il26r\, \I2.TDCDBSl26r_net_1\, 
        \I2.TDCDASl26r_net_1\, \I2.PIPE1_DT_752_net_1\, 
        \I2.PIPE1_DT_42_1_iv_i_0l25r\, \I2.PIPE1_DTl25r_net_1\, 
        \I2.PIPE1_DT_42_1_iv_2l25r_net_1\, \I2.TDCDBSl25r_net_1\, 
        \I2.PIPE1_DT_42_1_iv_1_il25r\, \I2.TDCDASl25r_net_1\, 
        \I2.STATE1l18r_net_1\, \I2.PIPE1_DT_751_net_1\, 
        \I2.PIPE1_DT_42_1_iv_i_0l24r\, \I2.PIPE1_DTl24r_net_1\, 
        \I2.EVNT_NUM_i_m_il8r\, \I2.PIPE1_DT_42_1_iv_1_il24r\, 
        \I2.PIPE1_DT_42_1_iv_0_il24r\, \I2.TDCDASl24r_net_1\, 
        \I2.TDCDBSl24r_net_1\, \I2.PIPE1_DT_750_net_1\, 
        \I2.PIPE1_DT_42l23r\, \I2.PIPE1_DTl23r_net_1\, 
        \I2.TDCDASl23r_net_1\, \I2.TDCDBSl23r_net_1\, 
        \I2.PIPE1_DT_749_net_1\, \I2.PIPE1_DT_42l22r\, 
        \I2.PIPE1_DTl22r_net_1\, \I2.TDCDASl22r_net_1\, 
        \I2.TDCDBSl22r_net_1\, \I2.PIPE1_DT_748_net_1\, 
        \I2.PIPE1_DT_42l21r\, \I2.PIPE1_DTl21r_net_1\, 
        \I2.TDCDASl21r_net_1\, \I2.TDCDBSl21r_net_1\, 
        \I2.PIPE1_DT_747_net_1\, \I2.PIPE1_DT_42l20r\, 
        \I2.PIPE1_DTl20r_net_1\, \I2.TDCDASl20r_net_1\, 
        \I2.TDCDBSl20r_net_1\, \I2.PIPE1_DT_746_net_1\, 
        \I2.PIPE1_DT_42l19r\, \I2.PIPE1_DTl19r_net_1\, 
        \I2.TDCDASl19r_net_1\, \I2.TDCDBSl19r_net_1\, 
        \I2.PIPE1_DT_745_net_1\, \I2.PIPE1_DT_42l18r\, 
        \I2.PIPE1_DTl18r_net_1\, \I2.PIPE1_DT_744_net_1\, 
        \I2.PIPE1_DT_42l17r\, \I2.PIPE1_DTl17r_net_1\, 
        \I2.PIPE1_DT_743_net_1\, \I2.PIPE1_DT_42l16r\, 
        \I2.PIPE1_DTl16r_net_1\, \I2.STATE1l11r_net_1\, 
        \I2.PIPE1_DT_1_sqmuxa\, \I2.TOKOUTAS_net_1\, 
        \I2.TOKOUTBS_net_1\, \I2.N_3902\, 
        \I2.MIC_ERR_REGSl48r_net_1\, \I2.PIPE1_DT_742_net_1\, 
        \I2.PIPE1_DT_42l15r\, \I2.PIPE1_DTl15r_net_1\, 
        \I2.MIC_ERR_REGSl15r_net_1\, \I2.MIC_ERR_REGSl31r_net_1\, 
        \I2.MIC_ERR_REGSl47r_net_1\, \I2.BNCID_VECTrxl11r\, 
        \I2.BNCID_VECTror_net_1\, \I2.N_3238\, \I2.DOUT_TMPl3r\, 
        \I2.DIN_REG1l3r\, \I2.N_13\, \I2.PIPE1_DT_741_net_1\, 
        \I2.PIPE1_DT_42l14r\, \I2.PIPE1_DTl14r_net_1\, 
        \I2.MIC_ERR_REGSl14r_net_1\, \I2.MIC_ERR_REGSl30r_net_1\, 
        \I2.MIC_ERR_REGSl46r_net_1\, \I2.BNCID_VECTrxl10r\, 
        \I2.DOUT_TMPl2r\, \I2.DIN_REG1l2r\, 
        \I2.PIPE1_DT_740_net_1\, \I2.PIPE1_DT_42l13r\, 
        \I2.PIPE1_DTl13r_net_1\, \I2.MIC_ERR_REGSl13r_net_1\, 
        \I2.MIC_ERR_REGSl29r_net_1\, \I2.MIC_ERR_REGSl45r_net_1\, 
        \I2.BNCID_VECTrxl9r\, \I2.DOUT_TMPl1r\, \I2.DIN_REG1l1r\, 
        \I2.PIPE1_DT_739_net_1\, \I2.PIPE1_DT_42l12r\, 
        \I2.PIPE1_DTl12r_net_1\, \I2.MIC_ERR_REGSl12r_net_1\, 
        \I2.MIC_ERR_REGSl28r_net_1\, \I2.MIC_ERR_REGSl44r_net_1\, 
        \I2.BNCID_VECTrxl8r\, \I2.DOUT_TMPl0r\, \I2.DIN_REG1l0r\, 
        \I2.PIPE1_DT_738_net_1\, \I2.PIPE1_DT_42l11r\, 
        \I2.PIPE1_DTl11r_net_1\, \I2.MIC_ERR_REGSl11r_net_1\, 
        \I2.MIC_ERR_REGSl27r_net_1\, \I2.MIC_ERR_REGSl43r_net_1\, 
        \I2.BNCID_VECTrxl7r\, \I2.DOUT_TMPl7r\, \I2.DIN_REG1l7r\, 
        \I2.PIPE1_DT_737_net_1\, \I2.PIPE1_DT_42l10r\, 
        \I2.PIPE1_DTl10r_net_1\, \I2.MIC_ERR_REGSl10r_net_1\, 
        \I2.MIC_ERR_REGSl26r_net_1\, \I2.MIC_ERR_REGSl42r_net_1\, 
        \I2.BNCID_VECTrxl6r\, \I2.DOUT_TMPl6r\, \I2.DIN_REG1l6r\, 
        \I2.PIPE1_DT_736_net_1\, \I2.PIPE1_DT_42l9r\, 
        \I2.PIPE1_DTl9r_net_1\, \I2.TDCDBSl7r_net_1\, 
        \I2.MIC_ERR_REGSl9r_net_1\, \I2.MIC_ERR_REGSl25r_net_1\, 
        \I2.MIC_ERR_REGSl41r_net_1\, \I2.TDCDASl7r_net_1\, 
        \I2.BNCID_VECTrxl5r\, \I2.DOUT_TMPl5r\, \I2.DIN_REG1l5r\, 
        \I2.PIPE1_DT_735_net_1\, \I2.PIPE1_DT_42l8r\, 
        \I2.PIPE1_DTl8r_net_1\, \I2.TDCDBSl6r_net_1\, 
        \I2.MIC_ERR_REGSl8r_net_1\, \I2.MIC_ERR_REGSl24r_net_1\, 
        \I2.MIC_ERR_REGSl40r_net_1\, \I2.TDCDASl6r_net_1\, 
        \I2.BNCID_VECTrxl4r\, \I2.DOUT_TMPl4r\, \I2.DIN_REG1l4r\, 
        \I2.PIPE1_DT_734_net_1\, \I2.PIPE1_DT_42l7r\, 
        \I2.PIPE1_DTl7r_net_1\, \I2.TDCDBSl5r_net_1\, 
        \I2.MIC_ERR_REGSl7r_net_1\, \I2.MIC_ERR_REGSl23r_net_1\, 
        \I2.MIC_ERR_REGSl39r_net_1\, \I2.TDCDASl5r_net_1\, 
        \I2.BNCID_VECTrxl3r\, \I2.DOUT_TMP_0l3r\, 
        \I2.DIN_REG1_0l3r\, \I2.PIPE1_DT_733_net_1\, 
        \I2.PIPE1_DT_42l6r\, \I2.PIPE1_DTl6r_net_1\, 
        \I2.TDCDBSl4r_net_1\, \I2.MIC_ERR_REGSl6r_net_1\, 
        \I2.MIC_ERR_REGSl22r_net_1\, \I2.STATE1l3r_net_1\, 
        \I2.MIC_ERR_REGSl38r_net_1\, \I2.STATE1l0r_net_1\, 
        \I2.TDCDASl4r_net_1\, \I2.BNCID_VECTrxl2r\, 
        \I2.DOUT_TMP_0l2r\, \I2.DIN_REG1_0l2r\, 
        \I2.PIPE1_DT_732_net_1\, \I2.PIPE1_DT_42l5r\, 
        \I2.PIPE1_DTl5r_net_1\, \I2.TDCDBSl3r_net_1\, 
        \I2.MIC_ERR_REGSl5r_net_1\, \I2.MIC_ERR_REGSl21r_net_1\, 
        \I2.MIC_ERR_REGSl37r_net_1\, \I2.TDCDASl3r_net_1\, 
        \I2.BNCID_VECTrxl1r\, \I2.DOUT_TMP_0l1r\, 
        \I2.DIN_REG1_0l1r\, \I2.PIPE1_DT_731_net_1\, 
        \I2.PIPE1_DT_42l4r\, \I2.PIPE1_DTl4r_net_1\, 
        \I2.TDCDBSl2r_net_1\, \I2.MIC_ERR_REGSl4r_net_1\, 
        \I2.MIC_ERR_REGSl20r_net_1\, \I2.MIC_ERR_REGSl36r_net_1\, 
        \I2.TDCDASl2r_net_1\, \I2.BNCID_VECTrxl0r\, 
        \I2.DOUT_TMP_0l0r\, \I2.DIN_REG1_0l0r\, \I2.I_6_0_i_0_i\, 
        \I2.I_6_2_i_0_i\, \I2.WADDR_REG1l2r\, \I2.WADDR_REG1l0r\, 
        \I2.I_6_1_i_0_i\, \I2.I_6_3_i_0_i\, \I2.N_11\, 
        \I2.WADDR_REG1l3r\, \I2.TRGSERVl3r_net_1\, 
        \I2.WADDR_REG1l1r\, \I2.BNCID_VECTror_10_tz_0_net_1\, 
        \I2.BNCID_VECTria_7_0_net_1\, \I2.BNCID_VECTro_6\, 
        \I2.BNCID_VECTro_7\, \I2.BNCID_VECTro_4\, 
        \I2.BNCID_VECTro_5\, \I2.BNCID_VECTro_0\, 
        \I2.BNCID_VECTro_1\, \I2.BNCID_VECTro_3\, 
        \I2.BNCID_VECTro_2\, \I2.BNCID_VECTror_8_tz_0_i\, 
        \I2.BNCID_VECTria_11_0_i\, \I2.BNCID_VECTro_10\, 
        \I2.BNCID_VECTro_11\, \I2.BNCID_VECTro_8\, 
        \I2.BNCID_VECTro_9\, \I2.BNCID_VECTro_14\, 
        \I2.BNCID_VECTro_15\, \I2.BNCID_VECTro_12\, 
        \I2.BNCID_VECTro_13\, \I2.PIPE1_DT_730_net_1\, 
        \I2.PIPE1_DT_42l3r\, \I2.PIPE1_DTl3r_net_1\, 
        \I2.TDCDASl1r_net_1\, \I2.TDCDBSl1r_net_1\, 
        \I2.MIC_ERR_REGSl3r_net_1\, \I2.MIC_ERR_REGSl19r_net_1\, 
        \I2.MIC_ERR_REGSl35r_net_1\, \I2.PIPE1_DT_729_net_1\, 
        \I2.PIPE1_DT_42l2r\, \I2.PIPE1_DTl2r_net_1\, 
        \I2.TDCDASl0r_net_1\, \I2.TDCDBSl0r_net_1\, 
        \I2.MIC_ERR_REGSl2r_net_1\, \I2.MIC_ERR_REGSl18r_net_1\, 
        \I2.MIC_ERR_REGSl34r_net_1\, \I2.PIPE1_DT_728_net_1\, 
        \I2.PIPE1_DT_42l1r\, \I2.PIPE1_DTl1r_net_1\, 
        \I2.MIC_ERR_REGSl1r_net_1\, \I2.MIC_ERR_REGSl17r_net_1\, 
        \I2.MIC_ERR_REGSl33r_net_1\, \I2.N_148\, \I2.N_3891\, 
        \I2.PIPE1_DT_727_net_1\, \I2.PIPE1_DT_42l0r\, 
        \I2.PIPE1_DTl0r_net_1\, \I2.N_3885\, \I2.N_3898_i\, 
        \I2.STATE1_i_0_il15r\, \I2.STATE1_i_0_il16r\, 
        \I2.STATE1l6r_net_1\, \I2.MIC_ERR_REGSl0r_net_1\, 
        \I2.STATE1l9r_net_1\, \I2.MIC_ERR_REGSl16r_net_1\, 
        \I2.MIC_ERR_REGSl32r_net_1\, \I2.NWPIPE1_726_net_1\, 
        \I2.NWPIPE1_net_1\, \I2.un1_STATE1_39_i_0\, 
        \I2.un1_STATE1_38\, \I2.N_3292\, \I2.un1_STATE1_39_6_i\, 
        \I2.un5_tdcgda1_net_1\, \I2.EVNT_WORDl12r_net_1\, 
        \I2.EVNT_WORDl11r_net_1\, \I2.EVNT_WORDl10r_net_1\, 
        \I2.EVNT_WORDl9r_net_1\, \I2.EVNT_WORDl8r_net_1\, 
        \I2.EVNT_WORDl7r_net_1\, \I2.EVNT_WORDl6r_net_1\, 
        \I2.EVNT_WORDl5r_net_1\, \I2.EVNT_WORDl4r_net_1\, 
        \I2.EVNT_WORDl3r_net_1\, \I2.EVNT_WORDl2r_net_1\, 
        \I2.EVNT_WORDl1r_net_1\, \I2.EVNT_WORDl0r_net_1\, 
        \I2.ENDF_712_net_1\, \I2.un1_STATE2_9\, \I2.un1_STATE2_7\, 
        \I2.END_TDC1_711_net_1\, \I2.END_TDC1_net_1\, \I2.N_3281\, 
        \I2.STATE1l7r_net_1\, \I2.N_3273\, \I2.N_3344_i\, 
        \I2.END_EVNT1_710_net_1\, \I2.END_EVNT1_net_1\, 
        \I2.END_CHAINB1_709_net_1\, \I2.N_3883\, 
        \I2.END_CHAINA1_708_net_1\, \I2.PIPE5_DT_707_net_1\, 
        \I2.PIPE5_DT_706_net_1\, \I2.PIPE5_DT_705_net_1\, 
        \I2.PIPE4_DTl29r_net_1\, \I2.PIPE5_DT_704_net_1\, 
        \I2.PIPE5_DT_6l28r\, \I2.PIPE4_DTl28r_net_1\, 
        \I2.PIPE5_DT_703_net_1\, \I2.PIPE4_DTl27r_net_1\, 
        \I2.PIPE5_DT_702_net_1\, \I2.PIPE4_DTl26r_net_1\, 
        \I2.PIPE5_DT_701_net_1\, \I2.PIPE4_DTl25r_net_1\, 
        \I2.PIPE5_DT_700_net_1\, \I2.PIPE4_DTl24r_net_1\, 
        \I2.PIPE5_DT_699_net_1\, \I2.PIPE5_DT_697_net_1\, 
        \I2.PIPE5_DT_696_net_1\, \I2.PIPE5_DT_6l20r_net_1\, 
        \I2.PIPE5_DT_6_dl20r_net_1\, \I2.PIPE5_DT_6_sl19r_net_1\, 
        \I2.PIPE4_DTl20r_net_1\, \I2.PIPE4_DTl19r_net_1\, 
        \I2.PIPE5_DT_695_net_1\, \I2.PIPE5_DT_6l19r_net_1\, 
        \I2.PIPE5_DT_6_dl19r_net_1\, \I2.PIPE4_DTl18r_net_1\, 
        \I2.PIPE5_DT_694_net_1\, \I2.PIPE5_DT_6l18r_net_1\, 
        \I2.PIPE5_DT_6_dl18r_net_1\, \I2.PIPE4_DTl17r_net_1\, 
        \I2.PIPE5_DT_693_net_1\, \I2.PIPE5_DT_6l17r_net_1\, 
        \I2.PIPE5_DT_6_dl17r_net_1\, \I2.PIPE4_DTl16r_net_1\, 
        \I2.PIPE5_DT_692_net_1\, \I2.PIPE5_DT_6l16r_net_1\, 
        \I2.PIPE4_DTl15r_net_1\, \I2.PIPE5_DT_691_net_1\, 
        \I2.PIPE5_DT_6l15r_net_1\, \I2.PIPE4_DTl14r_net_1\, 
        \I2.PIPE5_DT_690_net_1\, \I2.PIPE5_DT_6l14r_net_1\, 
        \I2.PIPE4_DTl13r_net_1\, \I2.PIPE5_DT_689_net_1\, 
        \I2.PIPE5_DT_6l13r_net_1\, \I2.PIPE4_DTl12r_net_1\, 
        \I2.PIPE5_DT_688_net_1\, \I2.PIPE5_DT_6l12r_net_1\, 
        \I2.PIPE4_DTl11r_net_1\, \I2.PIPE5_DT_687_net_1\, 
        \I2.PIPE5_DT_6l11r_net_1\, \I2.PIPE5_DT_686_net_1\, 
        \I2.PIPE5_DT_6l10r_net_1\, \I2.PIPE5_DT_685_net_1\, 
        \I2.PIPE5_DT_6l9r_net_1\, \I2.PIPE5_DT_684_net_1\, 
        \I2.PIPE5_DT_6l8r_net_1\, \I2.PIPE5_DT_683_net_1\, 
        \I2.PIPE5_DT_6l7r_net_1\, \I2.PIPE5_DT_682_net_1\, 
        \I2.PIPE5_DT_6l6r_net_1\, \I2.PIPE5_DT_681_net_1\, 
        \I2.PIPE5_DT_6l5r_net_1\, \I2.PIPE5_DT_680_net_1\, 
        \I2.PIPE5_DT_6l4r_net_1\, \I2.PIPE5_DT_679_net_1\, 
        \I2.PIPE5_DT_6l3r_net_1\, \I2.PIPE4_DTl2r_net_1\, 
        \I2.PIPE5_DT_678_net_1\, \I2.PIPE5_DT_6l2r_net_1\, 
        \I2.PIPE5_DT_677_net_1\, \I2.PIPE5_DT_6l1r_net_1\, 
        \I2.PIPE4_DTl0r_net_1\, \I2.PIPE5_DT_676_net_1\, 
        \I2.PIPE5_DT_6l0r_net_1\, \I2.FIRST_TDC_675_net_1\, 
        \I2.FIRST_TDC_i_0_i\, \I2.TOKOUT_FL_674_net_1\, 
        \I2.TOKOUT_FL_net_1\, \I2.N_3881\, \I2.TDCGDBi_673_net_1\, 
        \I2.un1_STATE1_24\, \I2.N_3866\, \I2.un6_tdcgdb1_3_net_1\, 
        \I2.un6_tdcgdb1_2_net_1\, \I2.TDCl2r_net_1\, 
        \I2.TDCl3r_net_1\, \I2.un6_tdcgdb1_1_net_1\, 
        \I2.un6_tdcgdb1_0_net_1\, \I2.TDCl0r_net_1\, 
        \I2.TDCl1r_net_1\, \I2.TDCGDAi_672_net_1\, 
        \I2.un1_STATE1_23_net_1\, \I2.un1_STATE1_30_net_1\, 
        \I2.END_TDC1_0_sqmuxa_1_net_1\, \I2.un7_tdcgda1_3_i_i\, 
        \I2.un7_tdcgda1_2_i_i\, \I2.un7_tdcgda1_1_i_i\, 
        \I2.un7_tdcgda1_0_i_i\, \I2.RAMAD1_671_net_1\, 
        \I2.RAMAD1l17r_net_1\, \I2.RAMAD1_670_net_1\, 
        \I2.RAMAD1l16r_net_1\, \I2.RAMAD1_12l16r_net_1\, 
        \I2.RAMAD1_669_net_1\, \I2.RAMAD1l15r_net_1\, 
        \I2.RAMAD1_12l15r_net_1\, \I2.RAMAD1_668_net_1\, 
        \I2.RAMAD1l14r_net_1\, \I2.RAMAD1_12l14r_net_1\, 
        \I2.RAMAD1_667_net_1\, \I2.RAMAD1l13r_net_1\, 
        \I2.RAMAD1_12l13r_net_1\, \I2.RAMAD1_666_net_1\, 
        \I2.RAMAD1l12r_net_1\, \I2.RAMAD1_12l12r_net_1\, 
        \I2.RAMAD1_665_net_1\, \I2.RAMAD1l11r_net_1\, 
        \I2.RAMAD1_12l11r_net_1\, \I2.RAMAD1_664_net_1\, 
        \I2.RAMAD1l10r_net_1\, \I2.RAMAD1_12l10r_net_1\, 
        \I2.RAMAD1_663_net_1\, \I2.RAMAD1l9r_net_1\, 
        \I2.RAMAD1_12l9r_net_1\, \I2.RAMAD1_662_net_1\, 
        \I2.RAMAD1l8r_net_1\, \I2.RAMAD1_12l8r_net_1\, 
        \I2.RAMAD1_661_net_1\, \I2.RAMAD1l7r_net_1\, 
        \I2.RAMAD1_12l7r_net_1\, \I2.RAMAD1_660_net_1\, 
        \I2.RAMAD1l6r_net_1\, \I2.RAMAD1_12l6r_net_1\, 
        \I2.RAMAD1_659_net_1\, \I2.RAMAD1l5r_net_1\, 
        \I2.RAMAD1_12l5r_net_1\, \I2.RAMAD1_658_net_1\, 
        \I2.RAMAD1l4r_net_1\, \I2.RAMAD1_12l4r_net_1\, 
        \I2.RAMAD1_657_net_1\, \I2.RAMAD1l3r_net_1\, 
        \I2.RAMAD1_12l3r_net_1\, \I2.RAMAD1_656_net_1\, 
        \I2.RAMAD1l2r_net_1\, \I2.RAMAD1_12l2r_net_1\, 
        \I2.RAMAD1_655_net_1\, \I2.RAMAD1l1r_net_1\, 
        \I2.RAMAD1_12l1r_net_1\, \I2.STATE1l12r_net_1\, 
        \I2.RAMAD1_654_net_1\, \I2.RAMAD1l0r_net_1\, 
        \I2.RAMAD1_12l0r_net_1\, \I2.TDC_653_net_1\, 
        \I2.TDC_652_net_1\, \I2.TDC_651_net_1\, 
        \I2.TDC_650_net_1\, \I2.TOKENTOB_RES_649_net_1\, 
        \I2.N_3302\, \I2.STATE1l8r_net_1\, 
        \I2.TOKENTOA_RES_648_net_1\, \I2.N_3306\, 
        \I2.NLD_647_net_1\, \I2.un1_STATE3_3\, 
        \I2.EVNT_REJ_646_net_1\, \I2.EVNT_REJ_net_1\, 
        \I2.L2TYPEl0r_net_1\, \I2.L2TYPEl8r_net_1\, 
        \I2.L2TYPEl4r_net_1\, \I2.L2TYPEl12r_net_1\, 
        \I2.L2TYPEl2r_net_1\, \I2.L2TYPEl10r_net_1\, 
        \I2.L2TYPEl6r_net_1\, \I2.L2TYPEl14r_net_1\, 
        \I2.RPAGEl15r\, \I2.L2TYPE_i_0_il1r\, 
        \I2.L2TYPE_i_0_il9r\, \I2.L2TYPE_i_0_il5r\, 
        \I2.L2TYPE_i_0_il13r\, \I2.L2TYPEl3r_net_1\, 
        \I2.L2TYPEl11r_net_1\, \I2.L2TYPEl7r_net_1\, 
        \I2.L2TYPEl15r_net_1\, \I2.LEAD_FLAG6_644_net_1\, 
        \I2.N_4527\, \I2.N_222\, \I2.LEAD_FLAG6_643_net_1\, 
        \I2.LEAD_FLAG6_642_net_1\, \I2.LEAD_FLAG6_641_net_1\, 
        \I2.LEAD_FLAG6_640_net_1\, \I2.PIPE5_DTl22r_net_1\, 
        \I2.LEAD_FLAG6_639_net_1\, \I2.LEAD_FLAG6_638_net_1\, 
        \I2.LEAD_FLAG6_637_net_1\, \I2.PIPE10_DT_636_net_1\, 
        \I2.PIPE9_DTl31r_net_1\, \I2.PIPE10_DT_635_net_1\, 
        \I2.PIPE9_DTl30r_net_1\, \I2.PIPE10_DT_634_net_1\, 
        \I2.PIPE9_DTl29r_net_1\, \I2.SUB9l20r_net_1\, 
        \I2.PIPE10_DT_633_net_1\, \I2.PIPE9_DTl28r_net_1\, 
        \I2.PIPE10_DT_632_net_1\, \I2.PIPE9_DTl27r_net_1\, 
        \I2.PIPE10_DT_631_net_1\, \I2.PIPE9_DTl26r_net_1\, 
        \I2.PIPE10_DT_630_net_1\, \I2.PIPE9_DTl25r_net_1\, 
        \I2.PIPE10_DT_629_net_1\, \I2.PIPE9_DTl24r_net_1\, 
        \I2.PIPE10_DT_628_net_1\, \I2.PIPE9_DTl23r_net_1\, 
        \I2.PIPE10_DT_627_net_1\, \I2.PIPE9_DTl22r_net_1\, 
        \I2.PIPE10_DT_626_net_1\, \I2.PIPE9_DTl21r_net_1\, 
        \I2.PIPE10_DT_625_net_1\, \I2.SUB9l7r_net_1\, 
        \I2.PIPE9_DTl20r_net_1\, \I2.PIPE10_DT_624_net_1\, 
        \I2.SUB9l6r_net_1\, \I2.PIPE9_DTl19r_net_1\, 
        \I2.PIPE10_DT_623_net_1\, \I2.SUB9l5r_net_1\, 
        \I2.PIPE9_DTl18r_net_1\, \I2.PIPE10_DT_622_net_1\, 
        \I2.SUB9l4r_net_1\, \I2.PIPE9_DTl17r_net_1\, 
        \I2.PIPE10_DT_621_net_1\, \I2.SUB9l3r_net_1\, 
        \I2.PIPE9_DTl16r_net_1\, \I2.PIPE10_DT_620_net_1\, 
        \I2.SUB9l2r_net_1\, \I2.PIPE9_DTl15r_net_1\, 
        \I2.PIPE10_DT_619_net_1\, \I2.SUB9l1r_net_1\, 
        \I2.PIPE9_DTl14r_net_1\, \I2.PIPE10_DT_618_net_1\, 
        \I2.SUB9l0r_net_1\, \I2.SUB9_i_0_il17r\, 
        \I2.SUB9l16r_net_1\, \I2.SUB9_i_0_il19r\, 
        \I2.SUB9l18r_net_1\, \I2.SUB9_i_0_il9r\, 
        \I2.SUB9l8r_net_1\, \I2.SUB9_i_0_il11r\, 
        \I2.SUB9l10r_net_1\, \I2.SUB9_i_0_il13r\, 
        \I2.SUB9l12r_net_1\, \I2.SUB9_i_0_il15r\, 
        \I2.SUB9l14r_net_1\, \I2.PIPE9_DTl13r_net_1\, 
        \I2.PIPE10_DT_617_net_1\, \I2.PIPE9_DTl12r_net_1\, 
        \I2.PIPE10_DT_616_net_1\, \I2.PIPE9_DTl11r_net_1\, 
        \I2.PIPE10_DT_615_net_1\, \I2.PIPE9_DTl10r_net_1\, 
        \I2.PIPE10_DT_614_net_1\, \I2.PIPE9_DTl9r_net_1\, 
        \I2.NWPIPE9_0_7\, \I2.PIPE10_DT_613_net_1\, 
        \I2.PIPE9_DTl8r_net_1\, \I2.PIPE10_DT_612_net_1\, 
        \I2.PIPE9_DTl7r_net_1\, \I2.PIPE10_DT_611_net_1\, 
        \I2.PIPE9_DTl6r_net_1\, \I2.PIPE10_DT_610_net_1\, 
        \I2.PIPE9_DTl5r_net_1\, \I2.PIPE10_DT_609_net_1\, 
        \I2.PIPE9_DTl4r_net_1\, \I2.PIPE10_DT_608_net_1\, 
        \I2.PIPE9_DTl3r_net_1\, \I2.PIPE10_DT_607_net_1\, 
        \I2.PIPE9_DTl2r_net_1\, \I2.PIPE10_DT_606_net_1\, 
        \I2.PIPE9_DTl1r_net_1\, \I2.PIPE10_DT_605_net_1\, 
        \I2.PIPE9_DTl0r_net_1\, \I2.L2TYPE_604_net_1\, 
        \I2.L2TYPE_4l15r\, \I2.L2TYPE_603_net_1\, \I2.N_4438\, 
        \I2.L2TYPE_602_net_1\, \I2.N_4439\, \I2.L2TYPE_601_net_1\, 
        \I2.N_4440\, \I2.L2TYPE_600_net_1\, \I2.N_4441\, 
        \I2.L2TYPE_599_net_1\, \I2.N_4442\, \I2.L2TYPE_598_net_1\, 
        \I2.N_4443\, \I2.L2TYPE_597_net_1\, \I2.N_4444\, 
        \I2.L2TYPE_596_net_1\, \I2.N_4445\, \I2.L2TYPE_595_net_1\, 
        \I2.N_4446\, \I2.L2TYPE_594_net_1\, \I2.N_4447\, 
        \I2.L2TYPE_593_net_1\, \I2.N_4448\, \I2.L2TYPE_592_net_1\, 
        \I2.N_4449\, \I2.L2TYPE_591_net_1\, \I2.N_4450\, 
        \I2.L2TYPE_590_net_1\, \I2.N_4451\, \I2.L2TYPE_589_net_1\, 
        \I2.N_4452\, \I2.SUB9_588_net_1\, \I2.SUB8l20r_net_1\, 
        \I2.SUB9_587_net_1\, \I2.N_3562_i\, \I2.SUB9_586_net_1\, 
        \I2.SUB9_585_net_1\, \I2.SUB9_584_net_1\, 
        \I2.SUB9_583_net_1\, \I2.SUB8l14r_net_1\, 
        \I2.SUB9_582_net_1\, \I2.SUB9_581_net_1\, 
        \I2.SUB9_580_net_1\, \I2.SUB8l11r_net_1\, 
        \I2.SUB9_579_net_1\, \I2.SUB9_578_net_1\, 
        \I2.SUB9_577_net_1\, \I2.SUB9_576_net_1\, 
        \I2.SUB9_575_net_1\, \I2.SUB9_574_net_1\, 
        \I2.SUB9_573_net_1\, \I2.SUB9_572_net_1\, 
        \I2.SUB9_571_net_1\, \I2.SUB9_570_net_1\, 
        \I2.SUB9_569_net_1\, \I2.SUB8l2r_net_1\, 
        \I2.SUB9_568_net_1\, \I2.SUB8l1r_net_1\, 
        \I2.PIPE8_DTl29r_net_1\, \I2.PIPE8_DTl31r_net_1\, 
        \I2.OFFSET_567_net_1\, \I2.OFFSET_37l7r\, 
        \I2.OFFSETl7r_net_1\, \I2.un1_NWPIPE7_2_net_1\, 
        \I2.N_746\, \I2.N_858\, \I2.CHA_DATA8_net_1\, \I2.N_690\, 
        \I2.N_738\, \I2.N_658\, \I2.N_682\, \I2.N_642\, 
        \I2.N_650\, \I2.N_666\, \I2.N_674\, \I2.N_714\, 
        \I2.N_730\, \I2.N_698\, \I2.N_706\, \I2.N_722\, 
        \I2.N_802\, \I2.N_850\, \I2.N_770\, \I2.N_794\, 
        \I2.N_754\, \I2.N_762\, \I2.N_778\, \I2.N_786\, 
        \I2.N_826\, \I2.N_842\, \I2.N_810\, \I2.N_818\, 
        \I2.N_834\, \I2.OFFSET_566_net_1\, \I2.OFFSET_37l6r\, 
        \I2.OFFSETl6r_net_1\, \I2.N_745\, \I2.N_857\, \I2.N_689\, 
        \I2.N_737\, \I2.N_657\, \I2.N_681\, \I2.N_641\, 
        \I2.N_649\, \I2.N_665\, \I2.N_673\, \I2.N_713\, 
        \I2.N_729\, \I2.N_697\, \I2.N_705\, \I2.N_721\, 
        \I2.N_801\, \I2.N_849\, \I2.N_769\, \I2.N_793\, 
        \I2.N_753\, \I2.N_761\, \I2.N_777\, \I2.N_785\, 
        \I2.N_825\, \I2.N_841\, \I2.N_809\, \I2.N_817\, 
        \I2.N_833\, \I2.OFFSET_565_net_1\, \I2.OFFSET_37l5r\, 
        \I2.OFFSETl5r_net_1\, \I2.N_744\, \I2.N_856\, \I2.N_688\, 
        \I2.N_736\, \I2.N_656\, \I2.N_680\, \I2.N_640\, 
        \I2.N_648\, \I2.N_664\, \I2.N_672\, \I2.N_712\, 
        \I2.N_728\, \I2.N_696\, \I2.N_704\, \I2.N_720\, 
        \I2.N_800\, \I2.N_848\, \I2.N_768\, \I2.N_792\, 
        \I2.N_752\, \I2.N_760\, \I2.N_776\, \I2.N_784\, 
        \I2.N_824\, \I2.N_840\, \I2.N_808\, \I2.N_816\, 
        \I2.N_832\, \I2.OFFSET_564_net_1\, \I2.OFFSET_37l4r\, 
        \I2.OFFSETl4r_net_1\, \I2.N_743\, \I2.N_855\, \I2.N_687\, 
        \I2.N_735\, \I2.N_655\, \I2.N_679\, \I2.N_639\, 
        \I2.N_647\, \I2.N_663\, \I2.N_671\, \I2.N_711\, 
        \I2.N_727\, \I2.N_695\, \I2.N_703\, \I2.N_719\, 
        \I2.N_799\, \I2.N_847\, \I2.N_767\, \I2.N_791\, 
        \I2.N_751\, \I2.N_759\, \I2.N_775\, \I2.N_783\, 
        \I2.N_823\, \I2.N_839\, \I2.N_807\, \I2.N_815\, 
        \I2.N_831\, \I2.OFFSET_563_net_1\, \I2.OFFSET_37l3r\, 
        \I2.OFFSETl3r_net_1\, \I2.N_742\, \I2.N_854\, \I2.N_686\, 
        \I2.N_734\, \I2.N_654\, \I2.N_678\, \I2.N_638\, 
        \I2.N_646\, \I2.N_662\, \I2.N_670\, \I2.N_710\, 
        \I2.N_726\, \I2.N_694\, \I2.N_702\, \I2.N_718\, 
        \I2.N_798\, \I2.N_846\, \I2.PIPE7_DTl24r_net_1\, 
        \I2.N_766\, \I2.N_790\, \I2.N_750\, \I2.N_758\, 
        \I2.N_774\, \I2.N_782\, \I2.N_822\, \I2.N_838\, 
        \I2.N_806\, \I2.N_814\, \I2.N_830\, \I2.OFFSET_562_net_1\, 
        \I2.OFFSET_37l2r\, \I2.OFFSETl2r_net_1\, \I2.N_741\, 
        \I2.N_853\, \I2.N_685\, \I2.N_733\, \I2.N_653\, 
        \I2.N_677\, \I2.N_637\, \I2.N_645\, \I2.N_661\, 
        \I2.N_669\, \I2.N_709\, \I2.N_725\, \I2.N_693\, 
        \I2.N_701\, \I2.N_717\, \I2.N_797\, \I2.N_845\, 
        \I2.N_765\, \I2.N_789\, \I2.N_749\, \I2.N_757\, 
        \I2.N_773\, \I2.N_781\, \I2.N_821\, \I2.N_837\, 
        \I2.N_805\, \I2.N_813\, \I2.N_829\, \I2.OFFSET_561_net_1\, 
        \I2.OFFSET_37l1r\, \I2.OFFSETl1r_net_1\, \I2.N_740\, 
        \I2.N_852\, \I2.N_684\, \I2.N_732\, \I2.N_652\, 
        \I2.N_676\, \I2.PIPE7_DTl25r_net_1\, \I2.N_636\, 
        \I2.N_644\, \I2.N_660\, \I2.N_668\, \I2.N_708\, 
        \I2.N_724\, \I2.N_692\, \I2.N_700\, \I2.N_716\, 
        \I2.N_796\, \I2.N_844\, \I2.N_764\, \I2.N_788\, 
        \I2.N_748\, \I2.N_756\, \I2.N_772\, \I2.N_780\, 
        \I2.N_820\, \I2.N_836\, \I2.N_804\, \I2.N_812\, 
        \I2.N_828\, \I2.OFFSET_560_net_1\, \I2.OFFSET_37l0r\, 
        \I2.CHB_DATA8_net_1\, \I2.N_739\, \I2.N_851\, \I2.N_683\, 
        \I2.N_731\, \I2.N_651\, \I2.N_675\, \I2.N_635\, 
        \I2.N_643\, \I2.N_659\, \I2.N_667\, \I2.N_707\, 
        \I2.N_723\, \I2.N_691\, \I2.N_699\, \I2.N_715\, 
        \I2.N_795\, \I2.N_843\, \I2.N_763\, \I2.N_787\, 
        \I2.N_747\, \I2.N_755\, \I2.N_771\, \I2.N_779\, 
        \I2.N_819\, \I2.N_835\, \I2.N_803\, \I2.N_811\, 
        \I2.N_827\, \I2.PIPE8_DT_559_net_1\, \I2.N_4418\, 
        \I2.PIPE8_DT_558_net_1\, \I2.PIPE8_DT_557_net_1\, 
        \I2.PIPE8_DT_21l29r\, \I2.PIPE7_DTl29r_net_1\, 
        \I2.PIPE8_DT_556_net_1\, \I2.N_4399\, 
        \I2.PIPE8_DTl28r_net_1\, \I2.PIPE7_DTl28r_net_1\, 
        \I2.PIPE8_DT_21_i_1l28r_net_1\, \I2.LSRAM_OUTl28r\, 
        \I2.PIPE8_DT_555_net_1\, \I2.PIPE8_DT_21l27r_net_1\, 
        \I2.PIPE8_DTl27r_net_1\, \I2.LSRAM_OUTl27r\, 
        \I2.PIPE8_DT_554_net_1\, \I2.PIPE8_DT_21l26r_net_1\, 
        \I2.PIPE8_DTl26r_net_1\, \I2.LSRAM_OUTl26r\, 
        \I2.PIPE8_DT_553_net_1\, \I2.PIPE8_DT_21l25r_net_1\, 
        \I2.PIPE8_DTl25r_net_1\, \I2.LSRAM_OUTl25r\, 
        \I2.PIPE8_DT_552_net_1\, \I2.PIPE8_DT_21l24r_net_1\, 
        \I2.PIPE8_DTl24r_net_1\, \I2.LSRAM_OUTl24r\, 
        \I2.PIPE8_DT_551_net_1\, \I2.PIPE8_DT_21l23r_net_1\, 
        \I2.PIPE8_DTl23r_net_1\, \I2.PIPE7_DTl23r_net_1\, 
        \I2.LSRAM_OUTl23r\, \I2.PIPE8_DT_550_net_1\, 
        \I2.PIPE8_DT_21l22r_net_1\, \I2.PIPE8_DTl22r_net_1\, 
        \I2.PIPE7_DTl22r_net_1\, \I2.LSRAM_OUTl22r\, 
        \I2.PIPE8_DT_549_net_1\, \I2.PIPE8_DT_21l21r_net_1\, 
        \I2.PIPE8_DTl21r_net_1\, \I2.PIPE7_DTl21r_net_1\, 
        \I2.LSRAM_OUTl21r\, \I2.PIPE8_DT_548_net_1\, 
        \I2.PIPE8_DT_21l20r_net_1\, \I2.PIPE8_DTl20r_net_1\, 
        \I2.PIPE8_DT_16l20r_net_1\, \I2.LSRAM_OUTl20r\, 
        \I2.PIPE7_DTl20r_net_1\, \I2.N_4681_i\, 
        \I2.PIPE8_DT_547_net_1\, \I2.PIPE8_DT_21l19r_net_1\, 
        \I2.PIPE8_DTl19r_net_1\, \I2.PIPE8_DT_16l19r_net_1\, 
        \I2.LSRAM_OUTl19r\, \I2.NWPIPE7_net_1\, 
        \I2.PIPE7_DTl19r_net_1\, \I2.PIPE8_DT_546_net_1\, 
        \I2.PIPE8_DT_21l18r_net_1\, \I2.PIPE8_DTl18r_net_1\, 
        \I2.PIPE8_DT_16l18r_net_1\, \I2.LSRAM_OUTl18r\, 
        \I2.PIPE7_DTl18r_net_1\, \I2.PIPE8_DT_545_net_1\, 
        \I2.PIPE8_DT_21l17r_net_1\, \I2.PIPE8_DTl17r_net_1\, 
        \I2.PIPE8_DT_16l17r_net_1\, \I2.LSRAM_OUTl17r\, 
        \I2.PIPE7_DTl17r_net_1\, \I2.PIPE8_DT_544_net_1\, 
        \I2.PIPE8_DT_21l16r_net_1\, \I2.PIPE8_DTl16r_net_1\, 
        \I2.PIPE8_DT_16l16r_net_1\, \I2.LSRAM_OUTl16r\, 
        \I2.PIPE7_DTl16r_net_1\, \I2.PIPE8_DT_543_net_1\, 
        \I2.PIPE8_DT_21l15r_net_1\, \I2.PIPE8_DTl15r_net_1\, 
        \I2.PIPE8_DT_16l15r_net_1\, \I2.LSRAM_OUTl15r\, 
        \I2.PIPE7_DTl15r_net_1\, \I2.PIPE8_DT_542_net_1\, 
        \I2.PIPE8_DT_21l14r_net_1\, \I2.PIPE8_DTl14r_net_1\, 
        \I2.PIPE8_DT_16l14r_net_1\, \I2.LSRAM_OUTl14r\, 
        \I2.PIPE7_DTl14r_net_1\, \I2.PIPE8_DT_541_net_1\, 
        \I2.PIPE8_DT_21l13r_net_1\, \I2.PIPE8_DTl13r_net_1\, 
        \I2.PIPE8_DT_16l13r_net_1\, \I2.LSRAM_OUTl13r\, 
        \I2.PIPE7_DTl13r_net_1\, \I2.PIPE8_DT_540_net_1\, 
        \I2.PIPE8_DT_21l12r_net_1\, \I2.PIPE8_DTl12r_net_1\, 
        \I2.LSRAM_OUTl12r\, \I2.PIPE7_DTl12r_net_1\, 
        \I2.PIPE8_DT_539_net_1\, \I2.PIPE8_DT_21l11r_net_1\, 
        \I2.PIPE8_DTl11r_net_1\, \I2.LSRAM_OUTl11r\, 
        \I2.PIPE7_DTl11r_net_1\, \I2.PIPE8_DT_538_net_1\, 
        \I2.PIPE8_DT_21l10r_net_1\, \I2.PIPE8_DTl10r_net_1\, 
        \I2.LSRAM_OUTl10r\, \I2.PIPE7_DTl10r_net_1\, 
        \I2.PIPE8_DT_537_net_1\, \I2.PIPE8_DT_21l9r_net_1\, 
        \I2.PIPE8_DTl9r_net_1\, \I2.LSRAM_OUTl9r\, 
        \I2.PIPE7_DTl9r_net_1\, \I2.PIPE8_DT_536_net_1\, 
        \I2.PIPE8_DT_21l8r_net_1\, \I2.PIPE8_DTl8r_net_1\, 
        \I2.LSRAM_OUTl8r\, \I2.PIPE7_DTl8r_net_1\, 
        \I2.PIPE8_DT_535_net_1\, \I2.PIPE8_DT_21l7r_net_1\, 
        \I2.PIPE8_DTl7r_net_1\, \I2.LSRAM_OUTl7r\, 
        \I2.PIPE7_DTl7r_net_1\, \I2.PIPE8_DT_534_net_1\, 
        \I2.PIPE8_DT_21l6r_net_1\, \I2.PIPE8_DTl6r_net_1\, 
        \I2.LSRAM_OUTl6r\, \I2.PIPE7_DTl6r_net_1\, 
        \I2.PIPE8_DT_533_net_1\, \I2.PIPE8_DT_21l5r_net_1\, 
        \I2.PIPE8_DTl5r_net_1\, \I2.LSRAM_OUTl5r\, 
        \I2.PIPE7_DTl5r_net_1\, \I2.PIPE8_DT_532_net_1\, 
        \I2.PIPE8_DT_21l4r_net_1\, \I2.PIPE8_DTl4r_net_1\, 
        \I2.LSRAM_OUTl4r\, \I2.PIPE7_DTl4r_net_1\, 
        \I2.PIPE8_DT_531_net_1\, \I2.PIPE8_DT_21l3r_net_1\, 
        \I2.PIPE8_DTl3r_net_1\, \I2.LSRAM_OUTl3r\, 
        \I2.PIPE7_DTl3r_net_1\, \I2.PIPE8_DT_530_net_1\, 
        \I2.PIPE8_DT_21l2r_net_1\, \I2.PIPE8_DTl2r_net_1\, 
        \I2.LSRAM_OUTl2r\, \I2.PIPE7_DTl2r_net_1\, 
        \I2.PIPE8_DT_529_net_1\, \I2.PIPE8_DT_21l1r_net_1\, 
        \I2.PIPE8_DTl1r_net_1\, \I2.LSRAM_OUTl1r\, 
        \I2.PIPE7_DTl1r_net_1\, \I2.PIPE8_DT_528_net_1\, 
        \I2.PIPE8_DT_21l0r_net_1\, \I2.PIPE8_DTl0r_net_1\, 
        \I2.LSRAM_OUTl0r\, \I2.PIPE7_DTl0r_net_1\, 
        \I2.INT_ERRBS_527_net_1\, \I2.INT_ERRBF1_net_1\, 
        \I2.INT_ERRBS_i_i\, \I2.INT_ERRAS_526_net_1\, 
        \I2.INT_ERRAF1_net_1\, \I2.INT_ERRAS_net_1\, 
        \I2.CHAINB_ERRS_525_net_1\, \I2.CHAINB_ERRF1_net_1\, 
        \I2.CHAINA_ERRS_524_net_1\, \I2.CHAINA_ERRF1_net_1\, 
        \I2.SUB8_523_net_1\, \I2.SUB_21x21_fast_I216_Y_0\, 
        \I2.N296_0\, \I2.N288_0\, \I2.N411\, \I2.N297_0\, 
        \I2.N285\, \I2.SUB8l19r_net_1\, 
        \I2.SUB_21x21_fast_I215_Y_0\, \I2.N345\, \I2.N298_0\, 
        \I2.N346_0\, \I2.N299_0\, \I2.N282\, \I2.SUB8_521_net_1\, 
        \I2.SUB8_2l18r\, \I2.N479\, \I2.SUB_21x21_fast_I214_Y_0\, 
        \I2.N300_0\, \I2.N348\, \I2.N301_2\, \I2.N279\, 
        \I2.N_3560_i_net_1\, \I2.SUB_21x21_fast_I213_Y_0\, 
        \I2.N349\, \I2.N302_0\, \I2.N350\, \I2.N303_0\, \I2.N276\, 
        \I2.N_3558_i_net_1\, \I2.SUB8_2_i_i_0l16r\, 
        \I2.I180_un1_Y\, \I2.SUB_21x21_fast_I212_Y_0\, 
        \I2.N304_0\, \I2.N305_0\, \I2.N273\, \I2.SUB8l15r_net_1\, 
        \I2.SUB8_2l15r\, \I2.N486_i\, 
        \I2.SUB_21x21_fast_I211_Y_0\, \I2.I161_un1_Y\, 
        \I2.N306_i_i\, \I2.N353\, \I2.N510\, \I2.N307_2\, 
        \I2.N270_0\, \I2.SUB8_517_net_1\, \I2.SUB8_2l14r\, 
        \I2.N489_i\, \I2.SUB_21x21_fast_I210_Y_0\, 
        \I2.I162_un1_Y\, \I2.N308_0\, \I2.N355_0\, \I2.N513\, 
        \I2.N356\, \I2.N309_0\, \I2.N267_0\, \I2.SUB8l13r_net_1\, 
        \I2.SUB8_2l13r\, \I2.N492_i\, 
        \I2.SUB_21x21_fast_I209_Y_0\, \I2.I163_un1_Y\, 
        \I2.N310_0\, \I2.N357_1\, \I2.N516\, \I2.N311_0\, 
        \I2.N264_0\, \I2.SUB8l12r_net_1\, \I2.SUB8_2l12r\, 
        \I2.N495_i\, \I2.SUB_21x21_fast_I208_Y_0\, \I2.N313_1\, 
        \I2.N312_0\, \I2.N261_0\, \I2.SUB8_514_net_1\, 
        \I2.SUB8_2l11r\, \I2.N498_1\, 
        \I2.SUB_21x21_fast_I207_Y_0\, \I2.N315\, \I2.N314\, 
        \I2.N258_0\, \I2.SUB8_513_net_1\, \I2.SUB8l10r_net_1\, 
        \I2.SUB8_2l10r\, \I2.N501_i\, 
        \I2.SUB_21x21_fast_I206_Y_0\, \I2.N363\, \I2.N317\, 
        \I2.N316_i_i\, \I2.N255_0\, \I2.SUB8_512_net_1\, 
        \I2.SUB8l9r_net_1\, \I2.SUB8_2l9r\, \I2.N504\, 
        \I2.SUB_21x21_fast_I205_Y_0\, \I2.N319_0\, \I2.N318\, 
        \I2.N252_0\, \I2.SUB8_511_net_1\, \I2.SUB8l8r_net_1\, 
        \I2.SUB8_2_i_i_0l8r\, \I2.I168_un1_Y\, 
        \I2.SUB_21x21_fast_I204_Y_0\, \I2.N320\, \I2.N321_0\, 
        \I2.N249_0\, \I2.SUB8_510_net_1\, \I2.SUB8l7r_net_1\, 
        \I2.SUB8_2l7r\, \I2.SUB_21x21_fast_I203_Y_0\, \I2.N323_0\, 
        \I2.N322\, \I2.N246_0\, \I2.N245\, \I2.SUB8_509_net_1\, 
        \I2.SUB8l6r_net_1\, \I2.SUB8_2l6r\, 
        \I2.SUB_21x21_fast_I202_Y_0\, \I2.N325_0\, \I2.N324\, 
        \I2.N243_0\, \I2.N242\, \I2.SUB8_508_net_1\, 
        \I2.SUB8l5r_net_1\, \I2.SUB8_2l5r\, 
        \I2.SUB_21x21_fast_I201_Y_0\, \I2.N326_0\, \I2.N240_0\, 
        \I2.N239\, \I2.SUB8_507_net_1\, \I2.SUB8l4r_net_1\, 
        \I2.SUB8_2l4r\, \I2.SUB_21x21_fast_I200_Y_0\, \I2.N237_0\, 
        \I2.N236\, \I2.SUB8_506_net_1\, \I2.SUB8l3r_net_1\, 
        \I2.SUB8_2l3r\, \I2.SUB_21x21_fast_I199_Y_0\, \I2.N233\, 
        \I2.SUB8_505_net_1\, \I2.SUB8_2l2r\, 
        \I2.SUB_21x21_fast_I198_Y_0\, \I2.SUB8_504_net_1\, 
        \I2.SUB8_2l1r\, \I2.SUB_21x21_fast_I197_Y_0\, 
        \I2.CHB_DATA8_503_net_1\, \I2.CHA_DATA8_502_net_1\, 
        \I2.L_LUT_498_net_1\, \I2.INT_ERRBF1_495_net_1\, 
        \I2.INT_ERRAF1_494_net_1\, \I2.CHAINB_ERRF1_493_net_1\, 
        \I2.CHAINA_ERRF1_492_net_1\, \I2.CHAIN_RDY_490_net_1\, 
        \I2.CHAIN_RDY_net_1\, \I2.N_3494\, 
        \I2.FIFO_END_EVNT_489_net_1\, \I2.DTESl31r_net_1\, 
        \I2.DTESl29r_net_1\, \I2.DTESl28r_net_1\, 
        \I2.DTES_i_0_il30r\, \I2.DTOSl30r_net_1\, 
        \I2.DTOSl28r_net_1\, \I2.DTOS_i_il31r\, 
        \I2.DTOSl29r_net_1\, \I2.SRAM_FULL_488_net_1\, 
        \I2.START_GIRO_net_1\, \I2.N_3823\, \I2.N_132\, 
        \I2.N_128_1\, \I2.SRAM_EVNTl4r_net_1\, 
        \I2.PIPE6_DT_487_net_1\, \I2.LSRAM_RDi_486_net_1\, 
        \I2.LSRAM_RDi_net_1\, \I2.PIPE6_DT_485_net_1\, 
        \I2.PIPE6_DTl31r_net_1\, \I2.PIPE6_DT_484_net_1\, 
        \I2.PIPE6_DTl30r_net_1\, \I2.PIPE6_DT_483_net_1\, 
        \I2.PIPE6_DTl29r_net_1\, \I2.PIPE6_DT_482_net_1\, 
        \I2.PIPE6_DTl28r_net_1\, \I2.PIPE6_DT_481_net_1\, 
        \I2.PIPE6_DT_480_net_1\, \I2.PIPE6_DT_479_net_1\, 
        \I2.PIPE6_DT_478_net_1\, \I2.PIPE6_DT_477_net_1\, 
        \I2.PIPE6_DTl23r_net_1\, \I2.PIPE6_DT_476_net_1\, 
        \I2.PIPE6_DTl22r_net_1\, \I2.PIPE6_DT_475_net_1\, 
        \I2.PIPE6_DTl21r_net_1\, \I2.PIPE6_DT_474_net_1\, 
        \I2.PIPE6_DTl20r_net_1\, \I2.PIPE6_DT_473_net_1\, 
        \I2.PIPE6_DTl19r_net_1\, \I2.PIPE6_DT_472_net_1\, 
        \I2.PIPE6_DTl18r_net_1\, \I2.PIPE6_DT_471_net_1\, 
        \I2.PIPE6_DTl17r_net_1\, \I2.PIPE6_DT_470_net_1\, 
        \I2.PIPE6_DTl16r_net_1\, \I2.PIPE6_DT_469_net_1\, 
        \I2.PIPE6_DTl15r_net_1\, \I2.PIPE6_DT_468_net_1\, 
        \I2.PIPE6_DTl14r_net_1\, \I2.PIPE6_DT_467_net_1\, 
        \I2.PIPE6_DTl13r_net_1\, \I2.PIPE6_DT_466_net_1\, 
        \I2.PIPE6_DTl12r_net_1\, \I2.PIPE6_DT_465_net_1\, 
        \I2.PIPE6_DTl11r_net_1\, \I2.PIPE6_DT_464_net_1\, 
        \I2.PIPE6_DTl10r_net_1\, \I2.PIPE6_DT_463_net_1\, 
        \I2.PIPE6_DTl9r_net_1\, \I2.PIPE6_DT_462_net_1\, 
        \I2.PIPE6_DTl8r_net_1\, \I2.PIPE6_DT_461_net_1\, 
        \I2.PIPE6_DTl7r_net_1\, \I2.PIPE6_DT_460_net_1\, 
        \I2.PIPE6_DTl6r_net_1\, \I2.PIPE6_DT_459_net_1\, 
        \I2.PIPE6_DTl5r_net_1\, \I2.PIPE6_DT_458_net_1\, 
        \I2.PIPE6_DTl4r_net_1\, \I2.PIPE6_DT_457_net_1\, 
        \I2.PIPE6_DTl3r_net_1\, \I2.PIPE6_DT_456_net_1\, 
        \I2.PIPE6_DTl2r_net_1\, \I2.PIPE6_DT_455_net_1\, 
        \I2.PIPE6_DTl1r_net_1\, \I2.PIPE6_DT_454_net_1\, 
        \I2.PIPE6_DTl0r_net_1\, \I2.START_GIRO_451_net_1\, 
        \I2.un1_STATE1_21\, \I2.NWEN_450_net_1\, \I2.N_2989\, 
        \I2.STATE3_i_il10r\, \I2.STATE3_i_il12r\, 
        \I2.STATE3l11r_net_1\, \I2.STATE3l13r_net_1\, 
        \I2.NWPIPE6_449_net_1\, \I2.CHAIN_ERR_DIS_448_net_1\, 
        \I2.TOKENB_TIMOUT_i_i\, \I2.TOKENA_TIMOUT_net_1\, 
        \I2.DTOSl27r_net_1\, \I2.DTESl27r_net_1\, 
        \I2.DTOSl26r_net_1\, \I2.DTESl26r_net_1\, 
        \I2.DTOSl25r_net_1\, \I2.DTESl25r_net_1\, 
        \I2.DTOSl24r_net_1\, \I2.DTESl24r_net_1\, 
        \I2.DTOSl23r_net_1\, \I2.DTESl23r_net_1\, 
        \I2.DTOSl22r_net_1\, \I2.DTESl22r_net_1\, 
        \I2.DTOSl21r_net_1\, \I2.DTESl21r_net_1\, 
        \I2.DTOSl20r_net_1\, \I2.DTESl20r_net_1\, 
        \I2.DTOSl19r_net_1\, \I2.DTESl19r_net_1\, 
        \I2.DTOSl18r_net_1\, \I2.DTESl18r_net_1\, 
        \I2.DTOSl17r_net_1\, \I2.DTESl17r_net_1\, 
        \I2.DTOSl16r_net_1\, \I2.DTESl16r_net_1\, 
        \I2.DTOSl15r_net_1\, \I2.DTESl15r_net_1\, 
        \I2.DTOSl14r_net_1\, \I2.DTESl14r_net_1\, 
        \I2.DTOSl13r_net_1\, \I2.DTESl13r_net_1\, 
        \I2.DTOSl12r_net_1\, \I2.STATE3l2r_net_1\, 
        \I2.DTESl12r_net_1\, \I2.DTOSl11r_net_1\, 
        \I2.DTESl11r_net_1\, \I2.DTOSl10r_net_1\, 
        \I2.DTESl10r_net_1\, \I2.FID_425_net_1\, \I2.FID_7l9r\, 
        \I2.DTOSl9r_net_1\, \I2.DTESl9r_net_1\, 
        \I2.STATE3l3r_net_1\, \I2.FID_424_net_1\, \I2.FID_7l8r\, 
        \I2.DTOSl8r_net_1\, \I2.DTESl8r_net_1\, 
        \I2.FID_423_net_1\, \I2.FID_7l7r\, \I2.DTOSl7r_net_1\, 
        \I2.DTESl7r_net_1\, \I2.FID_422_net_1\, \I2.FID_7l6r\, 
        \I2.DTOSl6r_net_1\, \I2.DTESl6r_net_1\, 
        \I2.FID_421_net_1\, \I2.FID_7_0_ivl5r_net_1\, 
        \I2.DTOSl5r_net_1\, \I2.FID_7_0_iv_0l5r_net_1\, 
        \I2.DTESl5r_net_1\, \I2.FID_420_net_1\, \I2.FID_7l4r\, 
        \I2.DTESl4r_net_1\, \I2.DTOSl4r_net_1\, 
        \I2.FID_419_net_1\, \I2.FID_7l3r\, \I2.DTESl3r_net_1\, 
        \I2.DTOSl3r_net_1\, \I2.FID_418_net_1\, \I2.FID_7l2r\, 
        \I2.DTESl2r_net_1\, \I2.DTOSl2r_net_1\, 
        \I2.FID_417_net_1\, \I2.FID_7_0_ivl1r_net_1\, 
        \I2.DTOSl1r_net_1\, \I2.FID_7_0_iv_0l1r_net_1\, 
        \I2.DTESl1r_net_1\, \I2.FID_416_net_1\, \I2.FID_7l0r\, 
        \I2.DTOSl0r_net_1\, \I2.DTESl0r_net_1\, 
        \I2.ERR_WORDS_RDY_415_net_1\, \I2.LSRAM_IN_414_0_0_net_1\, 
        \I2.LSRAM_INl31r_net_1\, \I2.LSRAM_IN_413_net_1\, 
        \I2.LSRAM_INl29r_net_1\, \I2.LSRAM_IN_412_net_1\, 
        \I2.LSRAM_INl28r_net_1\, \I2.LSRAM_IN_411_net_1\, 
        \I2.LSRAM_INl27r_net_1\, \I2.LSRAM_IN_410_net_1\, 
        \I2.LSRAM_INl26r_net_1\, \I2.LSRAM_IN_409_net_1\, 
        \I2.LSRAM_INl25r_net_1\, \I2.LSRAM_IN_408_net_1\, 
        \I2.LSRAM_INl24r_net_1\, \I2.LSRAM_IN_407_net_1\, 
        \I2.LSRAM_INl23r_net_1\, \I2.LSRAM_IN_406_net_1\, 
        \I2.LSRAM_INl22r_net_1\, \I2.LSRAM_IN_405_net_1\, 
        \I2.LSRAM_INl21r_net_1\, \I2.LSRAM_IN_404_net_1\, 
        \I2.LSRAM_INl20r_net_1\, \I2.LSRAM_IN_403_net_1\, 
        \I2.LSRAM_INl19r_net_1\, \I2.LSRAM_IN_402_net_1\, 
        \I2.LSRAM_INl18r_net_1\, \I2.LSRAM_IN_401_net_1\, 
        \I2.LSRAM_INl17r_net_1\, \I2.LSRAM_IN_400_net_1\, 
        \I2.LSRAM_INl16r_net_1\, \I2.LSRAM_IN_399_net_1\, 
        \I2.LSRAM_INl15r_net_1\, \I2.LSRAM_IN_398_net_1\, 
        \I2.LSRAM_INl14r_net_1\, \I2.LSRAM_IN_397_net_1\, 
        \I2.LSRAM_INl13r_net_1\, \I2.LSRAM_IN_396_net_1\, 
        \I2.LSRAM_INl12r_net_1\, \I2.LSRAM_IN_395_net_1\, 
        \I2.LSRAM_INl11r_net_1\, \I2.LSRAM_IN_394_net_1\, 
        \I2.LSRAM_INl10r_net_1\, \I2.LSRAM_IN_393_net_1\, 
        \I2.LSRAM_INl9r_net_1\, \I2.LSRAM_IN_392_net_1\, 
        \I2.LSRAM_INl8r_net_1\, \I2.LSRAM_IN_391_net_1\, 
        \I2.LSRAM_INl7r_net_1\, \I2.LSRAM_IN_390_net_1\, 
        \I2.LSRAM_INl6r_net_1\, \I2.LSRAM_IN_389_net_1\, 
        \I2.LSRAM_INl5r_net_1\, \I2.LSRAM_IN_388_net_1\, 
        \I2.LSRAM_INl4r_net_1\, \I2.LSRAM_IN_387_net_1\, 
        \I2.LSRAM_INl3r_net_1\, \I2.LSRAM_IN_386_net_1\, 
        \I2.LSRAM_INl2r_net_1\, \I2.LSRAM_IN_385_net_1\, 
        \I2.LSRAM_INl1r_net_1\, \I2.LSRAM_IN_384_net_1\, 
        \I2.LSRAM_INl0r_net_1\, \I2.LSRAM_WADDR_383_net_1\, 
        \I2.LSRAM_WADDRl2r_net_1\, \I2.LSRAM_WADDR_382_net_1\, 
        \I2.LSRAM_WADDRl1r_net_1\, \I2.LSRAM_WADDR_381_net_1\, 
        \I2.LSRAM_WADDRl0r_net_1\, \I2.LSRAM_WR_380_net_1\, 
        \I2.LSRAM_WR_net_1\, \I2.MTDCRESB_379_net_1\, 
        \I2.MTDCRESA_378_net_1\, \I2.NPRSFIF_328_net_1\, 
        \I2.PIPE9_DT_300_net_1\, \I2.PIPE9_DT_299_net_1\, 
        \I2.PIPE9_DT_298_net_1\, \I2.PIPE9_DT_297_net_1\, 
        \I2.PIPE9_DT_296_net_1\, \I2.PIPE9_DT_295_net_1\, 
        \I2.PIPE9_DT_294_net_1\, \I2.PIPE9_DT_293_net_1\, 
        \I2.PIPE9_DT_292_net_1\, \I2.PIPE9_DT_291_net_1\, 
        \I2.PIPE9_DT_290_net_1\, \I2.PIPE9_DT_289_net_1\, 
        \I2.PIPE9_DT_288_net_1\, \I2.PIPE9_DT_287_net_1\, 
        \I2.PIPE9_DT_286_net_1\, \I2.PIPE9_DT_285_net_1\, 
        \I2.PIPE9_DT_284_net_1\, \I2.PIPE9_DT_283_net_1\, 
        \I2.PIPE9_DT_282_net_1\, \I2.PIPE9_DT_281_net_1\, 
        \I2.PIPE9_DT_280_net_1\, \I2.PIPE9_DT_279_net_1\, 
        \I2.PIPE9_DT_278_net_1\, \I2.PIPE9_DT_277_net_1\, 
        \I2.PIPE9_DT_276_net_1\, \I2.PIPE9_DT_275_net_1\, 
        \I2.PIPE9_DT_274_net_1\, \I2.PIPE9_DT_273_net_1\, 
        \I2.PIPE9_DT_272_net_1\, \I2.PIPE9_DT_271_net_1\, 
        \I2.PIPE9_DT_270_net_1\, \I2.PIPE9_DT_269_net_1\, 
        \I2.END_EVNT6_net_1\, \I2.TDCTRGi_266_net_1\, 
        \I2.STATE4_il0r\, \I2.TRGARRl3r_net_1\, 
        \I2.TRGARRl0r_net_1\, \I2.TRGCNT_n0_net_1\, 
        \I2.TRGCNT_n0_0_net_1\, \I2.SRAM_EVNT_n4_net_1\, 
        \I2.N_3828\, \I2.SRAM_EVNT_n4_0_net_1\, 
        \I2.SRAM_EVNTl3r_net_1\, \I2.SRAM_EVNT_n3_net_1\, 
        \I2.N_3827\, \I2.SRAM_EVNT_n3_0_net_1\, 
        \I2.SRAM_EVNTl2r_net_1\, \I2.N_135\, 
        \I2.SRAM_EVNT_n2_net_1\, \I2.N_3826\, 
        \I2.SRAM_EVNT_n2_0_net_1\, \I2.SRAM_EVNTl0r_net_1\, 
        \I2.SRAM_EVNTl1r_net_1\, \I2.SRAM_EVNT_n1_net_1\, 
        \I2.N_3825\, \I2.SRAM_EVNT_n1_0_net_1\, 
        \I2.SRAM_EVNT_n0_net_1\, \I2.SRAM_EVNT_n0_0_net_1\, 
        \I2.RAMAD_4l17r_net_1\, \I2.N_544\, 
        \I2.RAMAD_4l16r_net_1\, \I2.N_543\, 
        \I2.RAMAD_4l15r_net_1\, \I2.N_542\, 
        \I2.RAMAD_4l14r_net_1\, \I2.N_541\, 
        \I2.RAMAD_4l13r_net_1\, \I2.N_540\, 
        \I2.RAMAD_4l12r_net_1\, \I2.N_539\, 
        \I2.RAMAD_4l11r_net_1\, \I2.N_538\, 
        \I2.RAMAD_4l10r_net_1\, \I2.N_537\, \I2.RAMAD_4l9r_net_1\, 
        \I2.N_536\, \I2.RAMAD_4l8r_net_1\, \I2.N_535\, 
        \I2.RAMAD_4l7r_net_1\, \I2.N_534\, \I2.RAMAD_4l6r_net_1\, 
        \I2.N_533\, \I2.RAMAD_4l5r_net_1\, \I2.N_532\, 
        \I2.RAMAD_4l4r_net_1\, \I2.N_531\, \I2.RAMAD_4l3r_net_1\, 
        \I2.N_530\, \I2.RAMAD_4l2r_net_1\, \I2.N_529\, 
        \I2.RAMAD_4l1r_net_1\, \I2.N_528\, \I2.RAMAD_4l0r_net_1\, 
        \I2.N_527\, \I2.TOKENB_CNT_3l1r\, \I2.I_10\, 
        \I2.TOKENB_CNT_3l0r\, \I2.DWACT_ADD_CI_0_partial_suml0r\, 
        \I2.TOKENA_CNT_4l1r_net_1\, \I2.I_10_0\, 
        \I2.TOKENA_CNT_4l0r_net_1\, 
        \I2.DWACT_ADD_CI_0_partial_sum_0l0r\, 
        \I2.TOKENB_TIMOUT_2\, \I2.TOKENB_CNTl0r_net_1\, 
        \I2.TOKENB_CNTl1r_net_1\, \I2.TOKENA_TIMOUT_2_net_1\, 
        \I2.TOKENA_CNTl0r_net_1\, \I2.TOKENA_CNTl1r_net_1\, 
        \I2.LSRAM_RD_net_1\, \I2.PLL_LOCK_sram\, 
        \I2.PLL_LOCK_tdc\, \I2.MSERCLKF1_net_1\, 
        \I2.MTDIAF1_net_1\, \I2.L1AF1_net_1\, \I2.L2AF1_net_1\, 
        \I2.L2RF1_net_1\, \I2.END_TDC2_net_1\, 
        \I2.END_EVNT4_net_1\, \I2.END_EVNT3_net_1\, 
        \I2.END_TDC4_net_1\, \I2.END_TDC3_net_1\, 
        \I2.END_EVNT9_net_1\, \I2.END_EVNT8_net_1\, 
        \I2.END_EVNT7_net_1\, \I2.I_5_1\, \I2.BNC_IDl2r_net_1\, 
        \I2.I_9_1\, \I2.I_13_2\, \I2.BNC_IDl4r_net_1\, 
        \I2.I_20_0\, \I2.BNC_IDl5r_net_1\, \I2.I_24_0\, 
        \I2.BNC_IDl6r_net_1\, \I2.I_31_0\, \I2.BNC_IDl7r_net_1\, 
        \I2.I_38_0\, \I2.I_45_0\, \I2.BNC_IDl9r_net_1\, 
        \I2.I_52_0\, \I2.BNC_IDl10r_net_1\, \I2.I_56_0\, 
        \I2.BNC_IDl11r_net_1\, \I2.I_66_0\, 
        \I2.STATEe_illegalpipe1_net_1\, \I2.N_3457_ip\, 
        \I2.PIPE3_DTl0r_net_1\, \I2.PIPE3_DTl1r_net_1\, 
        \I2.PIPE3_DTl2r_net_1\, \I2.PIPE3_DTl3r_net_1\, 
        \I2.PIPE3_DTl4r_net_1\, \I2.PIPE3_DTl5r_net_1\, 
        \I2.PIPE3_DTl6r_net_1\, \I2.PIPE3_DTl7r_net_1\, 
        \I2.PIPE3_DTl9r_net_1\, \I2.PIPE3_DTl10r_net_1\, 
        \I2.PIPE3_DTl11r_net_1\, \I2.PIPE3_DTl12r_net_1\, 
        \I2.PIPE3_DTl13r_net_1\, \I2.PIPE3_DTl14r_net_1\, 
        \I2.PIPE3_DTl15r_net_1\, \I2.PIPE3_DTl16r_net_1\, 
        \I2.PIPE3_DTl17r_net_1\, \I2.PIPE3_DTl18r_net_1\, 
        \I2.PIPE3_DTl19r_net_1\, \I2.PIPE3_DTl20r_net_1\, 
        \I2.PIPE3_DTl21r_net_1\, \I2.PIPE3_DTl22r_net_1\, 
        \I2.PIPE3_DTl23r_net_1\, \I2.PIPE3_DTl24r_net_1\, 
        \I2.PIPE3_DTl25r_net_1\, \I2.PIPE3_DTl26r_net_1\, 
        \I2.PIPE3_DTl27r_net_1\, \I2.PIPE3_DTl28r_net_1\, 
        \I2.PIPE3_DTl29r_net_1\, \I2.PIPE3_DTl30r_net_1\, 
        \I2.PIPE3_DTl31r_net_1\, \I2.DWACT_ADD_CI_0_TMP_1l0r\, 
        \I2.DWACT_ADD_CI_0_TMP_2l0r\, \I2.N_9_1\, \I2.N_16_1\, 
        \I2.N_29\, \I2.N_34\, \I2.N_39\, \I2.N_4_0\, \I2.N_11_1\, 
        \I2.N_24_1\, \I2.N_29_0\, \I2.N_34_0\, \I1.N_435_1\, 
        \FBOUTl0r\, \I1.sstate_ns_i_0_a4_0_1l0r\, \I1.N_292\, 
        \I1.sstate_ns_il5r\, \I1.sstatel3r_net_1\, 
        \I1.sstatel6r_net_1\, \I1.sstatel4r_net_1\, 
        \I1.sstatel5r_net_1\, \I1.sstate_nsl4r\, 
        \I1.COMMAND_net_1\, \I1.sstate_nsl7r\, \I1.N_370\, 
        \I1.N_436_i_i\, \I1.N_186\, \I1.N_405\, 
        \I1.NWRLUTi_57_net_1\, \I1.NWRLUTi_net_1\, \I1.N_1192\, 
        \I1.COMMAND_52_0\, \I1.NOELUTi_51_net_1\, \I3.N_1311_0\, 
        \I3.N_1310_i_0\, \I3.ASBSF1_net_1\, \I3.STATE1_ipl9r\, 
        \I3.STATE1_nsl1r\, \I3.EVREAD_DS_124_net_1\, 
        \I3.STATE1_ipl8r\, \I3.STATE1_nsl2r\, \I3.STATE1_nsl8r\, 
        \I3.N_1906_i_0_0\, \I3.WRITES_net_1\, 
        \I3.PULSE_330_net_1\, \I3.DSS_net_1\, \I3.DSSF1_net_1\, 
        \I3.SINGCYC_115_net_1\, \I3.BLTCYC_113_net_1\, 
        \I3.WRITES_23_net_1\, \I3.REGMAPl10r_net_1\, 
        \I3.STATE2l0r_net_1\, \I3.NRDMEBi_0_sqmuxa_net_1\, 
        \I3.STATE2l2r_net_1\, \I3.N_1896\, \I3.N_90_i_0_1\, 
        \I3.REGMAPl0r_net_1\, \I3.TCNT_0_sqmuxa_0\, 
        \I3.REGMAPl51r_net_1\, \I3.N_276\, \I3.REGMAPl1r_net_1\, 
        \I3.N_12180_i\, \I3.N_1905_1\, \I3.N_98_0\, 
        \I3.REGMAPl13r_net_1\, \I3.REG3l7r_net_1\, 
        \I3.TCNTl4r_net_1\, \I3.VSEL_0\, \I3.N_1918\, 
        \I3.N_1463_i_1\, \I3.REG3l5r_net_1\, \I3.REG2l5r_net_1\, 
        \I3.un7_cycs_i_net_1\, \I3.un7_cycs_0_a3_0_a3_net_1\, 
        \I3.N_2137_i_0\, \I3.MBLTCYC_net_1\, \I3.ADACKCYC_net_1\, 
        \I3.N_290\, \I3.N_95\, \I3.CLOSEDTK_net_1\, \I3.N_284\, 
        \I3.VDBil5r_net_1\, \I3.PIPEBl5r_net_1\, 
        \I3.PIPEAl5r_net_1\, \I3.STATE1_tr24_i_0_net_1\, 
        \I3.STATE1_tr24_i_0_o2_1_i\, \I3.WRITES_8\, \I3.N_303\, 
        \I3.VDBil7r_net_1\, \I3.N_129\, \I3.PIPEBl7r_net_1\, 
        \I3.PIPEAl7r_net_1\, \I3.STATE2_ns_i_i_a5_0_a3l1r_net_1\, 
        \I3.N_258\, \I3.N_1622_1\, \I3.un6_asb_NE_net_1\, 
        \I3.N_262_i_0\, \I3.N_261_i_0\, \I3.N_260_i_0\, 
        \I3.N_186_i_0\, \I3.STATE1_nsl0r\, \I3.STATE1l10r_net_1\, 
        \I3.DSS_9\, \I3.STATE2_nsl4r\, \I3.N_1465\, 
        \I3.STATE2l1r_net_1\, \I3.N_1879\, 
        \I3.STATE2_nsl3r_net_1\, \I3.N_281\, \I3.STATE2_nsl0r\, 
        \I3.EVREAD_DS_net_1\, \I3.STATE1_nsl7r\, 
        \I3.STATE1_nsl6r\, \I3.N_1920\, \I3.STATE1_nsl5r\, 
        \I3.STATE1_nsl4r\, \I3.N_1516\, \I3.STATE1_nsl3r\, 
        \I3.N_1189\, \I3.N_1186\, \I3.STATE1_ipl1r\, \I3.N_1180\, 
        \I3.STATE1_ipl4r\, \I3.N_1174\, \I3.STATE1_ipl5r\, 
        \I3.STATE1_ipl6r\, \I3.N_1168\, \I3.STATE1_ipl7r\, 
        \I3.STATE1_IPL8R_10\, \I3.STATE1_IPL9R_11\, 
        \I3.TCNT_384_net_1\, \I3.TCNTl0r_net_1\, \I3.TCNT_n0\, 
        \I3.TCNTe\, \I3.un1_STATE1_10_i_0\, \I3.N_1966_1\, 
        \I3.TCNT_383_net_1\, \I3.TCNTl1r_net_1\, \I3.TCNT_n1\, 
        \I3.TCNT_382_net_1\, \I3.TCNTl2r_net_1\, \I3.TCNT_n2\, 
        \I3.TCNT_381_net_1\, \I3.TCNTl3r_net_1\, \I3.TCNT_n3\, 
        \I3.TCNT_380_net_1\, \I3.TCNT_n4\, \I3.REG_1_sqmuxa_3\, 
        \I3.VDBi_371_net_1\, \I3.VDBi_57l31r\, 
        \I3.VDBil31r_net_1\, \I3.VDBi_31l31r_net_1\, \I3.N_1905\, 
        \I3.VDBi_20l31r\, \I3.REGl164r\, \I3.PIPEAl31r_net_1\, 
        \I3.VDBi_370_net_1\, \I3.VDBi_57l30r\, 
        \I3.VDBil30r_net_1\, \I3.VDBi_31l30r_net_1\, 
        \I3.VDBi_20l30r\, \I3.REGl163r\, \I3.PIPEAl30r_net_1\, 
        \I3.VDBi_369_net_1\, \I3.VDBi_57l29r\, 
        \I3.VDBil29r_net_1\, \I3.VDBi_31l29r_net_1\, 
        \I3.VDBi_20l29r\, \I3.REGl162r\, \I3.PIPEAl29r_net_1\, 
        \I3.VDBi_368_net_1\, \I3.VDBi_57l28r\, 
        \I3.VDBil28r_net_1\, \I3.VDBi_31l28r_net_1\, 
        \I3.VDBi_20l28r\, \I3.REGl161r\, \I3.PIPEAl28r_net_1\, 
        \I3.VDBi_367_net_1\, \I3.VDBi_57l27r\, 
        \I3.VDBil27r_net_1\, \I3.N_1839\, \I3.REGl160r\, 
        \I3.N_1917\, \I3.PIPEAl27r_net_1\, \I3.VDBi_366_net_1\, 
        \I3.VDBi_57l26r\, \I3.VDBil26r_net_1\, 
        \I3.VDBi_31l26r_net_1\, \I3.VDBi_20l26r\, \I3.REGl159r\, 
        \I3.PIPEAl26r_net_1\, \I3.VDBi_365_net_1\, 
        \I3.VDBi_57l25r\, \I3.VDBil25r_net_1\, 
        \I3.VDBi_31l25r_net_1\, \I3.VDBi_20l25r\, \I3.REGl158r\, 
        \I3.PIPEAl25r_net_1\, \I3.VDBi_364_net_1\, 
        \I3.VDBi_57l24r\, \I3.VDBil24r_net_1\, \I3.REGl157r\, 
        \I3.PIPEAl24r_net_1\, \I3.VDBi_363_net_1\, 
        \I3.VDBi_57l23r\, \I3.VDBil23r_net_1\, 
        \I3.VDBi_31l23r_net_1\, \I3.VDBi_20l23r\, \I3.REGl156r\, 
        \I3.PIPEAl23r_net_1\, \I3.VDBi_362_net_1\, 
        \I3.VDBi_57l22r\, \I3.VDBil22r_net_1\, 
        \I3.VDBi_31l22r_net_1\, \I3.VDBi_20l22r\, \I3.REGl155r\, 
        \I3.PIPEAl22r_net_1\, \I3.VDBi_361_net_1\, 
        \I3.VDBi_57l21r\, \I3.VDBil21r_net_1\, \I3.REGl154r\, 
        \I3.PIPEAl21r_net_1\, \I3.VDBi_360_net_1\, 
        \I3.VDBi_57l20r\, \I3.VDBil20r_net_1\, \I3.REGl153r\, 
        \I3.PIPEAl20r_net_1\, \I3.VDBi_359_net_1\, 
        \I3.VDBi_57l19r\, \I3.VDBil19r_net_1\, \I3.REGl152r\, 
        \I3.PIPEAl19r_net_1\, \I3.VDBi_358_net_1\, 
        \I3.VDBi_57l18r\, \I3.VDBil18r_net_1\, \I3.REGl151r\, 
        \I3.PIPEAl18r_net_1\, \I3.VDBi_357_net_1\, 
        \I3.VDBi_57l17r\, \I3.VDBil17r_net_1\, 
        \I3.VDBi_31l17r_net_1\, \I3.VDBi_20l17r\, \I3.REGl150r\, 
        \I3.PIPEAl17r_net_1\, \I3.VDBi_356_net_1\, 
        \I3.VDBi_57l16r\, \I3.VDBil16r_net_1\, 
        \I3.VDBi_31l16r_net_1\, \I3.VDBi_20l16r\, \I3.REGl149r\, 
        \I3.PIPEAl16r_net_1\, \I3.VDBi_355_net_1\, 
        \I3.VDBi_57l15r\, \I3.VDBil15r_net_1\, \I3.N_403_1\, 
        \I3.N_402_1\, \I3.PIPEAl15r_net_1\, \I3.REGl148r\, 
        \I3.N_2058\, \I3.VDBi_354_net_1\, \I3.VDBi_57l14r\, 
        \I3.VDBil14r_net_1\, \I3.PIPEAl14r_net_1\, \I3.N_352\, 
        \I3.VDBi_31l14r_net_1\, \I3.VDBi_20l14r\, \I3.REGl147r\, 
        \I3.VDBi_353_net_1\, \I3.VDBi_57l13r\, 
        \I3.VDBil13r_net_1\, \I3.N_2034\, \I3.RAMDTSl13r_net_1\, 
        \I3.REGl146r\, \I3.PIPEAl13r_net_1\, \I3.N_2276\, 
        \I3.N_56\, \I3.VDBi_352_net_1\, \I3.VDBi_57l12r\, 
        \I3.VDBil12r_net_1\, \I3.VDBi_40l12r_net_1\, \I3.N_1857\, 
        \I3.N_350\, \I3.VDBi_31l12r_net_1\, \I3.VDBi_20l12r\, 
        \I3.REGl145r\, \I3.N_280\, \I3.PIPEAl12r_net_1\, 
        \I3.VDBi_351_net_1\, \I3.VDBi_57l11r\, 
        \I3.VDBil11r_net_1\, \I3.VDBi_43l11r_net_1\, 
        \I3.VDBi_40l11r_net_1\, \I3.N_1856\, \I3.N_349\, 
        \I3.VDBi_31l11r_net_1\, \I3.VDBi_20l11r\, \I3.REGl144r\, 
        \I3.N_278\, \I3.PIPEAl11r_net_1\, \I3.VDBi_350_net_1\, 
        \I3.VDBi_57l10r\, \I3.VDBil10r_net_1\, 
        \I3.VDBi_43l10r_net_1\, \I3.VDBi_40l10r_net_1\, 
        \I3.N_1855\, \I3.N_348\, \I3.VDBi_31l10r_net_1\, 
        \I3.VDBi_20l10r\, \I3.REGl143r\, \I3.N_2261\, 
        \I3.PIPEAl10r_net_1\, \I3.VDBi_349_net_1\, 
        \I3.VDBi_57l9r\, \I3.VDBil9r_net_1\, 
        \I3.VDBi_43l9r_net_1\, \I3.VDBi_40l9r_net_1\, \I3.N_1854\, 
        \I3.N_347\, \I3.VDBi_31l9r_net_1\, \I3.VDBi_29l9r\, 
        \I3.REGl142r\, \I3.REGl100r\, \I3.REGMAPl14r_net_1\, 
        \I3.N_90_i_0\, \I3.PIPEAl9r_net_1\, \I3.VDBi_348_net_1\, 
        \I3.VDBi_57l8r\, \I3.VDBil8r_net_1\, \I3.RAMDTSl8r_net_1\, 
        \I3.PIPEAl8r_net_1\, \I3.N_2271\, \I3.REGl141r\, 
        \I3.VDBi_29l8r_net_1\, \I3.VDBi_20l8r\, \I3.REGl99r\, 
        \I3.VDBi_16l8r_net_1\, \I3.VDBi_10l8r_net_1\, 
        \I3.REGMAPl2r_net_1\, \I3.VDBi_347_net_1\, 
        \I3.VDBi_57l7r\, \I3.VDBoffl7r_net_1\, 
        \I3.RAMDTSl7r_net_1\, \I3.N_2047\, \I3.N_2048\, 
        \I3.REGl98r\, \I3.REGl140r\, \I3.N_2270\, 
        \I3.REG1l7r_net_1\, \I3.REG2l7r_net_1\, 
        \I3.VDBi_346_net_1\, \I3.VDBi_57l6r\, \I3.VDBil6r_net_1\, 
        \I3.VDBoffl6r_net_1\, \I3.PIPEAl6r_net_1\, 
        \I3.RAMDTSl6r_net_1\, \I3.REGl97r\, \I3.REGl139r\, 
        \I3.N_2269\, \I3.REG3l6r_net_1\, \I3.REG1l6r_net_1\, 
        \I3.REG2l6r_net_1\, \I3.VDBi_345_net_1\, \I3.VDBi_57l5r\, 
        \I3.VDBoffl5r_net_1\, \I3.RAMDTSl5r_net_1\, 
        \I3.VDBi_43l5r_net_1\, \I3.VDBi_40l5r\, \I3.N_137\, 
        \I3.N_1948\, \I3.REGl96r\, \I3.N_282_i_i\, \I3.N_283\, 
        \I3.REG1l5r_net_1\, \I3.REGl138r\, \I3.VDBi_344_net_1\, 
        \I3.VDBi_57l4r\, \I3.VDBil4r_net_1\, 
        \I3.VDBi_43l4r_net_1\, \I3.VDBi_40l4r_net_1\, \I3.N_136\, 
        \I3.N_342\, \I3.VDBi_31l4r_net_1\, \I3.VDBi_29l4r_net_1\, 
        \I3.REGl137r\, \I3.REGl95r\, \I3.REGMAPl3r_net_1\, 
        \I3.VDBoffl4r_net_1\, \I3.PIPEAl4r_net_1\, 
        \I3.VDBi_343_net_1\, \I3.VDBi_57l3r\, \I3.VDBil3r_net_1\, 
        \I3.VDBi_43l3r_net_1\, \I3.VDBi_40l3r_net_1\, \I3.N_135\, 
        \I3.N_341\, \I3.VDBi_31l3r_net_1\, \I3.VDBi_29l3r_net_1\, 
        \I3.REGl136r\, \I3.REGl94r\, \I3.VDBoffl3r_net_1\, 
        \I3.PIPEAl3r_net_1\, \I3.VDBi_342_net_1\, \I3.VDBi_57l2r\, 
        \I3.VDBil2r_net_1\, \I3.VDBoffl2r_net_1\, 
        \I3.PIPEAl2r_net_1\, \I3.REGMAPl8r_net_1\, 
        \I3.RAMDTSl2r_net_1\, \I3.REGl93r\, \I3.REGl135r\, 
        \I3.N_134\, \I3.REG1l2r_net_1\, \I3.REG3l2r_net_1\, 
        \I3.REG2l2r_net_1\, \I3.VDBi_341_net_1\, \I3.VDBi_57l1r\, 
        \I3.VDBil1r_net_1\, \I3.VDBi_43l1r_net_1\, 
        \I3.VDBi_40l1r_net_1\, \I3.N_133\, \I3.N_339\, 
        \I3.VDBi_31l1r_net_1\, \I3.REGl134r\, \I3.REGl92r\, 
        \I3.REGMAPl11r_net_1\, \I3.REG1l1r_net_1\, 
        \I3.REG3l1r_net_1\, \I3.REG2l1r_net_1\, 
        \I3.VDBoffl1r_net_1\, \I3.PIPEAl1r_net_1\, 
        \I3.VDBi_340_net_1\, \I3.VDBi_57l0r\, \I3.VDBil0r_net_1\, 
        \I3.REGMAPl50r_net_1\, \I3.REGMAP_i_0_il5r\, 
        \I3.REGMAPl4r_net_1\, \I3.REGMAP_i_0_il15r\, 
        \I3.REGMAPl6r_net_1\, \I3.REGMAPl56r_net_1\, 
        \I3.VDBoffl0r_net_1\, \I3.PIPEAl0r_net_1\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r\, 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_net_1\, \I3.N_1923\, 
        \I3.N_2063_i\, \I3.REG1l0r_net_1\, \I3.REG2l0r_net_1\, 
        \I3.REG3l0r_net_1\, \I3.REG1l405r_net_1\, 
        \I3.REG3l405r_net_1\, \I3.REG2l405r_net_1\, \I3.REGl91r\, 
        \I3.REGl133r\, \I3.N_132\, \I3.REGMAPl12r_net_1\, 
        \I3.RAMDTSl0r_net_1\, \I3.PULSE_339_net_1\, 
        \I3.PULSE_46l9r\, \I3.PULSE_338_net_1\, \I3.PULSE_46l8r\, 
        \I3.PULSE_337_net_1\, \I3.N_1897\, \I3.N_318\, 
        \I3.PULSE_336_net_1\, \I3.PULSE_46l6r\, 
        \I3.PULSE_335_net_1\, \I3.PULSE_46l5r\, 
        \I3.PULSE_334_net_1\, \I3.N_55\, \I3.PULSE_333_net_1\, 
        \I3.N_49\, \I3.PULSE_332_net_1\, \I3.PULSE_331_net_1\, 
        \I3.PIPEA1_329_net_1\, \I3.PIPEA1_12l31r_net_1\, 
        \I3.PIPEA1l31r_net_1\, \I3.PIPEA1_328_net_1\, 
        \I3.PIPEA1_12l30r_net_1\, \I3.PIPEA1l30r_net_1\, 
        \I3.PIPEA1_327_net_1\, \I3.PIPEA1_12l29r_net_1\, 
        \I3.PIPEA1l29r_net_1\, \I3.PIPEA1_326_net_1\, 
        \I3.PIPEA1_12l28r_net_1\, \I3.PIPEA1l28r_net_1\, 
        \I3.PIPEA1_325_net_1\, \I3.PIPEA1_12l27r_net_1\, 
        \I3.PIPEA1l27r_net_1\, \I3.PIPEA1_324_net_1\, 
        \I3.PIPEA1_12l26r_net_1\, \I3.PIPEA1l26r_net_1\, 
        \I3.PIPEA1_323_net_1\, \I3.PIPEA1_12l25r_net_1\, 
        \I3.PIPEA1l25r_net_1\, \I3.PIPEA1_322_net_1\, 
        \I3.PIPEA1_12l24r_net_1\, \I3.PIPEA1l24r_net_1\, 
        \I3.PIPEA1_321_net_1\, \I3.PIPEA1_12l23r_net_1\, 
        \I3.PIPEA1l23r_net_1\, \I3.PIPEA1_320_net_1\, 
        \I3.PIPEA1_12l22r_net_1\, \I3.PIPEA1l22r_net_1\, 
        \I3.PIPEA1_319_net_1\, \I3.PIPEA1_12l21r_net_1\, 
        \I3.PIPEA1l21r_net_1\, \I3.PIPEA1_318_net_1\, 
        \I3.PIPEA1_12l20r_net_1\, \I3.PIPEA1l20r_net_1\, 
        \I3.PIPEA1_317_net_1\, \I3.PIPEA1_12l19r_net_1\, 
        \I3.PIPEA1l19r_net_1\, \I3.PIPEA1_316_net_1\, 
        \I3.PIPEA1_12l18r_net_1\, \I3.PIPEA1l18r_net_1\, 
        \I3.PIPEA1_315_net_1\, \I3.PIPEA1_12l17r_net_1\, 
        \I3.PIPEA1l17r_net_1\, \I3.PIPEA1_314_net_1\, 
        \I3.PIPEA1_12l16r_net_1\, \I3.PIPEA1l16r_net_1\, 
        \I3.PIPEA1_313_net_1\, \I3.PIPEA1_12l15r_net_1\, 
        \I3.PIPEA1l15r_net_1\, \I3.PIPEA1_312_net_1\, 
        \I3.PIPEA1_12l14r_net_1\, \I3.PIPEA1l14r_net_1\, 
        \I3.PIPEA1_311_net_1\, \I3.PIPEA1_12l13r_net_1\, 
        \I3.PIPEA1l13r_net_1\, \I3.PIPEA1_310_net_1\, 
        \I3.PIPEA1_12l12r_net_1\, \I3.PIPEA1l12r_net_1\, 
        \I3.PIPEA1_309_net_1\, \I3.PIPEA1_12l11r_net_1\, 
        \I3.PIPEA1l11r_net_1\, \I3.PIPEA1_308_net_1\, 
        \I3.PIPEA1_12l10r_net_1\, \I3.PIPEA1l10r_net_1\, 
        \I3.PIPEA1_307_net_1\, \I3.PIPEA1_12l9r_net_1\, 
        \I3.PIPEA1l9r_net_1\, \I3.PIPEA1_306_net_1\, 
        \I3.PIPEA1_12l8r_net_1\, \I3.PIPEA1l8r_net_1\, 
        \I3.PIPEA1_305_net_1\, \I3.PIPEA1_12l7r_net_1\, 
        \I3.PIPEA1l7r_net_1\, \I3.PIPEA1_304_net_1\, 
        \I3.PIPEA1_12l6r_net_1\, \I3.PIPEA1l6r_net_1\, 
        \I3.PIPEA1_303_net_1\, \I3.PIPEA1_12l5r_net_1\, 
        \I3.PIPEA1l5r_net_1\, \I3.PIPEA1_302_net_1\, 
        \I3.PIPEA1_12l4r_net_1\, \I3.PIPEA1l4r_net_1\, 
        \I3.PIPEA1_301_net_1\, \I3.PIPEA1_12l3r_net_1\, 
        \I3.PIPEA1l3r_net_1\, \I3.PIPEA1_300_net_1\, 
        \I3.PIPEA1_12l2r_net_1\, \I3.PIPEA1l2r_net_1\, 
        \I3.PIPEA1_299_net_1\, \I3.PIPEA1_12l1r_net_1\, 
        \I3.PIPEA1l1r_net_1\, \I3.PIPEA1_298_net_1\, 
        \I3.PIPEA1_12l0r_net_1\, \I3.PIPEA1l0r_net_1\, 
        \I3.STATE2l4r_net_1\, \I3.REG_1_297_0\, \I3.REG_1_296_0\, 
        \I3.REG_1_295_0\, \I3.REG_1_294_0\, \I3.REG_1_293_0\, 
        \I3.REG_1_292_0\, \I3.REG_1_291_0\, \I3.REG_1_290_0\, 
        \I3.REG_1_284_0\, \I3.REG_1_283_0\, \I3.REG_1_282_0\, 
        \I3.REG_1_281_0\, \I3.N_2297_i\, \I3.REG_1_280_0\, 
        \I3.REG_1_279_0\, \I3.REG_1_278_0\, \I3.REG_1_277_0\, 
        \I3.REG_1_276_0\, \I3.REG_1_275_0\, \I3.REG_1_274_0\, 
        \I3.REG_1_273_0\, \I3.REG_1_272_0\, \I3.N_127\, 
        \I3.REG_1_271_0\, \I3.N_1636\, \I3.REG_1_270_0\, 
        \I3.N_1635\, \I3.N_1673\, \I3.N_98\, \I3.REG_1_269_0\, 
        \I3.N_1634\, \I3.N_1671\, \I3.REG_1_268_0\, \I3.N_1633\, 
        \I3.N_1669\, \I3.REG_1_267_0\, \I3.N_1632\, \I3.N_1667\, 
        \I3.REG_1_266_0\, \I3.N_1631\, \I3.N_1665\, 
        \I3.REG_1_265_0\, \I3.N_1630\, \I3.N_1663\, 
        \I3.REG_1_264_0\, \I3.N_1629\, \I3.N_327\, 
        \I3.REG_1_263_0\, \I3.N_2277_i\, \I3.PIPEA_262_net_1\, 
        \I3.PIPEA_8l31r_net_1\, \I3.N_240\, \I3.PIPEA_261_net_1\, 
        \I3.PIPEA_8l30r_net_1\, \I3.N_239\, \I3.PIPEA_260_net_1\, 
        \I3.PIPEA_8l29r_net_1\, \I3.N_238\, \I3.PIPEA_259_net_1\, 
        \I3.PIPEA_8l28r_net_1\, \I3.N_237\, \I3.PIPEA_258_net_1\, 
        \I3.PIPEA_8l27r_net_1\, \I3.N_236\, \I3.PIPEA_257_net_1\, 
        \I3.PIPEA_8l26r_net_1\, \I3.N_235\, \I3.PIPEA_256_net_1\, 
        \I3.PIPEA_8l25r_net_1\, \I3.N_234\, \I3.PIPEA_255_net_1\, 
        \I3.PIPEA_8l24r_net_1\, \I3.N_233\, \I3.PIPEA_254_net_1\, 
        \I3.PIPEA_8l23r_net_1\, \I3.N_232\, \I3.PIPEA_253_net_1\, 
        \I3.PIPEA_8l22r_net_1\, \I3.N_231\, \I3.PIPEA_252_net_1\, 
        \I3.PIPEA_8l21r_net_1\, \I3.N_230\, \I3.PIPEA_251_net_1\, 
        \I3.PIPEA_8l20r_net_1\, \I3.N_229\, \I3.PIPEA_250_net_1\, 
        \I3.PIPEA_8l19r_net_1\, \I3.N_228\, \I3.PIPEA_249_net_1\, 
        \I3.PIPEA_8l18r_net_1\, \I3.N_227\, \I3.PIPEA_248_net_1\, 
        \I3.PIPEA_8l17r_net_1\, \I3.N_226\, \I3.PIPEA_247_net_1\, 
        \I3.PIPEA_8l16r_net_1\, \I3.N_225\, \I3.PIPEA_246_net_1\, 
        \I3.PIPEA_8l15r_net_1\, \I3.N_224\, \I3.PIPEA_245_net_1\, 
        \I3.PIPEA_8l14r_net_1\, \I3.N_223\, \I3.PIPEA_244_net_1\, 
        \I3.PIPEA_8l13r_net_1\, \I3.N_222\, \I3.PIPEA_243_net_1\, 
        \I3.PIPEA_8l12r_net_1\, \I3.N_221\, \I3.PIPEA_242_net_1\, 
        \I3.PIPEA_8l11r_net_1\, \I3.N_220\, \I3.PIPEA_241_net_1\, 
        \I3.PIPEA_8l10r_net_1\, \I3.N_219\, \I3.PIPEA_240_net_1\, 
        \I3.PIPEA_8l9r_net_1\, \I3.N_218\, \I3.PIPEA_239_net_1\, 
        \I3.PIPEA_8l8r_net_1\, \I3.N_217\, \I3.PIPEA_238_net_1\, 
        \I3.PIPEA_8l7r_net_1\, \I3.N_216\, \I3.PIPEA_237_net_1\, 
        \I3.PIPEA_8l6r_net_1\, \I3.N_215\, \I3.PIPEA_236_net_1\, 
        \I3.PIPEA_8l5r_net_1\, \I3.N_214\, \I3.PIPEA_235_net_1\, 
        \I3.PIPEA_8l4r_net_1\, \I3.N_213\, \I3.PIPEA_234_net_1\, 
        \I3.PIPEA_8l3r_net_1\, \I3.N_212\, \I3.PIPEA_233_net_1\, 
        \I3.PIPEA_8l2r_net_1\, \I3.N_211\, \I3.PIPEA_232_net_1\, 
        \I3.PIPEA_8l1r_net_1\, \I3.N_210\, \I3.PIPEA_231_net_1\, 
        \I3.PIPEA_8l0r_net_1\, \I3.N_209\, \I3.NRDMEBi_230_net_1\, 
        \I3.un1_NRDMEBi_2_sqmuxa_3_net_1\, \I3.EFS_net_1\, 
        \I3.REG1l4r_net_1\, \I3.REG2l4r_net_1\, 
        \I3.REG3l4r_net_1\, \I3.N_297\, \I3.END_PK_229_net_1\, 
        \I3.END_PK_net_1\, \I3.un1_STATE2_11\, 
        \I3.STATE2l3r_net_1\, \I3.un15_anycyc_net_1\, 
        \I3.REG2_228_net_1\, \I3.REG2_15l405r\, \I3.N_1563\, 
        \I3.REG1_227_net_1\, \I3.REG3_226_net_1\, 
        \I3.EVREADi_225_net_1\, \I3.N_1860_2\, 
        \I3.un1_STATE2_9_net_1\, \I3.N_1861\, \I3.REG_1_224_0\, 
        \I3.REG_0_sqmuxa_3\, \I3.REG_1_223_0\, \I3.REG_1_222_0\, 
        \I3.REG_1_221_0\, \I3.REG_1_220_0\, \I3.REG_1_219_0\, 
        \I3.REG_1_218_0\, \I3.REG_1_217_0\, \I3.REG_1_216_0\, 
        \I3.REG_1_215_0\, \I3.REG_1_214_0\, \I3.REG_1_213_0\, 
        \I3.REG_1_212_0\, \I3.REG_1_211_0\, \I3.REG_1_210_0\, 
        \I3.REG_1_209_0\, \I3.REG_1_208_0\, \I3.REG_1_207_0\, 
        \I3.REG_1_206_0\, \I3.REG_1_205_0\, \I3.REG_1_204_0\, 
        \I3.REG_1_203_0\, \I3.REG_1_202_0\, \I3.REG_1_201_0\, 
        \I3.REG_1_200_0\, \I3.REG_1_199_0\, \I3.REG_1_198_0\, 
        \I3.REG_1_197_0\, \I3.REG_1_196_0\, \I3.REG_1_195_0\, 
        \I3.REG_1_194_0\, \I3.REG_1_193_0\, \I3.REG_1_192_0\, 
        \I3.REG_1_191_0\, \I3.REG_1_190_0\, \I3.REG_0_sqmuxa_2\, 
        \I3.REG_1_189_0\, \I3.REG_1_188_0\, \I3.REG_1_187_0\, 
        \I3.REG_1_186_0\, \I3.REG_1_185_0\, \I3.REG_1_184_0\, 
        \I3.REG_1_183_0\, \I3.REG_1_182_0\, \I3.REG_1_181_0\, 
        \I3.REG_1_180_0\, \I3.REG_1_179_0\, \I3.REG_1_178_0\, 
        \I3.REG_1_177_0\, \I3.REG_1_176_0\, \I3.REG_1_175_0\, 
        \I3.REG_1_174_0\, \I3.REG_1_173_0\, \I3.REG_1_172_0\, 
        \I3.REG_1_171_0\, \I3.REG_1_170_0\, \I3.REG_1_169_0\, 
        \I3.REG_1_168_0\, \I3.REG_1_167_0\, \I3.REG_1_166_0\, 
        \I3.REG_1_165_0\, \I3.REG_1_164_0\, \I3.REG_1_163_0\, 
        \I3.REG_1_162_0\, \I3.REG_1_161_0\, \I3.REG_1_160_0\, 
        \I3.REG_1_159_0\, \I3.N_1935\, \I3.REG_1_158_0\, 
        \I3.REG_1_157_0\, \I3.REG_1_156_0\, \I3.REG_1_155_0\, 
        \I3.REG_1_154_0\, \I3.REG_1_153_0\, \I3.REG_1_152_0\, 
        \I3.REG_1_151_0\, \I3.REG_1_150_0\, \I3.REG_1_149_0\, 
        \I3.REG2_148_net_1\, \I3.REG2_147_net_1\, 
        \I3.REG2_146_net_1\, \I3.REG2_145_net_1\, 
        \I3.REG2_144_net_1\, \I3.REG2_143_net_1\, 
        \I3.REG2_142_net_1\, \I3.REG2_141_net_1\, 
        \I3.REG1_140_net_1\, \I3.REG1_139_net_1\, 
        \I3.REG1_138_net_1\, \I3.REG1_137_net_1\, 
        \I3.REG1_136_net_1\, \I3.REG3_0_sqmuxa\, 
        \I3.REG1_135_net_1\, \I3.REG1_134_net_1\, 
        \I3.REG1_133_net_1\, \I3.REG3_132_net_1\, 
        \I3.REG3_131_net_1\, \I3.REG3_130_net_1\, 
        \I3.REG3_129_net_1\, \I3.REG3_128_net_1\, 
        \I3.REG3_127_net_1\, \I3.REG3_126_net_1\, 
        \I3.REG3_125_net_1\, \I3.un1_EVREAD_DS_1_sqmuxa_1_net_1\, 
        \I3.PIPEBl30r_net_1\, \I3.PIPEBl28r_net_1\, 
        \I3.PIPEB_i_0_il31r\, \I3.PIPEBl29r_net_1\, 
        \I3.VDBoff_123_net_1\, \I3.N_81\, \I3.VDBoffal7r_net_1\, 
        \I3.VDBoffbl7r_net_1\, \I3.VDBoff_122_net_1\, \I3.N_79\, 
        \I3.VDBoffal6r_net_1\, \I3.VDBoffbl6r_net_1\, 
        \I3.VDBoff_121_net_1\, \I3.N_77\, \I3.VDBoffal5r_net_1\, 
        \I3.VDBoffbl5r_net_1\, \I3.VDBoff_120_net_1\, \I3.N_2068\, 
        \I3.VDBoffal4r_net_1\, \I3.VDBoffbl4r_net_1\, 
        \I3.VDBoff_119_net_1\, \I3.N_2067\, \I3.VDBoffal3r_net_1\, 
        \I3.VDBoffbl3r_net_1\, \I3.VDBoff_118_net_1\, \I3.N_2066\, 
        \I3.VDBoffal2r_net_1\, \I3.VDBoffbl2r_net_1\, 
        \I3.VDBoff_117_net_1\, \I3.N_2065\, \I3.VDBoffal1r_net_1\, 
        \I3.VDBoffbl1r_net_1\, \I3.VDBoff_116_net_1\, \I3.N_2064\, 
        \I3.VDBoffal0r_net_1\, \I3.VDBoffbl0r_net_1\, \I3.N_1510\, 
        \I3.ASBS_net_1\, \I3.MBLTCYC_114_net_1\, \I3.N_80\, 
        \I3.N_1508\, \I3.N_2055\, \I3.CYCS_net_1\, 
        \I3.ADACKCYC_112_net_1\, \I3.N_1509\, 
        \I3.SELBASE32_net_1\, \I3.NOEDTKi_111_net_1\, 
        \I3.un1_NOEDTKi_0_sqmuxa\, \I3.un1_NOEDTKi_0_sqmuxa_1\, 
        \I3.PURGED_net_1\, \I3.PIPEB_110_net_1\, 
        \I3.PIPEB_109_net_1\, \I3.PIPEB_4l30r_net_1\, 
        \I3.PIPEB_108_net_1\, \I3.PIPEB_4l29r_net_1\, 
        \I3.PIPEB_107_net_1\, \I3.PIPEB_4l28r_net_1\, 
        \I3.PIPEB_106_net_1\, \I3.PIPEBl27r_net_1\, 
        \I3.PIPEB_105_net_1\, \I3.PIPEBl26r_net_1\, 
        \I3.PIPEB_104_net_1\, \I3.PIPEBl25r_net_1\, 
        \I3.PIPEB_103_net_1\, \I3.PIPEBl24r_net_1\, 
        \I3.PIPEB_102_net_1\, \I3.PIPEBl23r_net_1\, 
        \I3.PIPEB_101_net_1\, \I3.PIPEBl22r_net_1\, 
        \I3.PIPEB_100_net_1\, \I3.PIPEBl21r_net_1\, 
        \I3.PIPEB_99_net_1\, \I3.PIPEBl20r_net_1\, 
        \I3.PIPEB_98_net_1\, \I3.PIPEBl19r_net_1\, 
        \I3.PIPEB_97_net_1\, \I3.PIPEBl18r_net_1\, 
        \I3.PIPEB_96_net_1\, \I3.PIPEBl17r_net_1\, 
        \I3.PIPEB_95_net_1\, \I3.PIPEBl16r_net_1\, 
        \I3.PIPEB_94_net_1\, \I3.PIPEBl15r_net_1\, 
        \I3.PIPEB_93_net_1\, \I3.PIPEBl14r_net_1\, 
        \I3.PIPEB_92_net_1\, \I3.PIPEBl13r_net_1\, 
        \I3.PIPEB_91_net_1\, \I3.PIPEBl12r_net_1\, 
        \I3.PIPEB_90_net_1\, \I3.PIPEBl11r_net_1\, 
        \I3.PIPEB_89_net_1\, \I3.PIPEBl10r_net_1\, 
        \I3.PIPEB_88_net_1\, \I3.PIPEBl9r_net_1\, 
        \I3.PIPEB_87_net_1\, \I3.PIPEBl8r_net_1\, 
        \I3.PIPEB_86_net_1\, \I3.PIPEB_85_net_1\, 
        \I3.PIPEBl6r_net_1\, \I3.PIPEB_84_net_1\, 
        \I3.PIPEB_83_net_1\, \I3.PIPEBl4r_net_1\, 
        \I3.PIPEB_82_net_1\, \I3.PIPEBl3r_net_1\, 
        \I3.PIPEB_81_net_1\, \I3.PIPEBl2r_net_1\, 
        \I3.PIPEB_80_net_1\, \I3.PIPEBl1r_net_1\, 
        \I3.PIPEB_79_net_1\, \I3.PIPEBl0r_net_1\, 
        \I3.STBMIC_78_net_1\, \I3.N_1902\, \I3.VAS_77_net_1\, 
        \I3.VAS_i_0_il15r\, \I3.VAS_76_net_1\, \I3.VAS_i_0_il14r\, 
        \I3.VAS_75_net_1\, \I3.VAS_i_0_il13r\, \I3.VAS_74_net_1\, 
        \I3.VASl12r_net_1\, \I3.VAS_73_net_1\, \I3.VASl11r_net_1\, 
        \I3.VAS_72_net_1\, \I3.VAS_i_0_il10r\, \I3.VAS_71_net_1\, 
        \I3.VASl9r_net_1\, \I3.VAS_70_net_1\, \I3.VASl8r_net_1\, 
        \I3.VAS_69_net_1\, \I3.VAS_i_0_il7r\, \I3.VAS_68_net_1\, 
        \I3.VASl6r_net_1\, \I3.VAS_67_net_1\, \I3.VASl5r_net_1\, 
        \I3.VAS_66_net_1\, \I3.VASl4r_net_1\, \I3.VAS_65_net_1\, 
        \I3.VASl3r_net_1\, \I3.VAS_64_net_1\, \I3.VASl2r_net_1\, 
        \I3.VAS_63_net_1\, \I3.VASl1r_net_1\, 
        \I3.MYBERRi_62_net_1\, \I3.un1_MYBERRi_1_sqmuxa\, 
        \I3.LWORDS_61_net_1\, \I3.CYCSF1_60_net_1\, 
        \I3.CYCSF1_net_1\, \I3.VDBoffb_59_net_1\, 
        \I3.VDBoffb_58_net_1\, \I3.VDBoffb_57_net_1\, 
        \I3.VDBoffb_56_net_1\, \I3.VDBoffb_55_net_1\, 
        \I3.VDBoffb_54_net_1\, \I3.VDBoffb_53_net_1\, 
        \I3.VDBoffb_52_net_1\, \I3.VDBoffa_51_net_1\, 
        \I3.VDBoffa_50_net_1\, \I3.VDBoffa_49_net_1\, 
        \I3.VDBoffa_48_net_1\, \I3.VDBoffa_47_net_1\, 
        \I3.VDBoffa_46_net_1\, \I3.VDBoffa_45_net_1\, 
        \I3.VDBoffa_44_net_1\, \I3.PURGED_43_net_1\, 
        \I3.DSSF1_42_net_1\, \I3.N_306\, \I3.N_1512\, 
        \I3.RAMAD_VME_41_net_1\, \I3.RAMAD_VME_40_net_1\, 
        \I3.RAMAD_VME_39_net_1\, \I3.RAMAD_VME_38_net_1\, 
        \I3.RAMAD_VME_37_net_1\, \I3.RAMAD_VME_36_net_1\, 
        \I3.RAMAD_VME_35_net_1\, \I3.RAMAD_VME_34_net_1\, 
        \I3.RAMAD_VME_33_net_1\, \I3.RAMAD_VME_32_net_1\, 
        \I3.TCNT_0_sqmuxa\, \I3.RAMAD_VME_31_net_1\, 
        \I3.RAMAD_VME_30_net_1\, \I3.RAMAD_VME_29_net_1\, 
        \I3.RAMAD_VME_28_net_1\, \I3.RAMAD_VME_27_net_1\, 
        \I3.RAMAD_VME_26_net_1\, \I3.RAMAD_VME_25_net_1\, 
        \I3.RAMAD_VME_24_net_1\, \I3.CYCS1_i_0\, \I3.N_173\, 
        \I3.N_172\, \I3.N_171\, \I3.N_170\, \I3.N_169\, 
        \I3.N_168\, \I3.N_167\, \I3.N_166\, \I3.N_165\, 
        \I3.N_164\, \I3.N_163\, \I3.N_162\, \I3.N_161\, 
        \I3.N_160\, \I3.N_159\, \I3.N_158\, \I3.N_157\, 
        \I3.N_156\, \I3.N_155\, \I3.N_154\, \I3.N_153\, 
        \I3.N_152\, \I3.SINGCYC_net_1\, \I3.N_151\, 
        \I3.BLTCYC_net_1\, \I3.N_150\, \I3.N_148\, \I3.N_146\, 
        \I3.N_145\, \I3.N_144\, \I3.N_143\, \I3.N_142\, 
        \I3.N_1193_ip\, \HWRES_3_adt_net_738__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__net_1\, 
        \I2.DTO_16_1l18r_adt_net_756__net_1\, 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, 
        \I2.N_2826_1_adt_net_794__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__net_1\, 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, 
        \I2.DTO_9_iv_ml28r_adt_net_857__net_1\, 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_888__net_1\, 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_904__net_1\, 
        \I5.REG_2_sqmuxa_0_adt_net_975__net_1\, 
        \I5.N_155_0_adt_net_983__net_1\, 
        \I5.SDAnoe_8_adt_net_991__net_1\, 
        \I2.un1_STATE3_10_1_adt_net_999__net_1\, 
        \I2.N_182_adt_net_1007__net_1\, 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\, 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_1038__net_1\, 
        \I2.N_4667_1_adt_net_1046__net_1\, 
        \I2.N_199_0_adt_net_1054__net_1\, 
        \I2.N_2828_adt_net_1062__net_1\, 
        \I2.STOP_RDSRAM_453_i_adt_net_1077__net_1\, 
        \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_1085__net_1\, 
        \I2.TOKOUT_FL_674_adt_net_1115__net_1\, 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, 
        \I2.N_587_adt_net_1201__net_1\, 
        \I2.N_4547_1_adt_net_1209__net_1\, 
        \I2.N_1170_adt_net_1217__net_1\, 
        \I2.PIPE8_DT_21_i_1l28r_adt_net_1233__net_1\, 
        \I3.N_1463_i_adt_net_1279__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__net_1\, 
        \I3.un1_STATE2_15_1_adt_net_1342__net_1\, 
        \I3.un1_STATE1_13_1_adt_net_1351__net_1\, 
        \I3.un1_STATE2_11_adt_net_1401__net_1\, 
        \I1.N_50_0_adt_net_1409__net_1\, 
        \I3.un1_STATE2_7_1_adt_net_1473__net_1\, 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, 
        \I3.N_1186_adt_net_1488__net_1\, 
        \I3.N_1174_adt_net_1495__net_1\, 
        \I3.N_1180_adt_net_1502__net_1\, 
        \I3.N_1168_adt_net_1509__net_1\, 
        \I3.STATE1_nsl2r_adt_net_1586__net_1\, 
        \I3.VDBi_29l9r_adt_net_1596__net_1\, 
        \I3.VDBi_57l8r_adt_net_1606__net_1\, 
        \I3.VDBi_57l2r_adt_net_1614__net_1\, 
        \I3.VDBi_57l0r_adt_net_1621__net_1\, 
        \I2.N_4646_1_adt_net_1645_Rd1__net_1\, 
        \I2.END_CHAINB1_709_adt_net_2397__net_1\, 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_a5_2_i_adt_net_2404__net_1\, 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\, 
        \I3.VDBi_57l7r_adt_net_3750__net_1\, 
        \I3.VDBi_57l6r_adt_net_3761__net_1\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_4066__net_1\, 
        \I2.N411_adt_net_4092__net_1\, 
        \I3.un1_NOEDTKi_0_sqmuxa_adt_net_4101__net_1\, 
        \I2.N475_adt_net_4127__net_1\, 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_4146__net_1\, 
        \I3.N_290_adt_net_4891_\, 
        \I5.sstate1_ns_el0r_adt_net_8036_\, 
        \I5.sstate2_ns_el1r_adt_net_8563_\, 
        \I5.sstate1_ns_el8r_adt_net_8891_\, 
        \I5.N_75_adt_net_8973_\, 
        \I5.sstate1_ns_el5r_adt_net_9070_\, 
        \I5.sstate1_ns_el1r_adt_net_9243_\, 
        \I5.BITCNTe_adt_net_9456_\, \I5.N_52_adt_net_9528_\, 
        \I5.N_54_adt_net_9598_\, \I5.SDAnoe_8_adt_net_9738_\, 
        \I5.SDAnoe_8_adt_net_9739_\, \I5.N_150_adt_net_9846_\, 
        \I5.N_150_adt_net_9847_\, \I5.SDAout_12_adt_net_9915_\, 
        \I5.SDAout_12_adt_net_9916_\, 
        \I5.SBYTE_9l0r_adt_net_11050_\, 
        \I5.un1_sstate2_3_0_adt_net_11182_\, 
        \I5.REG_1_54_adt_net_11847_\, 
        \I5.DATA_12_ivl1r_adt_net_14302_\, 
        \I4.FLUSH_3_adt_net_15593_\, \I0.CLEAR_adt_net_15816_\, 
        \I0.CLEAR_adt_net_15818_\, \I2.N_3760_adt_net_15910_\, 
        \I2.N_3763_adt_net_16097_\, \I2.N_3764_adt_net_16233_\, 
        \I2.N_4524_adt_net_16803_\, \I2.N_4524_adt_net_16804_\, 
        \I2.FID_7l20r_adt_net_17380_\, 
        \I2.FID_7l20r_adt_net_17388_\, 
        \I2.un1_STATE3_10_1_adt_net_17431__net_1\, 
        \I2.FID_7l19r_adt_net_17517_\, 
        \I2.FID_7l19r_adt_net_17525_\, 
        \I2.FID_7l18r_adt_net_17611_\, 
        \I2.FID_7l18r_adt_net_17619_\, 
        \I2.FID_7l17r_adt_net_17705_\, 
        \I2.FID_7l17r_adt_net_17713_\, 
        \I2.FID_7l16r_adt_net_17799_\, 
        \I2.FID_7l16r_adt_net_17807_\, 
        \I2.FID_7l15r_adt_net_17893_\, 
        \I2.FID_7l15r_adt_net_17901_\, 
        \I2.FID_7l14r_adt_net_17987_\, 
        \I2.FID_7l14r_adt_net_17995_\, 
        \I2.FID_7l13r_adt_net_18081_\, 
        \I2.FID_7l13r_adt_net_18089_\, 
        \I2.FID_7l12r_adt_net_18175_\, 
        \I2.FID_7l12r_adt_net_18183_\, 
        \I2.FID_7l11r_adt_net_18269_\, 
        \I2.FID_7l11r_adt_net_18277_\, 
        \I2.FID_7l10r_adt_net_18363_\, 
        \I2.FID_7l10r_adt_net_18371_\, 
        \I2.FID_7l31r_adt_net_18457_\, 
        \I2.FID_7l31r_adt_net_18465_\, 
        \I2.FID_7l30r_adt_net_18551_\, 
        \I2.FID_7l30r_adt_net_18559_\, 
        \I2.FID_7l29r_adt_net_18645_\, 
        \I2.FID_7l29r_adt_net_18653_\, 
        \I2.FID_7l28r_adt_net_18739_\, 
        \I2.FID_7l28r_adt_net_18747_\, 
        \I2.FID_7l27r_adt_net_18833_\, 
        \I2.FID_7l27r_adt_net_18841_\, 
        \I2.FID_7l26r_adt_net_18927_\, 
        \I2.FID_7l26r_adt_net_18935_\, 
        \I2.FID_7l25r_adt_net_19021_\, 
        \I2.FID_7l25r_adt_net_19029_\, 
        \I2.FID_7l24r_adt_net_19115_\, 
        \I2.FID_7l24r_adt_net_19123_\, 
        \I2.FID_7l23r_adt_net_19209_\, 
        \I2.FID_7l23r_adt_net_19217_\, 
        \I2.FID_7l22r_adt_net_19303_\, 
        \I2.FID_7l22r_adt_net_19311_\, 
        \I2.FID_7l21r_adt_net_19397_\, 
        \I2.FID_7l21r_adt_net_19405_\, 
        \I2.N_4646_1_adt_net_19637_Rd1__net_1\, 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_adt_net_19813_\, 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_19952__net_1\, 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20049__net_1\, 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20059__net_1\, 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20061__net_1\, 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149__net_1\, 
        \I2.N_12169_i_adt_net_20407_\, \I2.N_3902_adt_net_20437_\, 
        \I2.un1_PIPE1_DT_1_sqmuxa_2_adt_net_20482_\, 
        \I2.N_4030_adt_net_20660_\, 
        \I2.SUB9_0_sqmuxa_0_adt_net_20771_\, 
        \I2.N_4273_adt_net_20831_\, \I2.N_4273_adt_net_20928_\, 
        \I2.N_3234_adt_net_21449_\, 
        \I2.STATE2_ns_i_0_1_il0r_adt_net_21493_\, 
        \I2.N_2796_i_0_adt_net_21536_\, 
        \I2.N_2796_i_0_adt_net_21575_\, 
        \I2.un5_tdcgda1_adt_net_21623_\, 
        \I2.un5_tdcgda1_adt_net_21626_\, 
        \I2.N_3887_adt_net_21857_\, \I2.N_3887_adt_net_21862_\, 
        \I2.N_3887_adt_net_21865_\, \I2.N_3347_1_adt_net_21905_\, 
        \I2.N_3214_i_0_adt_net_22011_\, 
        \I2.un1_DTO_cl_1_sqmuxa_2_adt_net_22202_\, 
        \I2.un1_DTO_cl_0_sqmuxa_adt_net_22686_\, 
        \I2.INT_ERRS_adt_net_22801_\, 
        \I2.STATEe_nsl4r_adt_net_22922_\, 
        \I2.STATEe_nsl3r_adt_net_22965_\, 
        \I2.STATEe_nsl3r_adt_net_22967_\, 
        \I2.STATEe_nsl0r_adt_net_23014_\, 
        \I2.N_3457_ip_adt_net_23079_\, 
        \I2.N_3457_ip_adt_net_23080_\, 
        \I2.N_3457_ip_adt_net_23081_\, 
        \I2.STATE1_nsl11r_adt_net_23385_\, 
        \I2.STATE1_nsl11r_adt_net_23387_\, 
        \I2.STATE1_nsl6r_adt_net_23511_\, 
        \I2.N_3012_adt_net_24321_\, \I2.N_3012_adt_net_24327_\, 
        \I2.N_12254_i_adt_net_24491_\, 
        \I2.STATE3_nsl8r_adt_net_24815_\, 
        \I2.STATE3_nsl6r_adt_net_24857_\, 
        \I2.STATE2_nsl2r_adt_net_24907_\, 
        \I2.STATE2_nsl2r_adt_net_24911_\, 
        \I2.STATE2_nsl2r_adt_net_24916_\, 
        \I2.STATE2_nsl1r_adt_net_24963_\, 
        \I2.STATE2_nsl1r_adt_net_24965_\, 
        \I2.N_3267_adt_net_25763_\, \I2.N_4344_adt_net_26298_\, 
        \I2.G_EVNT_NUM_n11_adt_net_26872_\, 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26950_\, 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26951_\, 
        \I2.L2SERVe_adt_net_26991_\, 
        \I2.ROFFSETe_0_adt_net_27175__net_1\, 
        \I2.ROFFSETe_0_adt_net_27185__net_1\, 
        \I2.ROFFSETe_0_adt_net_27187__net_1\, 
        \I2.DTO_9l31r_adt_net_27894_\, 
        \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_28030__net_1\, 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_28083__net_1\, 
        \I2.DTO_16_1l31r_adt_net_28246_\, 
        \I2.DTO_16_1l31r_adt_net_28248_\, 
        \I2.DTO_16_1l31r_adt_net_28255_\, 
        \I2.DTO_16_1l31r_adt_net_28256_\, 
        \I2.DTO_16_1_iv_1l30r_adt_net_28466_\, 
        \I2.DTO_16_1_iv_1l30r_adt_net_28472_\, 
        \I2.N_4159_adt_net_28676_\, 
        \I2.DTO_16_1l29r_adt_net_28730_\, 
        \I2.DTO_16_1l29r_adt_net_28732_\, 
        \I2.DTO_16_1l29r_adt_net_28739_\, 
        \I2.DTO_16_1l29r_adt_net_28740_\, 
        \I2.DTO_9_iv_ml28r_adt_net_28906__net_1\, 
        \I2.DTO_16_1_iv_0l28r_adt_net_28950_\, 
        \I2.DTO_16_1_ivl28r_adt_net_28982_\, 
        \I2.N_4647_adt_net_29104_\, 
        \I2.DTO_16_1l27r_adt_net_29240_\, 
        \I2.DTO_16_1l27r_adt_net_29242_\, 
        \I2.DTO_16_1l27r_adt_net_29251_\, 
        \I2.DTO_16_1l27r_adt_net_29252_\, 
        \I2.DTO_16_1l26r_adt_net_29426_\, 
        \I2.DTO_16_1l26r_adt_net_29428_\, 
        \I2.DTO_16_1l26r_adt_net_29437_\, 
        \I2.DTO_16_1l26r_adt_net_29438_\, 
        \I2.DTO_16_1l25r_adt_net_29612_\, 
        \I2.DTO_16_1l25r_adt_net_29614_\, 
        \I2.DTO_16_1l25r_adt_net_29623_\, 
        \I2.DTO_16_1l25r_adt_net_29624_\, 
        \I2.DTO_9l24r_adt_net_29794_\, 
        \I2.DTO_9l24r_adt_net_29802_\, 
        \I2.DTO_16_1l24r_adt_net_29854_\, 
        \I2.DTO_16_1l24r_adt_net_29860_\, 
        \I2.DTO_16_1l24r_adt_net_29868_\, 
        \I2.DTO_16_1l24r_adt_net_29869_\, 
        \I2.DTO_16_1l24r_adt_net_29870_\, 
        \I2.DTO_9l23r_adt_net_30040_\, 
        \I2.DTO_9l23r_adt_net_30048_\, 
        \I2.DTO_16_1l23r_adt_net_30100_\, 
        \I2.DTO_16_1l23r_adt_net_30106_\, 
        \I2.DTO_16_1l23r_adt_net_30114_\, 
        \I2.DTO_16_1l23r_adt_net_30115_\, 
        \I2.DTO_16_1l23r_adt_net_30116_\, 
        \I2.DTO_9l22r_adt_net_30286_\, 
        \I2.DTO_9l22r_adt_net_30294_\, 
        \I2.DTO_16_1l22r_adt_net_30346_\, 
        \I2.DTO_16_1l22r_adt_net_30352_\, 
        \I2.DTO_16_1l22r_adt_net_30360_\, 
        \I2.DTO_16_1l22r_adt_net_30361_\, 
        \I2.DTO_16_1l22r_adt_net_30362_\, 
        \I2.DTO_16_1l21r_adt_net_30536_\, 
        \I2.DTO_16_1l21r_adt_net_30538_\, 
        \I2.DTO_16_1l21r_adt_net_30547_\, 
        \I2.DTO_16_1l21r_adt_net_30548_\, 
        \I2.DTO_9l20r_adt_net_30718_\, 
        \I2.DTO_9l20r_adt_net_30726_\, 
        \I2.DTO_16_1l20r_adt_net_30778_\, 
        \I2.DTO_16_1l20r_adt_net_30786_\, 
        \I2.DTO_16_1l20r_adt_net_30792_\, 
        \I2.DTO_16_1l20r_adt_net_30793_\, 
        \I2.DTO_16_1l20r_adt_net_30794_\, 
        \I2.DTO_16_1l19r_adt_net_30968_\, 
        \I2.DTO_16_1l19r_adt_net_30970_\, 
        \I2.DTO_16_1l19r_adt_net_30979_\, 
        \I2.DTO_16_1l19r_adt_net_30980_\, 
        \I2.DTO_16_1l18r_adt_net_31333_\, 
        \I2.DTO_16_1l18r_adt_net_31339_\, 
        \I2.DTO_16_1l18r_adt_net_31345_\, 
        \I2.DTO_16_1l18r_adt_net_31346_\, 
        \I2.DTO_16_1l17r_adt_net_31520_\, 
        \I2.DTO_16_1l17r_adt_net_31522_\, 
        \I2.DTO_16_1l17r_adt_net_31531_\, 
        \I2.DTO_16_1l17r_adt_net_31532_\, 
        \I2.DTO_16_1l16r_adt_net_31706_\, 
        \I2.DTO_16_1l16r_adt_net_31708_\, 
        \I2.DTO_16_1l16r_adt_net_31717_\, 
        \I2.DTO_16_1l16r_adt_net_31718_\, 
        \I2.DTO_9l15r_adt_net_31888_\, 
        \I2.DTO_9l15r_adt_net_31896_\, 
        \I2.DTO_16_1l15r_adt_net_31948_\, 
        \I2.DTO_16_1l15r_adt_net_31956_\, 
        \I2.DTO_16_1l15r_adt_net_31962_\, 
        \I2.DTO_16_1l15r_adt_net_31963_\, 
        \I2.DTO_16_1l15r_adt_net_31964_\, 
        \I2.DTO_9l14r_adt_net_32134_\, 
        \I2.DTO_9l14r_adt_net_32142_\, 
        \I2.DTO_16_1l14r_adt_net_32194_\, 
        \I2.DTO_16_1l14r_adt_net_32202_\, 
        \I2.DTO_16_1l14r_adt_net_32208_\, 
        \I2.DTO_16_1l14r_adt_net_32209_\, 
        \I2.DTO_16_1l14r_adt_net_32210_\, 
        \I2.DTO_16_1l13r_adt_net_32384_\, 
        \I2.DTO_16_1l13r_adt_net_32386_\, 
        \I2.DTO_16_1l13r_adt_net_32395_\, 
        \I2.DTO_16_1l13r_adt_net_32396_\, 
        \I2.N_3966_adt_net_32562_\, 
        \I2.DTO_16_1l12r_adt_net_32622_\, 
        \I2.DTO_16_1l12r_adt_net_32624_\, 
        \I2.DTO_16_1l12r_adt_net_32632_\, 
        \I2.DTO_16_1l12r_adt_net_32633_\, 
        \I2.DTO_16_1l12r_adt_net_32634_\, 
        \I2.DTO_9l11r_adt_net_32804_\, 
        \I2.DTO_9l11r_adt_net_32812_\, 
        \I2.DTO_16_1l11r_adt_net_32864_\, 
        \I2.DTO_16_1l11r_adt_net_32872_\, 
        \I2.DTO_16_1l11r_adt_net_32878_\, 
        \I2.DTO_16_1l11r_adt_net_32879_\, 
        \I2.DTO_16_1l11r_adt_net_32880_\, 
        \I2.DTO_16_1l10r_adt_net_33054_\, 
        \I2.DTO_16_1l10r_adt_net_33056_\, 
        \I2.DTO_16_1l10r_adt_net_33065_\, 
        \I2.DTO_16_1l10r_adt_net_33066_\, 
        \I2.DTO_16_1l9r_adt_net_33240_\, 
        \I2.DTO_16_1l9r_adt_net_33242_\, 
        \I2.DTO_16_1l9r_adt_net_33251_\, 
        \I2.DTO_16_1l9r_adt_net_33252_\, 
        \I2.N_3967_adt_net_33418_\, 
        \I2.DTO_16_1l8r_adt_net_33478_\, 
        \I2.DTO_16_1l8r_adt_net_33480_\, 
        \I2.DTO_16_1l8r_adt_net_33488_\, 
        \I2.DTO_16_1l8r_adt_net_33489_\, 
        \I2.DTO_16_1l8r_adt_net_33490_\, 
        \I2.DTO_9l7r_adt_net_33660_\, 
        \I2.DTO_9l7r_adt_net_33668_\, 
        \I2.DTO_16_1l7r_adt_net_33720_\, 
        \I2.DTO_16_1l7r_adt_net_33728_\, 
        \I2.DTO_16_1l7r_adt_net_33734_\, 
        \I2.DTO_16_1l7r_adt_net_33735_\, 
        \I2.DTO_16_1l7r_adt_net_33736_\, 
        \I2.DTO_16_1l6r_adt_net_33910_\, 
        \I2.DTO_16_1l6r_adt_net_33912_\, 
        \I2.DTO_16_1l6r_adt_net_33921_\, 
        \I2.DTO_16_1l6r_adt_net_33922_\, 
        \I2.DTO_16_1l5r_adt_net_34192_\, 
        \I2.DTO_16_1l5r_adt_net_34198_\, 
        \I2.DTO_16_1l5r_adt_net_34199_\, 
        \I2.DTO_16_1l5r_adt_net_34200_\, 
        \I2.DTO_16_1l4r_adt_net_34374_\, 
        \I2.DTO_16_1l4r_adt_net_34376_\, 
        \I2.DTO_16_1l4r_adt_net_34385_\, 
        \I2.DTO_16_1l4r_adt_net_34386_\, 
        \I2.DTO_9_ivl3r_adt_net_34552_\, 
        \I2.DTO_16_1_iv_1l3r_adt_net_34602_\, 
        \I2.DTO_16_1_iv_1l3r_adt_net_34608_\, 
        \I2.DTO_9_ivl2r_adt_net_34812_\, 
        \I2.DTO_16_1_iv_0_1l2r_adt_net_34862_\, 
        \I2.DTO_16_1_iv_0_1l2r_adt_net_34868_\, 
        \I2.DTO_9_ivl1r_adt_net_35072_\, 
        \I2.DTO_16_1_iv_1l1r_adt_net_35122_\, 
        \I2.DTO_16_1_iv_1l1r_adt_net_35128_\, 
        \I2.DTO_9_ivl0r_adt_net_35332_\, 
        \I2.DTO_16_1_iv_0_0_1l0r_adt_net_35382_\, 
        \I2.DTO_16_1_iv_0_0_1l0r_adt_net_35388_\, 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35702__net_1\, 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35789__net_1\, 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35891_\, 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35893_\, 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35897_\, 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35904_\, 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35905_\, 
        \I2.DTE_21_1l17r_adt_net_36140_\, 
        \I2.DTE_21_1l17r_adt_net_36142_\, 
        \I2.DTE_21_1l17r_adt_net_36146_\, 
        \I2.DTE_21_1l17r_adt_net_36153_\, 
        \I2.DTE_21_1l17r_adt_net_36154_\, 
        \I2.DTE_21_1l31r_adt_net_36411_\, 
        \I2.DTE_21_1l31r_adt_net_36416_\, 
        \I2.DTE_21_1l31r_adt_net_36417_\, 
        \I2.DTE_21_1_0_iv_1l30r_adt_net_36505_\, 
        \I2.DTE_21_1_0_iv_1l30r_adt_net_36511_\, 
        \I2.DTE_21_1l29r_adt_net_36645_\, 
        \I2.DTE_21_1l29r_adt_net_36650_\, 
        \I2.DTE_21_1l29r_adt_net_36651_\, 
        \I2.DTE_21_1l28r_adt_net_36757_\, 
        \I2.DTE_21_1l28r_adt_net_36758_\, 
        \I2.DTE_21_1l28r_adt_net_36759_\, 
        \I2.DTE_21_1l27r_adt_net_36849_\, 
        \I2.DTE_21_1l27r_adt_net_36860_\, 
        \I2.DTE_21_1l27r_adt_net_36861_\, 
        \I2.DTE_21_1l26r_adt_net_36951_\, 
        \I2.DTE_21_1l26r_adt_net_36962_\, 
        \I2.DTE_21_1l26r_adt_net_36963_\, 
        \I2.N_4644_adt_net_37053_\, \I2.N_4644_adt_net_37064_\, 
        \I2.N_4644_adt_net_37065_\, 
        \I2.DTE_21_1l24r_adt_net_37173_\, 
        \I2.DTE_21_1l24r_adt_net_37174_\, 
        \I2.DTE_21_1l23r_adt_net_37283_\, 
        \I2.DTE_21_1l23r_adt_net_37284_\, 
        \I2.DTE_21_1l22r_adt_net_37393_\, 
        \I2.DTE_21_1l22r_adt_net_37394_\, 
        \I2.DTE_21_1l21r_adt_net_37485_\, 
        \I2.DTE_21_1l21r_adt_net_37496_\, 
        \I2.DTE_21_1l21r_adt_net_37497_\, 
        \I2.DTE_21_1l20r_adt_net_37603_\, 
        \I2.DTE_21_1l20r_adt_net_37605_\, 
        \I2.DTE_21_1l20r_adt_net_37612_\, 
        \I2.DTE_21_1l20r_adt_net_37614_\, 
        \I2.DTE_21_1l20r_adt_net_37615_\, 
        \I2.DTE_21_1l19r_adt_net_37713_\, 
        \I2.DTE_21_1l19r_adt_net_37715_\, 
        \I2.DTE_21_1l19r_adt_net_37723_\, 
        \I2.DTE_21_1l19r_adt_net_37724_\, 
        \I2.DTE_21_1l16r_adt_net_37823_\, 
        \I2.DTE_21_1l16r_adt_net_37825_\, 
        \I2.DTE_21_1l16r_adt_net_37833_\, 
        \I2.DTE_21_1l16r_adt_net_37834_\, 
        \I2.DTE_21_1l15r_adt_net_37943_\, 
        \I2.DTE_21_1l15r_adt_net_37950_\, 
        \I2.DTE_21_1l15r_adt_net_37952_\, 
        \I2.DTE_21_1l15r_adt_net_37953_\, 
        \I2.DTE_21_1l14r_adt_net_38061_\, 
        \I2.DTE_21_1l14r_adt_net_38068_\, 
        \I2.DTE_21_1l14r_adt_net_38070_\, 
        \I2.DTE_21_1l14r_adt_net_38071_\, 
        \I2.DTE_21_1l13r_adt_net_38169_\, 
        \I2.DTE_21_1l13r_adt_net_38171_\, 
        \I2.DTE_21_1l13r_adt_net_38179_\, 
        \I2.DTE_21_1l13r_adt_net_38180_\, 
        \I2.DTE_21_1l12r_adt_net_38279_\, 
        \I2.DTE_21_1l12r_adt_net_38283_\, 
        \I2.DTE_21_1l12r_adt_net_38296_\, 
        \I2.DTE_21_1l12r_adt_net_38297_\, 
        \I2.DTE_21_1l12r_adt_net_38298_\, 
        \I2.DTE_21_1l11r_adt_net_38407_\, 
        \I2.DTE_21_1l11r_adt_net_38414_\, 
        \I2.DTE_21_1l11r_adt_net_38416_\, 
        \I2.DTE_21_1l11r_adt_net_38417_\, 
        \I2.DTE_21_1l10r_adt_net_38515_\, 
        \I2.DTE_21_1l10r_adt_net_38517_\, 
        \I2.DTE_21_1l10r_adt_net_38525_\, 
        \I2.DTE_21_1l10r_adt_net_38526_\, 
        \I2.DTE_21_1l9r_adt_net_38625_\, 
        \I2.DTE_21_1l9r_adt_net_38627_\, 
        \I2.DTE_21_1l9r_adt_net_38635_\, 
        \I2.DTE_21_1l9r_adt_net_38636_\, 
        \I2.DTE_21_1l8r_adt_net_38735_\, 
        \I2.DTE_21_1l8r_adt_net_38739_\, 
        \I2.DTE_21_1l8r_adt_net_38752_\, 
        \I2.DTE_21_1l8r_adt_net_38753_\, 
        \I2.DTE_21_1l8r_adt_net_38754_\, 
        \I2.DTE_21_1l7r_adt_net_38863_\, 
        \I2.DTE_21_1l7r_adt_net_38870_\, 
        \I2.DTE_21_1l7r_adt_net_38872_\, 
        \I2.DTE_21_1l7r_adt_net_38873_\, 
        \I2.DTE_21_1l6r_adt_net_38971_\, 
        \I2.DTE_21_1l6r_adt_net_38973_\, 
        \I2.DTE_21_1l6r_adt_net_38981_\, 
        \I2.DTE_21_1l6r_adt_net_38982_\, 
        \I2.DTE_21_1l5r_adt_net_39091_\, 
        \I2.DTE_21_1l5r_adt_net_39098_\, 
        \I2.DTE_21_1l5r_adt_net_39100_\, 
        \I2.DTE_21_1l5r_adt_net_39101_\, 
        \I2.DTE_21_1l4r_adt_net_39199_\, 
        \I2.DTE_21_1l4r_adt_net_39201_\, 
        \I2.DTE_21_1l4r_adt_net_39209_\, 
        \I2.DTE_21_1l4r_adt_net_39210_\, 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39303_\, 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39312_\, 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39313_\, 
        \I2.DTE_21_1_iv_2_il2r_adt_net_39443_\, 
        \I2.DTE_21_1_iv_2_il2r_adt_net_39452_\, 
        \I2.DTE_21_1_iv_2_il2r_adt_net_39453_\, 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39583_\, 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39592_\, 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39593_\, 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39723_\, 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39732_\, 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39733_\, 
        \I2.N_4262_adt_net_39852_\, 
        \I2.N_2828_adt_net_39955__net_1\, 
        \I2.N_2828_adt_net_39957__net_1\, 
        \I2.N_2826_1_adt_net_40738__net_1\, 
        \I2.N_2826_1_adt_net_40744__net_1\, 
        \I2.N_230_i_i_adt_net_41076_\, \I2.N_3926_adt_net_42578_\, 
        \I2.N_3920_adt_net_43068_\, 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_44987__net_1\, 
        \I2.PIPE1_DT_42l31r_adt_net_45035_\, 
        \I2.PIPE1_DT_42l31r_adt_net_45041_\, 
        \I2.un1_STATE1_40_1_adt_net_45381__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45387__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45389__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45408__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45409__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45410__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45413__net_1\, 
        \I2.PIPE1_DT_42l30r_adt_net_45594_\, 
        \I2.PIPE1_DT_42l30r_adt_net_45595_\, 
        \I2.PIPE1_DT_42l29r_adt_net_45835_\, 
        \I2.PIPE1_DT_42l29r_adt_net_45836_\, 
        \I2.PIPE1_DT_42l29r_adt_net_45837_\, 
        \I2.PIPE1_DT_42l29r_adt_net_45838_\, 
        \I2.PIPE1_DT_42l29r_adt_net_45839_\, 
        \I2.PIPE1_DT_42l28r_adt_net_45929_\, 
        \I2.PIPE1_DT_42l28r_adt_net_45931_\, 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46027_\, 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46033_\, 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46038_\, 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46039_\, 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46167_\, 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46173_\, 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46178_\, 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46179_\, 
        \I2.PIPE1_DT_42_1_iv_1_il25r_adt_net_46307_\, 
        \I2.PIPE1_DT_42_1_iv_1_il25r_adt_net_46311_\, 
        \I2.PIPE1_DT_42_1_iv_1_il24r_adt_net_46469_\, 
        \I2.PIPE1_DT_42_1_iv_0_il24r_adt_net_46513_\, 
        \I2.PIPE1_DT_42l23r_adt_net_46639_\, 
        \I2.PIPE1_DT_42l23r_adt_net_46641_\, 
        \I2.PIPE1_DT_42l23r_adt_net_46647_\, 
        \I2.PIPE1_DT_42l23r_adt_net_46653_\, 
        \I2.PIPE1_DT_42l23r_adt_net_46654_\, 
        \I2.PIPE1_DT_42l22r_adt_net_46749_\, 
        \I2.PIPE1_DT_42l22r_adt_net_46751_\, 
        \I2.PIPE1_DT_42l22r_adt_net_46757_\, 
        \I2.PIPE1_DT_42l22r_adt_net_46763_\, 
        \I2.PIPE1_DT_42l22r_adt_net_46764_\, 
        \I2.PIPE1_DT_42l21r_adt_net_46859_\, 
        \I2.PIPE1_DT_42l21r_adt_net_46861_\, 
        \I2.PIPE1_DT_42l21r_adt_net_46867_\, 
        \I2.PIPE1_DT_42l21r_adt_net_46873_\, 
        \I2.PIPE1_DT_42l21r_adt_net_46874_\, 
        \I2.PIPE1_DT_42l20r_adt_net_47053_\, 
        \I2.PIPE1_DT_42l20r_adt_net_47055_\, 
        \I2.PIPE1_DT_42l20r_adt_net_47061_\, 
        \I2.PIPE1_DT_42l20r_adt_net_47067_\, 
        \I2.PIPE1_DT_42l20r_adt_net_47068_\, 
        \I2.PIPE1_DT_42l19r_adt_net_47247_\, 
        \I2.PIPE1_DT_42l19r_adt_net_47249_\, 
        \I2.PIPE1_DT_42l19r_adt_net_47255_\, 
        \I2.PIPE1_DT_42l19r_adt_net_47261_\, 
        \I2.PIPE1_DT_42l19r_adt_net_47262_\, 
        \I2.PIPE1_DT_42l18r_adt_net_47441_\, 
        \I2.PIPE1_DT_42l18r_adt_net_47443_\, 
        \I2.PIPE1_DT_42l18r_adt_net_47449_\, 
        \I2.PIPE1_DT_42l18r_adt_net_47455_\, 
        \I2.PIPE1_DT_42l18r_adt_net_47456_\, 
        \I2.PIPE1_DT_42l17r_adt_net_47635_\, 
        \I2.PIPE1_DT_42l17r_adt_net_47637_\, 
        \I2.PIPE1_DT_42l17r_adt_net_47643_\, 
        \I2.PIPE1_DT_42l17r_adt_net_47649_\, 
        \I2.PIPE1_DT_42l17r_adt_net_47650_\, 
        \I2.PIPE1_DT_42l16r_adt_net_47833_\, 
        \I2.PIPE1_DT_42l16r_adt_net_47835_\, 
        \I2.PIPE1_DT_42l16r_adt_net_47837_\, 
        \I2.PIPE1_DT_42l16r_adt_net_47850_\, 
        \I2.PIPE1_DT_42l16r_adt_net_47851_\, 
        \I2.PIPE1_DT_42l16r_adt_net_47852_\, 
        \I2.N_13_adt_net_47925_\, 
        \I2.BNCID_VECTror_8_tz_0_i_adt_net_48007_\, 
        \I2.BNCID_VECTror_8_tz_i_adt_net_48039_\, 
        \I2.BNCID_VECTror_9_tz_adt_net_48087_\, 
        \I2.BNCID_VECTror_9_tz_adt_net_48091_\, 
        \I2.BNCID_VECTror_9_tz_adt_net_48098_\, 
        \I2.BNCID_VECTror_9_tz_adt_net_48099_\, 
        \I2.BNCID_VECTror_10_tz_0_adt_net_48139_\, 
        \I2.BNCID_VECTror_10_tz_adt_net_48171_\, 
        \I2.BNCID_VECTror_adt_net_48219__net_1\, 
        \I2.BNCID_VECTror_adt_net_48223__net_1\, 
        \I2.BNCID_VECTror_adt_net_48230__net_1\, 
        \I2.BNCID_VECTror_adt_net_48231__net_1\, 
        \I2.BNCID_VECTror_adt_net_48326_\, 
        \I2.BNCID_VECTror_adt_net_48365_\, 
        \I2.BNCID_VECTror_adt_net_48367_\, 
        \I2.BNCID_VECTror_adt_net_48422_\, 
        \I2.BNCID_VECTror_adt_net_48461_\, 
        \I2.BNCID_VECTror_adt_net_48463_\, 
        \I2.N_3238_adt_net_48555_\, 
        \I2.PIPE1_DT_42l15r_adt_net_48697_\, 
        \I2.PIPE1_DT_42l15r_adt_net_48701_\, 
        \I2.PIPE1_DT_42l15r_adt_net_48707_\, 
        \I2.PIPE1_DT_42l15r_adt_net_48714_\, 
        \I2.PIPE1_DT_42l15r_adt_net_48715_\, 
        \I2.PIPE1_DT_42l15r_adt_net_48716_\, 
        \I2.PIPE1_DT_42l15r_adt_net_48717_\, 
        \I2.PIPE1_DT_42l14r_adt_net_48944_\, 
        \I2.PIPE1_DT_42l14r_adt_net_48948_\, 
        \I2.PIPE1_DT_42l14r_adt_net_48954_\, 
        \I2.PIPE1_DT_42l14r_adt_net_48962_\, 
        \I2.PIPE1_DT_42l14r_adt_net_48963_\, 
        \I2.PIPE1_DT_42l14r_adt_net_48964_\, 
        \I2.PIPE1_DT_42l13r_adt_net_49191_\, 
        \I2.PIPE1_DT_42l13r_adt_net_49195_\, 
        \I2.PIPE1_DT_42l13r_adt_net_49201_\, 
        \I2.PIPE1_DT_42l13r_adt_net_49209_\, 
        \I2.PIPE1_DT_42l13r_adt_net_49210_\, 
        \I2.PIPE1_DT_42l13r_adt_net_49211_\, 
        \I2.PIPE1_DT_42l12r_adt_net_49438_\, 
        \I2.PIPE1_DT_42l12r_adt_net_49442_\, 
        \I2.PIPE1_DT_42l12r_adt_net_49448_\, 
        \I2.PIPE1_DT_42l12r_adt_net_49456_\, 
        \I2.PIPE1_DT_42l12r_adt_net_49457_\, 
        \I2.PIPE1_DT_42l12r_adt_net_49458_\, 
        \I2.PIPE1_DT_42l11r_adt_net_49685_\, 
        \I2.PIPE1_DT_42l11r_adt_net_49689_\, 
        \I2.PIPE1_DT_42l11r_adt_net_49695_\, 
        \I2.PIPE1_DT_42l11r_adt_net_49703_\, 
        \I2.PIPE1_DT_42l11r_adt_net_49704_\, 
        \I2.PIPE1_DT_42l11r_adt_net_49705_\, 
        \I2.PIPE1_DT_42l10r_adt_net_49932_\, 
        \I2.PIPE1_DT_42l10r_adt_net_49936_\, 
        \I2.PIPE1_DT_42l10r_adt_net_49942_\, 
        \I2.PIPE1_DT_42l10r_adt_net_49950_\, 
        \I2.PIPE1_DT_42l10r_adt_net_49951_\, 
        \I2.PIPE1_DT_42l10r_adt_net_49952_\, 
        \I2.PIPE1_DT_42l9r_adt_net_50179_\, 
        \I2.PIPE1_DT_42l9r_adt_net_50183_\, 
        \I2.PIPE1_DT_42l9r_adt_net_50189_\, 
        \I2.PIPE1_DT_42l9r_adt_net_50197_\, 
        \I2.PIPE1_DT_42l9r_adt_net_50198_\, 
        \I2.PIPE1_DT_42l9r_adt_net_50199_\, 
        \I2.PIPE1_DT_42l8r_adt_net_50426_\, 
        \I2.PIPE1_DT_42l8r_adt_net_50430_\, 
        \I2.PIPE1_DT_42l8r_adt_net_50436_\, 
        \I2.PIPE1_DT_42l8r_adt_net_50444_\, 
        \I2.PIPE1_DT_42l8r_adt_net_50445_\, 
        \I2.PIPE1_DT_42l8r_adt_net_50446_\, 
        \I2.PIPE1_DT_42l7r_adt_net_50673_\, 
        \I2.PIPE1_DT_42l7r_adt_net_50677_\, 
        \I2.PIPE1_DT_42l7r_adt_net_50683_\, 
        \I2.PIPE1_DT_42l7r_adt_net_50691_\, 
        \I2.PIPE1_DT_42l7r_adt_net_50692_\, 
        \I2.PIPE1_DT_42l7r_adt_net_50693_\, 
        \I2.PIPE1_DT_42l6r_adt_net_50920_\, 
        \I2.PIPE1_DT_42l6r_adt_net_50924_\, 
        \I2.PIPE1_DT_42l6r_adt_net_50930_\, 
        \I2.PIPE1_DT_42l6r_adt_net_50938_\, 
        \I2.PIPE1_DT_42l6r_adt_net_50939_\, 
        \I2.PIPE1_DT_42l6r_adt_net_50940_\, 
        \I2.PIPE1_DT_42l5r_adt_net_51167_\, 
        \I2.PIPE1_DT_42l5r_adt_net_51171_\, 
        \I2.PIPE1_DT_42l5r_adt_net_51177_\, 
        \I2.PIPE1_DT_42l5r_adt_net_51185_\, 
        \I2.PIPE1_DT_42l5r_adt_net_51186_\, 
        \I2.PIPE1_DT_42l5r_adt_net_51187_\, 
        \I2.PIPE1_DT_42l4r_adt_net_51414_\, 
        \I2.PIPE1_DT_42l4r_adt_net_51418_\, 
        \I2.PIPE1_DT_42l4r_adt_net_51424_\, 
        \I2.PIPE1_DT_42l4r_adt_net_51432_\, 
        \I2.PIPE1_DT_42l4r_adt_net_51433_\, 
        \I2.PIPE1_DT_42l4r_adt_net_51434_\, 
        \I2.PIPE1_DT_42l3r_adt_net_51617_\, 
        \I2.PIPE1_DT_42l3r_adt_net_51627_\, 
        \I2.PIPE1_DT_42l3r_adt_net_51634_\, 
        \I2.PIPE1_DT_42l3r_adt_net_51635_\, 
        \I2.PIPE1_DT_42l3r_adt_net_51636_\, 
        \I2.PIPE1_DT_42l3r_adt_net_51637_\, 
        \I2.PIPE1_DT_42l2r_adt_net_51819_\, 
        \I2.PIPE1_DT_42l2r_adt_net_51829_\, 
        \I2.PIPE1_DT_42l2r_adt_net_51836_\, 
        \I2.PIPE1_DT_42l2r_adt_net_51837_\, 
        \I2.PIPE1_DT_42l2r_adt_net_51838_\, 
        \I2.PIPE1_DT_42l2r_adt_net_51839_\, 
        \I2.PIPE1_DT_42l1r_adt_net_52027_\, 
        \I2.PIPE1_DT_42l1r_adt_net_52031_\, 
        \I2.PIPE1_DT_42l1r_adt_net_52043_\, 
        \I2.PIPE1_DT_42l1r_adt_net_52044_\, 
        \I2.PIPE1_DT_42l1r_adt_net_52045_\, 
        \I2.PIPE1_DT_42l1r_adt_net_52046_\, 
        \I2.PIPE1_DT_42l0r_adt_net_52231_\, 
        \I2.PIPE1_DT_42l0r_adt_net_52239_\, 
        \I2.PIPE1_DT_42l0r_adt_net_52246_\, 
        \I2.PIPE1_DT_42l0r_adt_net_52247_\, 
        \I2.PIPE1_DT_42l0r_adt_net_52248_\, 
        \I2.PIPE1_DT_42l0r_adt_net_52249_\, 
        \I2.N_3292_adt_net_52393_\, 
        \I2.un1_STATE1_39_6_i_adt_net_52471_\, 
        \I2.un1_STATE1_39_6_i_adt_net_52472_\, 
        \I2.un1_STATE1_39_6_i_adt_net_52473_\, 
        \I2.un1_STATE1_38_adt_net_52557_\, 
        \I2.un1_STATE1_38_adt_net_52564_\, 
        \I2.EVNT_WORD_713_adt_net_53148_\, 
        \I2.un1_STATE2_7_adt_net_53240_\, 
        \I2.N_3281_adt_net_53327_\, 
        \I2.END_CHAINB1_709_adt_net_53455_\, 
        \I2.END_CHAINB1_709_adt_net_53463_\, 
        \I2.END_CHAINA1_708_adt_net_53509_\, 
        \I2.END_CHAINA1_708_adt_net_53513_\, 
        \I2.FIRST_TDC_675_adt_net_61236_\, 
        \I2.TOKOUT_FL_674_adt_net_61290__net_1\, 
        \I2.TOKOUT_FL_674_adt_net_61319_\, 
        \I2.N_3866_adt_net_61369_\, \I2.N_4528_adt_net_63525_\, 
        \I2.N_4527_adt_net_63801_\, 
        \I2.LEAD_FLAG6_644_adt_net_63844_\, 
        \I2.N_4529_adt_net_63916_\, 
        \I2.LEAD_FLAG6_643_adt_net_63956_\, 
        \I2.N_4530_adt_net_64028_\, 
        \I2.LEAD_FLAG6_642_adt_net_64068_\, 
        \I2.N_4531_adt_net_64140_\, 
        \I2.LEAD_FLAG6_641_adt_net_64180_\, 
        \I2.N_4532_adt_net_64252_\, 
        \I2.LEAD_FLAG6_640_adt_net_64292_\, 
        \I2.N_4533_adt_net_64364_\, 
        \I2.LEAD_FLAG6_639_adt_net_64404_\, 
        \I2.N_4534_adt_net_64476_\, 
        \I2.LEAD_FLAG6_638_adt_net_64516_\, 
        \I2.N_4535_adt_net_64588_\, 
        \I2.LEAD_FLAG6_637_adt_net_64628_\, 
        \I2.L2TYPE_4l15r_adt_net_66837_\, 
        \I2.N_4441_adt_net_67338_\, \I2.N_4445_adt_net_67839_\, 
        \I2.N_4449_adt_net_68340_\, 
        \I2.PIPE8_DT_558_adt_net_82590_\, 
        \I2.PIPE8_DT_21l29r_adt_net_82644_\, 
        \I2.PIPE8_DT_21_i_1l28r_adt_net_82784_\, 
        \I2.PIPE8_DT_21_i_1l28r_adt_net_82871_\, 
        \I2.N296_0_adt_net_86398_\, \I2.N296_0_adt_net_86403_\, 
        \I2.N312_0_adt_net_86445_\, \I2.N312_0_adt_net_86450_\, 
        \I2.N308_0_adt_net_86492_\, \I2.N308_0_adt_net_86497_\, 
        \I2.N316_i_i_adt_net_86577_\, 
        \I2.N316_i_i_adt_net_86582_\, \I2.N359_adt_net_86622_\, 
        \I2.N304_0_adt_net_86999_\, \I2.N304_0_adt_net_87004_\, 
        \I2.N300_0_adt_net_87046_\, \I2.N300_0_adt_net_87051_\, 
        \I2.N475_adt_net_87328__net_1\, \I2.N475_adt_net_87372_\, 
        \I2.N516_adt_net_87903__net_1\, 
        \I2.N498_1_adt_net_88035_\, \I2.N400_adt_net_88380_\, 
        \I2.N501_i_adt_net_88539_\, \I2.N504_adt_net_88887_\, 
        \I2.N481_adt_net_88982_\, \I2.N486_i_adt_net_89208_\, 
        \I2.N489_i_adt_net_89351_\, \I2.N492_i_adt_net_89450_\, 
        \I2.L_LUT_498_adt_net_90208_\, 
        \I2.INT_ERRBF1_495_adt_net_90378_\, 
        \I2.INT_ERRAF1_494_adt_net_90420_\, 
        \I2.N_3494_adt_net_90556_\, \I2.N_3494_adt_net_90563_\, 
        \I2.N_3823_adt_net_90689_\, \I2.N_2989_adt_net_92424_\, 
        \I2.N_2989_adt_net_92425_\, 
        \I2.CHAIN_ERR_DIS_448_adt_net_92599_\, 
        \I2.FID_7l9r_adt_net_92645_\, 
        \I2.FID_7l9r_adt_net_92653_\, 
        \I2.FID_7l8r_adt_net_92739_\, 
        \I2.FID_7l8r_adt_net_92747_\, 
        \I2.FID_7l7r_adt_net_92833_\, 
        \I2.FID_7l7r_adt_net_92841_\, 
        \I2.FID_7l6r_adt_net_92927_\, 
        \I2.FID_7l6r_adt_net_92935_\, 
        \I2.FID_7_0_iv_0l5r_adt_net_93017_\, 
        \I2.FID_7l4r_adt_net_93151_\, 
        \I2.FID_7l4r_adt_net_93158_\, 
        \I2.FID_7l4r_adt_net_93159_\, 
        \I2.FID_7l3r_adt_net_93251_\, 
        \I2.FID_7l3r_adt_net_93258_\, 
        \I2.FID_7l3r_adt_net_93259_\, 
        \I2.FID_7l2r_adt_net_93351_\, 
        \I2.FID_7l2r_adt_net_93358_\, 
        \I2.FID_7l2r_adt_net_93359_\, 
        \I2.FID_7_0_iv_0l1r_adt_net_93441_\, 
        \I2.FID_7l0r_adt_net_93569_\, 
        \I2.FID_7l0r_adt_net_93577_\, 
        \I2.NPRSFIF_328_adt_net_97261_\, 
        \I2.N_3828_adt_net_101749_\, \I2.N_3827_adt_net_101792_\, 
        \I1.N_370_adt_net_106310_\, \I1.N_370_adt_net_106316_\, 
        \I1.un1_sbyte13_1_i_1_adt_net_106369_\, 
        \I1.PAGECNTe_adt_net_106660_\, 
        \I1.sstate_ns_i_0_a4_0_1l0r_adt_net_107171_\, 
        \I1.sstate_ns_il5r_adt_net_107266_\, 
        \I1.sstate_nsl7r_adt_net_107573_\, 
        \I1.sstate_nsl7r_adt_net_107578_\, 
        \I1.sstate_nsl1r_adt_net_107663_\, 
        \I1.N_50_0_adt_net_109751__net_1\, 
        \I1.NCS0_56_adt_net_133847_\, 
        \I3.STATE1_nsl1r_adt_net_134330_\, 
        \I3.STATE1_nsl1r_adt_net_134332_\, 
        \I3.STATE1_nsl1r_adt_net_134337_\, 
        \I3.STATE1_nsl2r_adt_net_134784_\, 
        \I3.STATE1_nsl2r_adt_net_134789_\, 
        \I3.N_116_adt_net_134828_\, 
        \I3.PULSE_330_adt_net_134909_\, 
        \I3.N_2055_adt_net_134991_\, \I3.N_2055_adt_net_134992_\, 
        \I3.N_1510_adt_net_135035_\, \I3.N_1508_adt_net_135122_\, 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135386_\, 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135633_\, 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135637_\, 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135642_\, 
        \I3.STATE2_ns_i_i_a5_0_a3l1r_adt_net_135757_\, 
        \I3.un6_asb_NE_adt_net_135785_\, 
        \I3.un1_NOEDTKi_0_sqmuxa_adt_net_135826__net_1\, 
        \I3.STATE1_nsl0r_adt_net_135920_\, 
        \I3.STATE2_nsl0r_adt_net_136048_\, 
        \I3.STATE1_nsl8r_adt_net_136092_\, 
        \I3.STATE1_nsl7r_adt_net_136170_\, 
        \I3.STATE1_nsl7r_adt_net_136177_\, 
        \I3.STATE1_nsl5r_adt_net_136318_\, 
        \I3.STATE1_nsl5r_adt_net_136320_\, 
        \I3.STATE1_nsl3r_adt_net_136439_\, 
        \I3.STATE1_nsl3r_adt_net_136441_\, 
        \I3.N_1193_ip_adt_net_136530_\, 
        \I3.N_1193_ip_adt_net_136550_\, 
        \I3.N_1193_ip_adt_net_136551_\, 
        \I3.N_1193_ip_adt_net_136552_\, 
        \I3.N_1193_ip_adt_net_136553_\, 
        \I3.N_1193_ip_adt_net_136554_\, 
        \I3.N_1193_ip_adt_net_136555_\, 
        \I3.N_1193_ip_adt_net_136556_\, 
        \I3.N_1193_ip_adt_net_136557_\, 
        \I3.N_1193_ip_adt_net_136558_\, 
        \I3.VDBi_57l31r_adt_net_137838_\, 
        \I3.VDBi_57l31r_adt_net_137844_\, 
        \I3.un1_STATE1_13_1_adt_net_137890__net_1\, 
        \I3.un1_STATE1_13_1_adt_net_137902__net_1\, 
        \I3.VDBi_57l30r_adt_net_138033_\, 
        \I3.VDBi_57l30r_adt_net_138039_\, 
        \I3.VDBi_57l29r_adt_net_138169_\, 
        \I3.VDBi_57l29r_adt_net_138175_\, 
        \I3.VDBi_57l28r_adt_net_138305_\, 
        \I3.VDBi_57l28r_adt_net_138311_\, 
        \I3.VDBi_57l27r_adt_net_138431_\, 
        \I3.VDBi_57l27r_adt_net_138433_\, 
        \I3.VDBi_57l27r_adt_net_138440_\, 
        \I3.VDBi_57l27r_adt_net_138441_\, 
        \I3.VDBi_57l26r_adt_net_138571_\, 
        \I3.VDBi_57l26r_adt_net_138577_\, 
        \I3.VDBi_57l25r_adt_net_138707_\, 
        \I3.VDBi_57l25r_adt_net_138713_\, 
        \I3.VDBi_57l24r_adt_net_138805_\, 
        \I3.VDBi_57l24r_adt_net_138807_\, 
        \I3.VDBi_57l24r_adt_net_138814_\, 
        \I3.VDBi_57l24r_adt_net_138815_\, 
        \I3.VDBi_57l23r_adt_net_138945_\, 
        \I3.VDBi_57l23r_adt_net_138951_\, 
        \I3.VDBi_57l22r_adt_net_139083_\, 
        \I3.VDBi_57l22r_adt_net_139087_\, 
        \I3.VDBi_57l21r_adt_net_139179_\, 
        \I3.VDBi_57l21r_adt_net_139183_\, 
        \I3.VDBi_57l21r_adt_net_139188_\, 
        \I3.VDBi_57l21r_adt_net_139189_\, 
        \I3.VDBi_57l20r_adt_net_139281_\, 
        \I3.VDBi_57l20r_adt_net_139285_\, 
        \I3.VDBi_57l20r_adt_net_139290_\, 
        \I3.VDBi_57l20r_adt_net_139291_\, 
        \I3.VDBi_57l19r_adt_net_139383_\, 
        \I3.VDBi_57l19r_adt_net_139387_\, 
        \I3.VDBi_57l19r_adt_net_139392_\, 
        \I3.VDBi_57l19r_adt_net_139393_\, 
        \I3.VDBi_57l18r_adt_net_139485_\, 
        \I3.VDBi_57l18r_adt_net_139489_\, 
        \I3.VDBi_57l18r_adt_net_139494_\, 
        \I3.VDBi_57l18r_adt_net_139495_\, 
        \I3.VDBi_57l17r_adt_net_139627_\, 
        \I3.VDBi_57l17r_adt_net_139631_\, 
        \I3.VDBi_57l16r_adt_net_139761_\, 
        \I3.VDBi_57l16r_adt_net_139767_\, 
        \I3.VDBi_57l15r_adt_net_139959_\, 
        \I3.VDBi_57l15r_adt_net_139961_\, 
        \I3.VDBi_57l15r_adt_net_139969_\, 
        \I3.VDBi_57l15r_adt_net_139970_\, 
        \I3.VDBi_57l15r_adt_net_139971_\, 
        \I3.VDBi_57l15r_adt_net_139972_\, 
        \I3.VDBi_20l14r_adt_net_140054_\, 
        \I3.VDBi_57l14r_adt_net_140190_\, 
        \I3.VDBi_57l14r_adt_net_140192_\, 
        \I3.VDBi_57l14r_adt_net_140197_\, 
        \I3.VDBi_57l13r_adt_net_140454_\, 
        \I3.VDBi_57l13r_adt_net_140499_\, 
        \I3.VDBi_57l13r_adt_net_140578_\, 
        \I3.VDBi_57l13r_adt_net_140582_\, 
        \I3.VDBi_57l13r_adt_net_140592_\, 
        \I3.VDBi_57l13r_adt_net_140593_\, 
        \I3.VDBi_57l13r_adt_net_140594_\, 
        \I3.VDBi_57l13r_adt_net_140595_\, 
        \I3.VDBi_57l13r_adt_net_140596_\, 
        \I3.VDBi_57l13r_adt_net_140597_\, 
        \I3.VDBi_20l12r_adt_net_140765_\, 
        \I3.VDBi_57l12r_adt_net_140988_\, 
        \I3.VDBi_57l12r_adt_net_140997_\, 
        \I3.VDBi_57l12r_adt_net_140998_\, 
        \I3.VDBi_20l11r_adt_net_141166_\, 
        \I3.VDBi_57l11r_adt_net_141431_\, 
        \I3.VDBi_57l11r_adt_net_141440_\, 
        \I3.VDBi_57l11r_adt_net_141441_\, 
        \I3.VDBi_20l10r_adt_net_141609_\, 
        \I3.VDBi_57l10r_adt_net_141874_\, 
        \I3.VDBi_57l10r_adt_net_141883_\, 
        \I3.VDBi_57l10r_adt_net_141884_\, 
        \I3.VDBi_29l9r_adt_net_142014__net_1\, 
        \I3.VDBi_29l9r_adt_net_142020__net_1\, 
        \I3.VDBi_57l9r_adt_net_142322_\, 
        \I3.VDBi_57l9r_adt_net_142331_\, 
        \I3.VDBi_57l9r_adt_net_142332_\, 
        \I3.VDBi_20l8r_adt_net_142456_\, 
        \I3.VDBi_57l8r_adt_net_142588__net_1\, 
        \I3.VDBi_57l8r_adt_net_142596__net_1\, 
        \I3.VDBi_57l8r_adt_net_142678_\, 
        \I3.VDBi_57l8r_adt_net_142723_\, 
        \I3.VDBi_57l8r_adt_net_142780_\, 
        \I3.VDBi_57l8r_adt_net_142784_\, 
        \I3.VDBi_57l8r_adt_net_142786_\, 
        \I3.VDBi_57l8r_adt_net_142792_\, 
        \I3.VDBi_57l8r_adt_net_142793_\, 
        \I3.VDBi_57l7r_adt_net_142952__net_1\, 
        \I3.VDBi_57l7r_adt_net_142961__net_1\, 
        \I3.VDBi_57l7r_adt_net_143017__net_1\, 
        \I3.VDBi_57l7r_adt_net_143023__net_1\, 
        \I3.VDBi_57l7r_adt_net_143034__net_1\, 
        \I3.VDBi_57l7r_adt_net_143035__net_1\, 
        \I3.VDBi_57l7r_adt_net_143036__net_1\, 
        \I3.VDBi_57l7r_adt_net_143037__net_1\, 
        \I3.VDBi_57l7r_adt_net_143093_\, 
        \I3.VDBi_57l7r_adt_net_143099_\, 
        \I3.VDBi_57l7r_adt_net_143103_\, 
        \I3.VDBi_57l7r_adt_net_143110_\, 
        \I3.VDBi_57l7r_adt_net_143111_\, 
        \I3.VDBi_57l7r_adt_net_143112_\, 
        \I3.VDBi_57l6r_adt_net_143243__net_1\, 
        \I3.VDBi_57l6r_adt_net_143252__net_1\, 
        \I3.VDBi_57l6r_adt_net_143308__net_1\, 
        \I3.VDBi_57l6r_adt_net_143314__net_1\, 
        \I3.VDBi_57l6r_adt_net_143325__net_1\, 
        \I3.VDBi_57l6r_adt_net_143326__net_1\, 
        \I3.VDBi_57l6r_adt_net_143327__net_1\, 
        \I3.VDBi_57l6r_adt_net_143328__net_1\, 
        \I3.VDBi_57l6r_adt_net_143384_\, 
        \I3.VDBi_57l6r_adt_net_143390_\, 
        \I3.VDBi_57l6r_adt_net_143394_\, 
        \I3.VDBi_57l6r_adt_net_143401_\, 
        \I3.VDBi_57l6r_adt_net_143402_\, 
        \I3.VDBi_57l6r_adt_net_143403_\, 
        \I3.N_283_adt_net_143528_\, 
        \I3.VDBi_31_i_a3_0_1l5r_adt_net_143649_\, 
        \I3.VDBi_31_i_a3_0_1l5r_adt_net_143654_\, 
        \I3.N_1772_adt_net_143698_\, \I3.N_1772_adt_net_143704_\, 
        \I3.VDBi_40l5r_adt_net_143744_\, 
        \I3.VDBi_57l5r_adt_net_143846_\, 
        \I3.VDBi_57l5r_adt_net_143850_\, 
        \I3.VDBi_57l5r_adt_net_143854_\, 
        \I3.VDBi_57l5r_adt_net_143861_\, 
        \I3.VDBi_57l5r_adt_net_143862_\, 
        \I3.VDBi_57l5r_adt_net_143863_\, 
        \I3.VDBi_29l4r_adt_net_144161_\, 
        \I3.VDBi_57l4r_adt_net_144429_\, 
        \I3.VDBi_57l4r_adt_net_144439_\, 
        \I3.VDBi_57l4r_adt_net_144440_\, 
        \I3.VDBi_57l4r_adt_net_144441_\, 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144601_\, 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144610_\, 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144611_\, 
        \I3.VDBi_20l3r_adt_net_144750_\, 
        \I3.VDBi_57l3r_adt_net_145062_\, 
        \I3.VDBi_57l3r_adt_net_145072_\, 
        \I3.VDBi_57l3r_adt_net_145073_\, 
        \I3.VDBi_57l3r_adt_net_145074_\, 
        \I3.VDBi_57l2r_adt_net_145218__net_1\, 
        \I3.VDBi_57l2r_adt_net_145225__net_1\, 
        \I3.VDBi_57l2r_adt_net_145226__net_1\, 
        \I3.VDBi_57l2r_adt_net_145227__net_1\, 
        \I3.VDBi_57l2r_adt_net_145285__net_1\, 
        \I3.VDBi_57l2r_adt_net_145295__net_1\, 
        \I3.VDBi_57l2r_adt_net_145303__net_1\, 
        \I3.VDBi_57l2r_adt_net_145304__net_1\, 
        \I3.VDBi_57l2r_adt_net_145305__net_1\, 
        \I3.VDBi_57l2r_adt_net_145306__net_1\, 
        \I3.VDBi_57l2r_adt_net_145362_\, 
        \I3.VDBi_57l2r_adt_net_145368_\, 
        \I3.VDBi_57l2r_adt_net_145372_\, 
        \I3.VDBi_57l2r_adt_net_145379_\, 
        \I3.VDBi_57l2r_adt_net_145380_\, 
        \I3.VDBi_57l2r_adt_net_145381_\, 
        \I3.VDBi_23l1r_adt_net_145526__net_1\, 
        \I3.VDBi_23l1r_adt_net_145528__net_1\, 
        \I3.VDBi_23l1r_adt_net_145530__net_1\, 
        \I3.VDBi_23l1r_adt_net_145532__net_1\, 
        \I3.VDBi_23l1r_adt_net_145541__net_1\, 
        \I3.VDBi_23l1r_adt_net_145542__net_1\, 
        \I3.VDBi_23l1r_adt_net_145581_\, 
        \I3.VDBi_57l1r_adt_net_145935_\, 
        \I3.VDBi_57l1r_adt_net_145945_\, 
        \I3.VDBi_57l1r_adt_net_145946_\, 
        \I3.VDBi_57l1r_adt_net_145947_\, 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_adt_net_146105_\, 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_adt_net_146111_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146197__net_1\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146205__net_1\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146304_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146347_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146420_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146422_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146424_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146426_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146432_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146446_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146447_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146448_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146450_\, 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146451_\, 
        \I3.VDBi_57l0r_adt_net_146601_\, 
        \I3.VDBi_57l0r_adt_net_146651_\, 
        \I3.VDBi_57l0r_adt_net_146655_\, 
        \I3.VDBi_57l0r_adt_net_146660_\, 
        \I3.PULSE_46l9r_adt_net_146747_\, 
        \I3.PULSE_46l8r_adt_net_146836_\, 
        \I3.PULSE_46l6r_adt_net_147009_\, 
        \I3.PULSE_46l6r_adt_net_147015_\, 
        \I3.PULSE_46l5r_adt_net_147097_\, 
        \I3.N_55_adt_net_147183_\, \I3.N_122_adt_net_147352_\, 
        \I3.PULSE_332_adt_net_147433_\, 
        \I3.N_118_adt_net_147476_\, 
        \I3.PULSE_331_adt_net_147557_\, 
        \I3.un15_anycyc_adt_net_147611_\, 
        \I3.un15_anycyc_adt_net_147613_\, 
        \I3.un15_anycyc_adt_net_147616_\, 
        \I3.un15_anycyc_adt_net_147620_\, 
        \I3.N_297_adt_net_147649_\, 
        \I3.un1_STATE2_15_1_adt_net_147708__net_1\, 
        \I3.N_1636_adt_net_150083_\, \I3.N_1635_adt_net_150153_\, 
        \I3.N_1634_adt_net_150223_\, \I3.N_1633_adt_net_150293_\, 
        \I3.N_1632_adt_net_150363_\, \I3.N_1631_adt_net_150433_\, 
        \I3.N_1630_adt_net_150503_\, 
        \I3.un1_STATE2_13_adt_net_150833__net_1\, 
        \I3.un1_STATE2_13_adt_net_150841__net_1\, 
        \I3.un1_NRDMEBi_2_sqmuxa_3_0_adt_net_153527_\, 
        \I3.un1_NRDMEBi_2_sqmuxa_3_adt_net_153598_\, 
        \I3.un1_STATE2_11_adt_net_153679__net_1\, 
        \I3.un1_STATE2_11_adt_net_153728_\, 
        \I3.un1_EVREAD_DS_1_sqmuxa_1_adt_net_158292_\, 
        \I3.N_80_adt_net_159051_\, 
        \I3.un1_NOEDTKi_0_sqmuxa_adt_net_159270_\, 
        \I3.un1_NOEDTKi_0_sqmuxa_1_adt_net_159322_\, 
        \I3.un1_NOEDTKi_0_sqmuxa_1_adt_net_159328_\, 
        \I3.PIPEB_110_adt_net_159411_\, 
        \I3.PIPEB_106_adt_net_159579_\, 
        \I3.PIPEB_105_adt_net_159621_\, 
        \I3.PIPEB_104_adt_net_159663_\, 
        \I3.PIPEB_103_adt_net_159705_\, 
        \I3.PIPEB_102_adt_net_159747_\, 
        \I3.PIPEB_101_adt_net_159789_\, 
        \I3.PIPEB_100_adt_net_159831_\, 
        \I3.PIPEB_99_adt_net_159873_\, 
        \I3.PIPEB_98_adt_net_159915_\, 
        \I3.PIPEB_97_adt_net_159957_\, 
        \I3.PIPEB_96_adt_net_159999_\, 
        \I3.PIPEB_95_adt_net_160041_\, 
        \I3.PIPEB_94_adt_net_160083_\, 
        \I3.PIPEB_93_adt_net_160125_\, 
        \I3.PIPEB_92_adt_net_160167_\, 
        \I3.PIPEB_91_adt_net_160209_\, 
        \I3.PIPEB_90_adt_net_160251_\, 
        \I3.PIPEB_89_adt_net_160293_\, 
        \I3.PIPEB_88_adt_net_160335_\, 
        \I3.PIPEB_87_adt_net_160377_\, 
        \I3.PIPEB_86_adt_net_160419_\, 
        \I3.PIPEB_85_adt_net_160461_\, 
        \I3.PIPEB_84_adt_net_160503_\, 
        \I3.PIPEB_83_adt_net_160545_\, 
        \I3.PIPEB_82_adt_net_160587_\, 
        \I3.PIPEB_81_adt_net_160629_\, 
        \I3.PIPEB_80_adt_net_160671_\, 
        \I3.PIPEB_79_adt_net_160713_\, 
        \I3.N_1902_adt_net_160759_\, 
        \I3.un1_MYBERRi_1_sqmuxa_adt_net_161480_\, 
        \I3.un1_MYBERRi_1_sqmuxa_adt_net_161483_\, 
        \I3.N_306_adt_net_161608_\, 
        \I3.VDBoffb_30l7r_adt_net_161744_\, 
        \I3.VDBoffb_30l7r_adt_net_161748_\, 
        \I3.VDBoffb_30l7r_adt_net_161752_\, 
        \I3.VDBoffb_30l7r_adt_net_161756_\, 
        \I3.VDBoffb_30l7r_adt_net_161760_\, 
        \I3.VDBoffb_30l7r_adt_net_161764_\, 
        \I3.VDBoffb_30l7r_adt_net_161768_\, 
        \I3.VDBoffb_30l7r_adt_net_161788_\, 
        \I3.VDBoffb_30l7r_adt_net_161789_\, 
        \I3.VDBoffb_30l7r_adt_net_161790_\, 
        \I3.VDBoffb_30l7r_adt_net_161791_\, 
        \I3.VDBoffb_30l7r_adt_net_161792_\, 
        \I3.VDBoffb_30l7r_adt_net_161793_\, 
        \I3.VDBoffb_30l7r_adt_net_161794_\, 
        \I3.VDBoffb_30l7r_adt_net_161795_\, 
        \I3.VDBoffb_30l7r_adt_net_161797_\, 
        \I3.VDBoffb_30l7r_adt_net_161799_\, 
        \I3.VDBoffb_30l7r_adt_net_161800_\, 
        \I3.VDBoffb_59_adt_net_161840_\, 
        \I3.VDBoffb_30l6r_adt_net_161934_\, 
        \I3.VDBoffb_30l6r_adt_net_161938_\, 
        \I3.VDBoffb_30l6r_adt_net_161942_\, 
        \I3.VDBoffb_30l6r_adt_net_161946_\, 
        \I3.VDBoffb_30l6r_adt_net_161950_\, 
        \I3.VDBoffb_30l6r_adt_net_161954_\, 
        \I3.VDBoffb_30l6r_adt_net_161958_\, 
        \I3.VDBoffb_30l6r_adt_net_161978_\, 
        \I3.VDBoffb_30l6r_adt_net_161979_\, 
        \I3.VDBoffb_30l6r_adt_net_161980_\, 
        \I3.VDBoffb_30l6r_adt_net_161981_\, 
        \I3.VDBoffb_30l6r_adt_net_161982_\, 
        \I3.VDBoffb_30l6r_adt_net_161983_\, 
        \I3.VDBoffb_30l6r_adt_net_161984_\, 
        \I3.VDBoffb_30l6r_adt_net_161985_\, 
        \I3.VDBoffb_30l6r_adt_net_161987_\, 
        \I3.VDBoffb_30l6r_adt_net_161989_\, 
        \I3.VDBoffb_30l6r_adt_net_161990_\, 
        \I3.VDBoffb_58_adt_net_162030_\, 
        \I3.VDBoffb_30l5r_adt_net_162124_\, 
        \I3.VDBoffb_30l5r_adt_net_162128_\, 
        \I3.VDBoffb_30l5r_adt_net_162132_\, 
        \I3.VDBoffb_30l5r_adt_net_162136_\, 
        \I3.VDBoffb_30l5r_adt_net_162140_\, 
        \I3.VDBoffb_30l5r_adt_net_162144_\, 
        \I3.VDBoffb_30l5r_adt_net_162148_\, 
        \I3.VDBoffb_30l5r_adt_net_162168_\, 
        \I3.VDBoffb_30l5r_adt_net_162169_\, 
        \I3.VDBoffb_30l5r_adt_net_162170_\, 
        \I3.VDBoffb_30l5r_adt_net_162171_\, 
        \I3.VDBoffb_30l5r_adt_net_162172_\, 
        \I3.VDBoffb_30l5r_adt_net_162173_\, 
        \I3.VDBoffb_30l5r_adt_net_162174_\, 
        \I3.VDBoffb_30l5r_adt_net_162175_\, 
        \I3.VDBoffb_30l5r_adt_net_162177_\, 
        \I3.VDBoffb_30l5r_adt_net_162179_\, 
        \I3.VDBoffb_30l5r_adt_net_162180_\, 
        \I3.VDBoffb_57_adt_net_162220_\, 
        \I3.VDBoffb_30l4r_adt_net_162314_\, 
        \I3.VDBoffb_30l4r_adt_net_162318_\, 
        \I3.VDBoffb_30l4r_adt_net_162322_\, 
        \I3.VDBoffb_30l4r_adt_net_162326_\, 
        \I3.VDBoffb_30l4r_adt_net_162330_\, 
        \I3.VDBoffb_30l4r_adt_net_162334_\, 
        \I3.VDBoffb_30l4r_adt_net_162338_\, 
        \I3.VDBoffb_30l4r_adt_net_162358_\, 
        \I3.VDBoffb_30l4r_adt_net_162359_\, 
        \I3.VDBoffb_30l4r_adt_net_162360_\, 
        \I3.VDBoffb_30l4r_adt_net_162361_\, 
        \I3.VDBoffb_30l4r_adt_net_162362_\, 
        \I3.VDBoffb_30l4r_adt_net_162363_\, 
        \I3.VDBoffb_30l4r_adt_net_162364_\, 
        \I3.VDBoffb_30l4r_adt_net_162365_\, 
        \I3.VDBoffb_30l4r_adt_net_162367_\, 
        \I3.VDBoffb_30l4r_adt_net_162369_\, 
        \I3.VDBoffb_30l4r_adt_net_162370_\, 
        \I3.VDBoffb_56_adt_net_162410_\, 
        \I3.VDBoffb_30l3r_adt_net_162504_\, 
        \I3.VDBoffb_30l3r_adt_net_162508_\, 
        \I3.VDBoffb_30l3r_adt_net_162512_\, 
        \I3.VDBoffb_30l3r_adt_net_162516_\, 
        \I3.VDBoffb_30l3r_adt_net_162520_\, 
        \I3.VDBoffb_30l3r_adt_net_162524_\, 
        \I3.VDBoffb_30l3r_adt_net_162528_\, 
        \I3.VDBoffb_30l3r_adt_net_162548_\, 
        \I3.VDBoffb_30l3r_adt_net_162549_\, 
        \I3.VDBoffb_30l3r_adt_net_162550_\, 
        \I3.VDBoffb_30l3r_adt_net_162551_\, 
        \I3.VDBoffb_30l3r_adt_net_162552_\, 
        \I3.VDBoffb_30l3r_adt_net_162553_\, 
        \I3.VDBoffb_30l3r_adt_net_162554_\, 
        \I3.VDBoffb_30l3r_adt_net_162555_\, 
        \I3.VDBoffb_30l3r_adt_net_162557_\, 
        \I3.VDBoffb_30l3r_adt_net_162559_\, 
        \I3.VDBoffb_30l3r_adt_net_162560_\, 
        \I3.VDBoffb_55_adt_net_162600_\, 
        \I3.VDBoffb_30l2r_adt_net_162694_\, 
        \I3.VDBoffb_30l2r_adt_net_162698_\, 
        \I3.VDBoffb_30l2r_adt_net_162702_\, 
        \I3.VDBoffb_30l2r_adt_net_162706_\, 
        \I3.VDBoffb_30l2r_adt_net_162710_\, 
        \I3.VDBoffb_30l2r_adt_net_162714_\, 
        \I3.VDBoffb_30l2r_adt_net_162718_\, 
        \I3.VDBoffb_30l2r_adt_net_162738_\, 
        \I3.VDBoffb_30l2r_adt_net_162739_\, 
        \I3.VDBoffb_30l2r_adt_net_162740_\, 
        \I3.VDBoffb_30l2r_adt_net_162741_\, 
        \I3.VDBoffb_30l2r_adt_net_162742_\, 
        \I3.VDBoffb_30l2r_adt_net_162743_\, 
        \I3.VDBoffb_30l2r_adt_net_162744_\, 
        \I3.VDBoffb_30l2r_adt_net_162745_\, 
        \I3.VDBoffb_30l2r_adt_net_162747_\, 
        \I3.VDBoffb_30l2r_adt_net_162749_\, 
        \I3.VDBoffb_30l2r_adt_net_162750_\, 
        \I3.VDBoffb_54_adt_net_162790_\, 
        \I3.VDBoffb_30l1r_adt_net_162884_\, 
        \I3.VDBoffb_30l1r_adt_net_162888_\, 
        \I3.VDBoffb_30l1r_adt_net_162892_\, 
        \I3.VDBoffb_30l1r_adt_net_162896_\, 
        \I3.VDBoffb_30l1r_adt_net_162900_\, 
        \I3.VDBoffb_30l1r_adt_net_162904_\, 
        \I3.VDBoffb_30l1r_adt_net_162908_\, 
        \I3.VDBoffb_30l1r_adt_net_162928_\, 
        \I3.VDBoffb_30l1r_adt_net_162929_\, 
        \I3.VDBoffb_30l1r_adt_net_162930_\, 
        \I3.VDBoffb_30l1r_adt_net_162931_\, 
        \I3.VDBoffb_30l1r_adt_net_162932_\, 
        \I3.VDBoffb_30l1r_adt_net_162933_\, 
        \I3.VDBoffb_30l1r_adt_net_162934_\, 
        \I3.VDBoffb_30l1r_adt_net_162935_\, 
        \I3.VDBoffb_30l1r_adt_net_162937_\, 
        \I3.VDBoffb_30l1r_adt_net_162939_\, 
        \I3.VDBoffb_30l1r_adt_net_162940_\, 
        \I3.VDBoffb_53_adt_net_162980_\, 
        \I3.VDBoffb_30l0r_adt_net_163074_\, 
        \I3.VDBoffb_30l0r_adt_net_163078_\, 
        \I3.VDBoffb_30l0r_adt_net_163082_\, 
        \I3.VDBoffb_30l0r_adt_net_163086_\, 
        \I3.VDBoffb_30l0r_adt_net_163090_\, 
        \I3.VDBoffb_30l0r_adt_net_163094_\, 
        \I3.VDBoffb_30l0r_adt_net_163098_\, 
        \I3.VDBoffb_30l0r_adt_net_163118_\, 
        \I3.VDBoffb_30l0r_adt_net_163119_\, 
        \I3.VDBoffb_30l0r_adt_net_163120_\, 
        \I3.VDBoffb_30l0r_adt_net_163121_\, 
        \I3.VDBoffb_30l0r_adt_net_163122_\, 
        \I3.VDBoffb_30l0r_adt_net_163123_\, 
        \I3.VDBoffb_30l0r_adt_net_163124_\, 
        \I3.VDBoffb_30l0r_adt_net_163125_\, 
        \I3.VDBoffb_30l0r_adt_net_163127_\, 
        \I3.VDBoffb_30l0r_adt_net_163129_\, 
        \I3.VDBoffb_30l0r_adt_net_163130_\, 
        \I3.VDBoffb_52_adt_net_163170_\, 
        \I3.VDBoffa_31l7r_adt_net_163264_\, 
        \I3.VDBoffa_31l7r_adt_net_163268_\, 
        \I3.VDBoffa_31l7r_adt_net_163272_\, 
        \I3.VDBoffa_31l7r_adt_net_163276_\, 
        \I3.VDBoffa_31l7r_adt_net_163280_\, 
        \I3.VDBoffa_31l7r_adt_net_163284_\, 
        \I3.VDBoffa_31l7r_adt_net_163288_\, 
        \I3.VDBoffa_31l7r_adt_net_163308_\, 
        \I3.VDBoffa_31l7r_adt_net_163309_\, 
        \I3.VDBoffa_31l7r_adt_net_163310_\, 
        \I3.VDBoffa_31l7r_adt_net_163311_\, 
        \I3.VDBoffa_31l7r_adt_net_163312_\, 
        \I3.VDBoffa_31l7r_adt_net_163313_\, 
        \I3.VDBoffa_31l7r_adt_net_163314_\, 
        \I3.VDBoffa_31l7r_adt_net_163315_\, 
        \I3.VDBoffa_31l7r_adt_net_163317_\, 
        \I3.VDBoffa_31l7r_adt_net_163319_\, 
        \I3.VDBoffa_31l7r_adt_net_163320_\, 
        \I3.VDBoffa_51_adt_net_163358_\, 
        \I3.N_2070_adt_net_163454_\, \I3.N_2070_adt_net_163458_\, 
        \I3.N_2070_adt_net_163462_\, \I3.N_2070_adt_net_163466_\, 
        \I3.N_2070_adt_net_163470_\, \I3.N_2070_adt_net_163474_\, 
        \I3.N_2070_adt_net_163478_\, \I3.N_2070_adt_net_163498_\, 
        \I3.N_2070_adt_net_163499_\, \I3.N_2070_adt_net_163500_\, 
        \I3.N_2070_adt_net_163501_\, \I3.N_2070_adt_net_163502_\, 
        \I3.N_2070_adt_net_163503_\, \I3.N_2070_adt_net_163504_\, 
        \I3.N_2070_adt_net_163505_\, \I3.N_2070_adt_net_163507_\, 
        \I3.N_2070_adt_net_163509_\, \I3.N_2070_adt_net_163510_\, 
        \I3.VDBoffa_50_adt_net_163548_\, 
        \I3.VDBoffa_31l5r_adt_net_163644_\, 
        \I3.VDBoffa_31l5r_adt_net_163648_\, 
        \I3.VDBoffa_31l5r_adt_net_163652_\, 
        \I3.VDBoffa_31l5r_adt_net_163656_\, 
        \I3.VDBoffa_31l5r_adt_net_163660_\, 
        \I3.VDBoffa_31l5r_adt_net_163664_\, 
        \I3.VDBoffa_31l5r_adt_net_163668_\, 
        \I3.VDBoffa_31l5r_adt_net_163688_\, 
        \I3.VDBoffa_31l5r_adt_net_163689_\, 
        \I3.VDBoffa_31l5r_adt_net_163690_\, 
        \I3.VDBoffa_31l5r_adt_net_163691_\, 
        \I3.VDBoffa_31l5r_adt_net_163692_\, 
        \I3.VDBoffa_31l5r_adt_net_163693_\, 
        \I3.VDBoffa_31l5r_adt_net_163694_\, 
        \I3.VDBoffa_31l5r_adt_net_163695_\, 
        \I3.VDBoffa_31l5r_adt_net_163697_\, 
        \I3.VDBoffa_31l5r_adt_net_163699_\, 
        \I3.VDBoffa_31l5r_adt_net_163700_\, 
        \I3.VDBoffa_49_adt_net_163738_\, 
        \I3.VDBoffa_31l4r_adt_net_163834_\, 
        \I3.VDBoffa_31l4r_adt_net_163838_\, 
        \I3.VDBoffa_31l4r_adt_net_163842_\, 
        \I3.VDBoffa_31l4r_adt_net_163846_\, 
        \I3.VDBoffa_31l4r_adt_net_163850_\, 
        \I3.VDBoffa_31l4r_adt_net_163854_\, 
        \I3.VDBoffa_31l4r_adt_net_163858_\, 
        \I3.VDBoffa_31l4r_adt_net_163878_\, 
        \I3.VDBoffa_31l4r_adt_net_163879_\, 
        \I3.VDBoffa_31l4r_adt_net_163880_\, 
        \I3.VDBoffa_31l4r_adt_net_163881_\, 
        \I3.VDBoffa_31l4r_adt_net_163882_\, 
        \I3.VDBoffa_31l4r_adt_net_163883_\, 
        \I3.VDBoffa_31l4r_adt_net_163884_\, 
        \I3.VDBoffa_31l4r_adt_net_163885_\, 
        \I3.VDBoffa_31l4r_adt_net_163887_\, 
        \I3.VDBoffa_31l4r_adt_net_163889_\, 
        \I3.VDBoffa_31l4r_adt_net_163890_\, 
        \I3.VDBoffa_48_adt_net_163928_\, 
        \I3.VDBoffa_31l3r_adt_net_164024_\, 
        \I3.VDBoffa_31l3r_adt_net_164028_\, 
        \I3.VDBoffa_31l3r_adt_net_164032_\, 
        \I3.VDBoffa_31l3r_adt_net_164036_\, 
        \I3.VDBoffa_31l3r_adt_net_164040_\, 
        \I3.VDBoffa_31l3r_adt_net_164044_\, 
        \I3.VDBoffa_31l3r_adt_net_164048_\, 
        \I3.VDBoffa_31l3r_adt_net_164068_\, 
        \I3.VDBoffa_31l3r_adt_net_164069_\, 
        \I3.VDBoffa_31l3r_adt_net_164070_\, 
        \I3.VDBoffa_31l3r_adt_net_164071_\, 
        \I3.VDBoffa_31l3r_adt_net_164072_\, 
        \I3.VDBoffa_31l3r_adt_net_164073_\, 
        \I3.VDBoffa_31l3r_adt_net_164074_\, 
        \I3.VDBoffa_31l3r_adt_net_164075_\, 
        \I3.VDBoffa_31l3r_adt_net_164077_\, 
        \I3.VDBoffa_31l3r_adt_net_164079_\, 
        \I3.VDBoffa_31l3r_adt_net_164080_\, 
        \I3.VDBoffa_47_adt_net_164118_\, 
        \I3.VDBoffa_31l2r_adt_net_164214_\, 
        \I3.VDBoffa_31l2r_adt_net_164218_\, 
        \I3.VDBoffa_31l2r_adt_net_164222_\, 
        \I3.VDBoffa_31l2r_adt_net_164226_\, 
        \I3.VDBoffa_31l2r_adt_net_164230_\, 
        \I3.VDBoffa_31l2r_adt_net_164234_\, 
        \I3.VDBoffa_31l2r_adt_net_164238_\, 
        \I3.VDBoffa_31l2r_adt_net_164258_\, 
        \I3.VDBoffa_31l2r_adt_net_164259_\, 
        \I3.VDBoffa_31l2r_adt_net_164260_\, 
        \I3.VDBoffa_31l2r_adt_net_164261_\, 
        \I3.VDBoffa_31l2r_adt_net_164262_\, 
        \I3.VDBoffa_31l2r_adt_net_164263_\, 
        \I3.VDBoffa_31l2r_adt_net_164264_\, 
        \I3.VDBoffa_31l2r_adt_net_164265_\, 
        \I3.VDBoffa_31l2r_adt_net_164267_\, 
        \I3.VDBoffa_31l2r_adt_net_164269_\, 
        \I3.VDBoffa_31l2r_adt_net_164270_\, 
        \I3.VDBoffa_46_adt_net_164308_\, 
        \I3.VDBoffa_31l1r_adt_net_164404_\, 
        \I3.VDBoffa_31l1r_adt_net_164408_\, 
        \I3.VDBoffa_31l1r_adt_net_164412_\, 
        \I3.VDBoffa_31l1r_adt_net_164416_\, 
        \I3.VDBoffa_31l1r_adt_net_164420_\, 
        \I3.VDBoffa_31l1r_adt_net_164424_\, 
        \I3.VDBoffa_31l1r_adt_net_164428_\, 
        \I3.VDBoffa_31l1r_adt_net_164448_\, 
        \I3.VDBoffa_31l1r_adt_net_164449_\, 
        \I3.VDBoffa_31l1r_adt_net_164450_\, 
        \I3.VDBoffa_31l1r_adt_net_164451_\, 
        \I3.VDBoffa_31l1r_adt_net_164452_\, 
        \I3.VDBoffa_31l1r_adt_net_164453_\, 
        \I3.VDBoffa_31l1r_adt_net_164454_\, 
        \I3.VDBoffa_31l1r_adt_net_164455_\, 
        \I3.VDBoffa_31l1r_adt_net_164457_\, 
        \I3.VDBoffa_31l1r_adt_net_164459_\, 
        \I3.VDBoffa_31l1r_adt_net_164460_\, 
        \I3.VDBoffa_45_adt_net_164498_\, 
        \I3.VDBoffa_31l0r_adt_net_164594_\, 
        \I3.VDBoffa_31l0r_adt_net_164598_\, 
        \I3.VDBoffa_31l0r_adt_net_164602_\, 
        \I3.VDBoffa_31l0r_adt_net_164606_\, 
        \I3.VDBoffa_31l0r_adt_net_164610_\, 
        \I3.VDBoffa_31l0r_adt_net_164614_\, 
        \I3.VDBoffa_31l0r_adt_net_164618_\, 
        \I3.VDBoffa_31l0r_adt_net_164638_\, 
        \I3.VDBoffa_31l0r_adt_net_164639_\, 
        \I3.VDBoffa_31l0r_adt_net_164640_\, 
        \I3.VDBoffa_31l0r_adt_net_164641_\, 
        \I3.VDBoffa_31l0r_adt_net_164642_\, 
        \I3.VDBoffa_31l0r_adt_net_164643_\, 
        \I3.VDBoffa_31l0r_adt_net_164644_\, 
        \I3.VDBoffa_31l0r_adt_net_164645_\, 
        \I3.VDBoffa_31l0r_adt_net_164647_\, 
        \I3.VDBoffa_31l0r_adt_net_164649_\, 
        \I3.VDBoffa_31l0r_adt_net_164650_\, 
        \I3.VDBoffa_44_adt_net_164688_\, 
        \I2.N411_adt_net_194931__net_1\, 
        \I2.N411_adt_net_194981__net_1\, 
        \I2.N495_i_adt_net_202032_\, \I2.N495_i_adt_net_202093_\, 
        \I2.N495_i_adt_net_202144_\, \I2.N495_i_adt_net_207682_\, 
        \I2.I180_un1_Y_adt_net_215260_\, 
        \I2.N510_adt_net_220872_\, \I2.N510_adt_net_220925_\, 
        \I2.N510_adt_net_232425_\, 
        \I2.I180_un1_Y_adt_net_240062_\, 
        \I2.I180_un1_Y_adt_net_240115_\, 
        \I2.I180_un1_Y_adt_net_252355_\, 
        \I3.VDBi_13l4r_adt_net_284333_\, 
        \I3.VDBi_13l4r_adt_net_284335_\, 
        \I2.N479_adt_net_296182__net_1\, 
        \I2.N477_adt_net_301898__net_1\, 
        \I2.N477_adt_net_302171__net_1\, 
        \I2.N477_adt_net_302175__net_1\, 
        \I2.N477_adt_net_302179__net_1\, 
        \I2.I180_un1_Y_adt_net_309337_\, 
        \I2.N477_adt_net_371248_\, \I2.N477_adt_net_371301_\, 
        \I2.N475_adt_net_378647__net_1\, 
        \I3.VDBi_29l1r_adt_net_411517_\, 
        \I3.VDBi_20l4r_adt_net_414879_\, 
        \I2.N481_adt_net_423940_\, \I2.N481_adt_net_424213_\, 
        \I2.N481_adt_net_424217_\, \I2.N481_adt_net_424221_\, 
        \I2.N477_adt_net_438351_\, 
        \I2.N475_adt_net_442369__net_1\, 
        \I2.N475_adt_net_442371__net_1\, 
        \I2.N475_adt_net_460353__net_1\, 
        \I3.VDBi_31l1r_adt_net_506164_\, 
        \I3.VDBi_29l3r_adt_net_510711_\, 
        \I3.VDBi_29l3r_adt_net_510792_\, 
        \I3.VDBi_20l4r_adt_net_514155_\, 
        \I2.SUB8_520_adt_net_531295_\, 
        \I2.SUB8_520_adt_net_531407_\, \I2.N479_adt_net_538167_\, 
        \I2.N479_adt_net_538220_\, \I2.N479_adt_net_538261_\, 
        \I2.SUB8_522_adt_net_551987_\, 
        \I2.SUB8_522_adt_net_552099_\, 
        \I2.SUB8_523_adt_net_566364_\, 
        \I2.SUB8_523_adt_net_566476_\, 
        \I3.VDBi_31l1r_adt_net_614331_\, 
        \I3.VDBi_29l3r_adt_net_618363_\, 
        \I3.VDBi_29l4r_adt_net_621921_\, 
        \I2.SUB8_520_adt_net_635603_\, 
        \I2.SUB8_520_adt_net_635605_\, 
        \I2.SUB8_520_adt_net_635607_\, 
        \I2.SUB8_520_adt_net_635612_\, \I2.N479_adt_net_642172_\, 
        \I2.N479_adt_net_642225_\, \I2.N479_adt_net_642266_\, 
        \I2.N479_adt_net_649015_\, \I2.SUB8_522_adt_net_659160_\, 
        \I2.SUB8_522_adt_net_659162_\, 
        \I2.SUB8_522_adt_net_659164_\, 
        \I2.SUB8_522_adt_net_659169_\, 
        \I2.SUB8_523_adt_net_670055_\, 
        \I2.SUB8_523_adt_net_670057_\, 
        \I2.SUB8_523_adt_net_670059_\, 
        \I2.SUB8_523_adt_net_670064_\, \I3.TCNT3_c1\, \I5.N_74\, 
        \I5.N_81_i_0_i\, \I5.AIR_WDATA_9l11r_net_1\, 
        \I5.AIR_WDATA_9l10r_net_1\, \I5.AIR_WDATA_9l9r_net_1\, 
        \I5.N_463\, \I5.N_480\, \I5.REG_12l431r_net_1\, 
        \I5.AIR_START_16_net_1\, \I4.N_1\, \I4.N_2\, \I4.N_4\, 
        \I4.N_5\, \I0.CLEARF1_i_net_1\, \I0.BNC_RESerr_1_net_1\, 
        \I0.EV_RESi_1_net_1\, \I2.N_2330_tz\, \I2.N_2328_tz\, 
        \I2.MIC_REG1_1_sqmuxa_0\, \I2.N_4327\, 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, \I2.un8_evread_1\, 
        \I2.MIC_REG1_0_sqmuxa_0_net_1\, \I2.TRAIL_MIS6_i_net_1\, 
        \I2.PIPE6_DT_il33r_net_1\, \I2.STATE3_il9r\, 
        \I2.TDCTRG_c_i_0\, \I2.BNC_ID_i_0l0r\, \I2.STATE5_nsl2r\, 
        \I2.L2ARR_n1_net_1\, \I2.N_4334\, \I2.N_4335\, 
        \I2.L2SERV_n1_net_1\, \I2.L2SERV_c1_net_1\, 
        \I2.ROFFSET_c2_net_1\, \I2.ROFFSET_c1_net_1\, 
        \I2.PIPE1_DT_42_1l29r\, \I2.N_4261\, \I2.N_3277\, 
        \I2.N_3351\, \I2.N_89_0\, \I2.N_64_0\, \I2.N_17\, 
        \I2.N_52\, \I2.N_52_0\, \I2.ADD_21x21_fast_I172_Y_0\, 
        \I2.ADD_21x21_fast_I172_Y_0_0\, \I2.N_85_0\, 
        \I2.un27_pipe5_dt0l0r\, \I2.un27_pipe5_dt1l0r\, 
        \I2.sram_empty_3_i_0_i\, \I2.un21_sram_empty_0_net_1\, 
        \I2.un21_sram_empty_1_net_1\, \I2.N_620\, \I2.N_621\, 
        \I2.N_623\, \I2.N_624\, \I2.N_627\, \I2.N_628\, 
        \I2.N_630\, \I2.N_631\, \I2.DTEST_FIFO_645_net_1\, 
        \I2.N_484\, \I2.N_483\, \I2.N_22_i_0\, \I2.N_4455\, 
        \I2.N_4459\, \I2.N_4460\, \I2.N_4454\, \I2.N_4456\, 
        \I2.N_4457\, \I2.N_4461\, \I2.N_4458\, 
        \I2.PIPE8_DT_21_i_0_il30r\, \I2.N_585\, \I2.N_584\, 
        \I2.N_583\, \I2.N_582\, \I2.N_581\, \I2.N_580\, 
        \I2.N_579\, \I2.N_578\, \I2.N_577\, \I2.N_576\, 
        \I2.N_575\, \I2.N_574\, \I2.N_573\, \I2.N_572\, 
        \I2.N_571\, \I2.N_570\, \I2.N_569\, \I2.N_568\, 
        \I2.N_567\, \I2.N_566\, \I2.un21_pipe5_dt_2_net_1\, 
        \I2.un21_pipe5_dt_0_net_1\, \I2.un21_pipe5_dt_1_net_1\, 
        \I2.un78_pipe5_dt_2_net_1\, \I2.un78_pipe5_dt_0_net_1\, 
        \I2.un78_pipe5_dt_1_net_1\, \I2.N_3019\, \I2.N_4673\, 
        \I2.N_4545\, \I2.N_219\, \I2.N_4542\, \I2.N_217\, 
        \I2.N_3890\, \I2.N_3882\, \I2.N_4676\, \I2.un1_STATE3\, 
        \I2.MIC_ERR_REGS_377_net_1\, \I2.MIC_ERR_REGS_376_net_1\, 
        \I2.MIC_ERR_REGS_375_net_1\, \I2.MIC_ERR_REGS_374_net_1\, 
        \I2.MIC_ERR_REGS_373_net_1\, \I2.MIC_ERR_REGS_372_net_1\, 
        \I2.MIC_ERR_REGS_371_net_1\, \I2.MIC_ERR_REGS_370_net_1\, 
        \I2.MIC_ERR_REGS_369_net_1\, \I2.MIC_ERR_REGS_368_net_1\, 
        \I2.MIC_ERR_REGS_367_net_1\, \I2.MIC_ERR_REGS_366_net_1\, 
        \I2.MIC_ERR_REGS_365_net_1\, \I2.MIC_ERR_REGS_364_net_1\, 
        \I2.MIC_ERR_REGS_363_net_1\, \I2.MIC_ERR_REGS_362_net_1\, 
        \I2.MIC_ERR_REGS_361_net_1\, \I2.MIC_ERR_REGS_360_net_1\, 
        \I2.MIC_ERR_REGS_359_net_1\, \I2.MIC_ERR_REGS_358_net_1\, 
        \I2.MIC_ERR_REGS_357_net_1\, \I2.MIC_ERR_REGS_356_net_1\, 
        \I2.MIC_ERR_REGS_355_net_1\, \I2.MIC_ERR_REGS_354_net_1\, 
        \I2.MIC_ERR_REGS_353_net_1\, \I2.MIC_ERR_REGS_352_net_1\, 
        \I2.MIC_ERR_REGS_351_net_1\, \I2.MIC_ERR_REGS_350_net_1\, 
        \I2.MIC_ERR_REGS_349_net_1\, \I2.MIC_ERR_REGS_348_net_1\, 
        \I2.MIC_ERR_REGS_347_net_1\, \I2.MIC_ERR_REGS_346_net_1\, 
        \I2.MIC_ERR_REGS_345_net_1\, \I2.MIC_ERR_REGS_344_net_1\, 
        \I2.MIC_ERR_REGS_343_net_1\, \I2.MIC_ERR_REGS_342_net_1\, 
        \I2.MIC_ERR_REGS_341_net_1\, \I2.MIC_ERR_REGS_340_net_1\, 
        \I2.MIC_ERR_REGS_339_net_1\, \I2.MIC_ERR_REGS_338_net_1\, 
        \I2.MIC_ERR_REGS_337_net_1\, \I2.MIC_ERR_REGS_336_net_1\, 
        \I2.MIC_ERR_REGS_335_net_1\, \I2.MIC_ERR_REGS_334_net_1\, 
        \I2.MIC_ERR_REGS_333_net_1\, \I2.MIC_ERR_REGS_332_net_1\, 
        \I2.MIC_ERR_REGS_331_net_1\, \I2.MIC_ERR_REGS_330_net_1\, 
        \I2.MIC_ERR_REGS_329_net_1\, \I2.W_ERR_WORDS_327_net_1\, 
        \I2.MIC_REG3_324_net_1\, \I2.MIC_REG3_323_net_1\, 
        \I2.MIC_REG3_322_net_1\, \I2.MIC_REG3_321_net_1\, 
        \I2.MIC_REG3_318_net_1\, \I2.MIC_REG3_317_net_1\, 
        \I2.MIC_REG2_316_net_1\, \I2.MIC_REG2_315_net_1\, 
        \I2.MIC_REG2_314_net_1\, \I2.MIC_REG2_313_net_1\, 
        \I2.MIC_REG2_310_net_1\, \I2.MIC_REG2_309_net_1\, 
        \I2.MIC_REG1_308_net_1\, \I2.MIC_REG1_307_net_1\, 
        \I2.MIC_REG1_306_net_1\, \I2.MIC_REG1_305_net_1\, 
        \I2.MIC_REG1_302_net_1\, \I2.MIC_REG1_301_net_1\, 
        \I2.END_TDC6_268_net_1\, \I2.END_EVNT6_267_net_1\, 
        \I2.BNCID_VECTrff_3_262_0_a2_0\, 
        \I2.BNCID_VECTrff_7_258_0_a2_0\, 
        \I2.BNCID_VECTrff_8_257_0_a2_0\, 
        \I2.BNCID_VECTrff_12_253_0_a2_0\, \I2.REG_1_n15_0_net_1\, 
        \I2.REG_1_n14_0_net_1\, \I2.REG_1_n13_0_net_1\, 
        \I2.REG_1_n12_0_net_1\, \I2.REG_1_n11_0_net_1\, 
        \I2.REG_1_n10_0_net_1\, \I2.REG_1_n9_0_net_1\, 
        \I2.REG_1_n8_0_net_1\, \I2.REG_1_n7_0_net_1\, 
        \I2.REG_1_n6_0_net_1\, \I2.REG_1_n5_0_net_1\, 
        \I2.REG_1_n4_0_net_1\, \I2.REG_1_n3_0_net_1\, \I2.N_119\, 
        \I2.N_3765\, \I2.N_3855\, \I2.N_3850\, \I2.N_3899\, 
        \I2.LSRAM_RADDRl2r_net_1\, \I2.LSRAM_RADDRl1r_net_1\, 
        \I2.LSRAM_RADDRl0r_net_1\, 
        \I2.DWACT_ADD_CI_0_partial_sum_2l0r\, 
        \I2.DWACT_ADD_CI_0_TMPl0r\, \I2.N_3547_i_i\, \I2.G_1_2\, 
        \I2.N_3539_i_i\, \I2.G_1_3\, \I2.N_3537_i_i\, \I2.G_1_4\, 
        \I2.ca_0_and2\, \I2.G_1_5\, \I2.SUB9_1l2r\, \I2.ca\, 
        \I3.TCNT1_i_0l0r\, CLEAR_STAT_i_0, NOEAD_c, 
        \I3.TCNT2_n1_net_1\, \I3.TCNT2_n2_net_1\, 
        \I3.TCNT4_388_net_1\, \I3.TCNT4_n1_net_1\, 
        \I3.TCNT4_c1_net_1\, \I3.TCNT3_379_net_1\, 
        \I3.TCNT3_n1_net_1\, \I3.TCNT3_n2_net_1\, \I3.un102_reg\, 
        \I3.N_1764\, \I3.N_1911\, \I3.N_291\, \I3.TCNT1_c1_net_1\, 
        \I3.TCNT1_n1_net_1\, \I3.N_558\, \I3.N_554\, \I3.N_555\, 
        \I3.N_551\, \I3.N_550\, \I3.N_552\, \I3.N_553\, 
        \I2.un3_tdcgda1_1_adt_net_821__net_1\, 
        \I2.un2_tdcgdb1_0_adt_net_830__net_1\, 
        \I2.N_3496_adt_net_926__net_1\, 
        \I2.N_4528_adt_net_1129__net_1\, 
        \I2.N_4529_adt_net_1136__net_1\, 
        \I2.N_4530_adt_net_1143__net_1\, 
        \I2.N_4531_adt_net_1150__net_1\, 
        \I2.N_4532_adt_net_1157__net_1\, 
        \I2.N_4533_adt_net_1164__net_1\, 
        \I2.N_4534_adt_net_1171__net_1\, 
        \I2.N_4535_adt_net_1178__net_1\, 
        \I3.N_243_4_adt_net_1290__net_1\, 
        \I5.sstate1_ns_el0r_adt_net_7898_\, 
        \REGl7r_adt_net_8466_\, 
        \I5.sstate1_ns_el3r_adt_net_9195_\, 
        \I5.SDAout_12_adt_net_9914_\, \REGl6r_adt_net_14043_\, 
        \I5.SENS_ADDR_1_sqmuxa_adt_net_14344_\, 
        \I4.un2_end_tdc_0_adt_net_15179_\, 
        \I4.un2_end_tdc_1_adt_net_15219_\, 
        \I4.END_FLUSH_2_adt_net_15635_\, \REGl18r_adt_net_15773_\, 
        \I0.TDC_RESi_1_adt_net_15858_\, 
        \I2.N_3760_adt_net_15913_\, \I2.N_3760_adt_net_15916_\, 
        \I2.N_2327_tz_adt_net_16395_\, 
        \I2.N_2329_tz_adt_net_16479_\, \I2.N_4524_adt_net_16635_\, 
        \I2.N_4273_adt_net_20927_\, \REGl1r_adt_net_21137_\, 
        \REGl2r_adt_net_21315_\, 
        \I2.un3_tdcgda1_1_adt_net_21664__net_1\, 
        \I2.un2_tdcgdb1_0_adt_net_21805__net_1\, 
        \I2.N_3457_ip_adt_net_23071_\, 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23152_\, 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23154_\, 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23155_\, 
        \I2.un21_sram_empty_NE_adt_net_24173_\, 
        \I2.N_118_i_1_adt_net_24217__net_1\, 
        \I3.N_203_adt_net_24459_\, 
        \I2.STATE3_0_sqmuxa_1_0_adt_net_24559_\, 
        \I2.ROFFSETe_0_adt_net_27184__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45405__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_45406__net_1\, 
        \I2.PIPE1_DT_42l29r_adt_net_45714_\, 
        \I2.un1_STATE1_39_6_i_adt_net_52470_\, 
        \REGl0r_adt_net_53773_\, \I2.N_128_adt_net_54290_\, 
        \I2.N_128_adt_net_54291_\, 
        \I2.N_2360_tz_tz_adt_net_54584_\, 
        \I2.N_108_0_adt_net_55153_\, \I2.N_222_adt_net_63455_\, 
        \I2.N_4551_adt_net_63758_\, \I2.N_4551_adt_net_63759_\, 
        \I2.N_3822_adt_net_64757_\, \I2.N_3822_adt_net_64759_\, 
        \I2.N_3822_adt_net_64761_\, \I2.N_3822_adt_net_64763_\, 
        \I2.N_3822_adt_net_64764_\, \I2.N_3822_adt_net_64765_\, 
        \I2.N_3822_adt_net_64766_\, \I2.N_4438_adt_net_66932_\, 
        \I2.N_4438_adt_net_66975_\, \I2.N_4439_adt_net_67071_\, 
        \I2.N_4439_adt_net_67114_\, \I2.N_4440_adt_net_67210_\, 
        \I2.N_4440_adt_net_67253_\, \I2.N_4442_adt_net_67433_\, 
        \I2.N_4442_adt_net_67476_\, \I2.N_4443_adt_net_67572_\, 
        \I2.N_4443_adt_net_67615_\, \I2.N_4444_adt_net_67711_\, 
        \I2.N_4444_adt_net_67754_\, \I2.N_4446_adt_net_67934_\, 
        \I2.N_4446_adt_net_67977_\, \I2.N_4447_adt_net_68073_\, 
        \I2.N_4447_adt_net_68116_\, \I2.N_4448_adt_net_68212_\, 
        \I2.N_4448_adt_net_68255_\, \I2.N_4450_adt_net_68435_\, 
        \I2.N_4450_adt_net_68478_\, \I2.N_4451_adt_net_68574_\, 
        \I2.N_4451_adt_net_68617_\, \I2.N_4452_adt_net_68713_\, 
        \I2.N_4452_adt_net_68756_\, \I2.N303_adt_net_69116_\, 
        \I2.N307_1_adt_net_69278_\, \I2.N309_adt_net_70030_\, 
        \I2.N305_adt_net_70150_\, \I2.N_3824_adt_net_90292_\, 
        \I2.N_3824_adt_net_90298_\, \I2.N_2989_adt_net_92422_\, 
        \I3.un6_tcnt1_adt_net_134941_\, 
        \I3.un6_tcnt1_adt_net_134944_\, 
        \I3.un10_tcnt2_adt_net_135286_\, 
        \I3.un10_tcnt2_adt_net_135288_\, 
        \I3.un10_tcnt2_adt_net_135290_\, 
        \I3.un10_tcnt2_adt_net_135291_\, 
        \I3.TCNT_n1_adt_net_137059_\, 
        \I3.TCNT_n2_adt_net_137234_\, 
        \I3.un1_STATE2_15_1_adt_net_147701__net_1\, 
        \I3.un1_STATE2_9_adt_net_154004_\, 
        \I3.N_544_adt_net_165558_\, 
        \I3.un7_ronly_0_a2_0_a3_adt_net_165586_\, 
        \I3.un12_tcnt3_adt_net_165616_\, 
        \I3.un12_tcnt3_adt_net_165618_\, 
        \I3.un12_tcnt3_adt_net_165620_\, 
        \I3.un12_tcnt3_adt_net_165621_\, 
        \I3.un15_tcnt4_adt_net_165650_\, 
        \I3.un15_tcnt4_adt_net_165652_\, 
        \I3.N_545_adt_net_165682_\, \I3.N_586_adt_net_165970_\, 
        \I3.un60_reg_ads_3_adt_net_166295_\, 
        \I2.N_107_adt_net_256840_\, \I2.N_107_adt_net_276024_\, 
        \I3.N_1309_i_net_1\, \I3.TCNT3_c2\, \I3.TCNT2_c2\, 
        \I5.SCL_1_i_a2_0_1_net_1\, \I5.N_479\, \I5.N_67\, 
        \I4.bcnt_7_net_1\, \I4.bcnt_6_net_1\, \I4.N_3\, \I4.N_6\, 
        \I4.FLUSH_1_sqmuxa\, \I4.un2_end_tdc_1_net_1\, 
        \I4.un2_end_tdc_0_net_1\, \I2.N_2329_tz\, \I2.N_4328\, 
        \I2.N_565_0\, \I2.DWACT_ADD_CI_0_g_array_1l0r\, 
        \I2.DWACT_ADD_CI_0_g_array_12l0r\, \I2.L1AF2_i_net_1\, 
        \I2.L2RF2_i_net_1\, \I2.N_4462\, \I2.EVNT_NUM_n2_tz_i\, 
        \I2.EVNT_NUM_c2_net_1\, \I2.L2ARR_n2_net_1\, 
        \I2.L2ARR_c2_net_1\, \I2.N_4336\, \I2.N_279\, \I2.N_317\, 
        \I2.N_189\, \I2.N_186\, \I2.L2SERV_n2_net_1\, 
        \I2.L2SERV_c2_net_1\, \I2.ROFFSET_n2_tz_i\, 
        \I2.ROFFSET_n3_tz_i\, \I2.ROFFSET_c3_net_1\, \I2.N_4182\, 
        \I2.PIPE1_DT_12l30r_net_1\, \I2.PIPE1_DT_30l30r_net_1\, 
        \I2.PIPE1_DT_12l20r_net_1\, \I2.PIPE1_DT_30l20r_net_1\, 
        \I2.PIPE1_DT_12l19r_net_1\, \I2.PIPE1_DT_30l19r_net_1\, 
        \I2.PIPE1_DT_12l18r_net_1\, \I2.PIPE1_DT_30l18r_net_1\, 
        \I2.PIPE1_DT_12l17r_net_1\, \I2.PIPE1_DT_30l17r_net_1\, 
        \I2.PIPE1_DT_12l16r_net_1\, \I2.PIPE1_DT_30l16r_net_1\, 
        \I2.PIPE1_DT_30l15r_net_1\, \I2.PIPE1_DT_12l15r_net_1\, 
        \I2.PIPE1_DT_30l14r_net_1\, \I2.PIPE1_DT_12l14r_net_1\, 
        \I2.PIPE1_DT_30l13r_net_1\, \I2.PIPE1_DT_12l13r_net_1\, 
        \I2.PIPE1_DT_30l12r_net_1\, \I2.PIPE1_DT_12l12r_net_1\, 
        \I2.PIPE1_DT_30l11r_net_1\, \I2.PIPE1_DT_12l11r_net_1\, 
        \I2.PIPE1_DT_30l10r_net_1\, \I2.PIPE1_DT_12l10r_net_1\, 
        \I2.PIPE1_DT_30l9r_net_1\, \I2.PIPE1_DT_12l9r_net_1\, 
        \I2.PIPE1_DT_30l8r_net_1\, \I2.PIPE1_DT_12l8r_net_1\, 
        \I2.PIPE1_DT_30l7r_net_1\, \I2.PIPE1_DT_12l7r_net_1\, 
        \I2.PIPE1_DT_30l6r_net_1\, \I2.PIPE1_DT_12l6r_net_1\, 
        \I2.PIPE1_DT_30l5r_net_1\, \I2.PIPE1_DT_12l5r_net_1\, 
        \I2.PIPE1_DT_30l4r_net_1\, \I2.PIPE1_DT_12l4r_net_1\, 
        \I2.PIPE1_DT_12l3r_net_1\, \I2.PIPE1_DT_30l3r_net_1\, 
        \I2.PIPE1_DT_12l2r_net_1\, \I2.PIPE1_DT_30l2r_net_1\, 
        \I2.PIPE1_DT_30l1r_net_1\, \I2.PIPE1_DT_12l1r_net_1\, 
        \I2.PIPE1_DT_12l0r_net_1\, \I2.PIPE1_DT_30l0r_net_1\, 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\, 
        \I2.N_80\, \I2.N_112_2\, \I2.N_95\, \I2.N_108\, 
        \I2.N_128\, \I2.N_95_0\, \I2.N_139_0\, \I2.N_140_0\, 
        \I2.N_84_0\, \I2.ADD_21x21_fast_I174_Y_0\, 
        \I2.ADD_21x21_fast_I174_Y_0_0\, \I2.N_28_0\, 
        \I2.ADD_21x21_fast_I173_Y_0\, 
        \I2.ADD_21x21_fast_I173_Y_0_0\, \I2.N357\, \I2.N357_0\, 
        \I2.ADD_21x21_fast_I171_Y_0\, 
        \I2.ADD_21x21_fast_I171_Y_0_0\, \I2.N_3870\, 
        \I2.un21_sram_empty_NE_net_1\, \I2.N_629\, \I2.N_632\, 
        \I2.N_3822\, \I2.N_26\, \I2.N_4468\, \I2.N_4467\, 
        \I2.N_4466\, \I2.N_4465\, \I2.L2AS_net_1\, 
        \I2.ADD_18x18_fast_I147_Y_0\, \I2.N241\, 
        \I2.ADD_18x18_fast_I145_Y_0\, \I2.N238\, 
        \I2.ADD_18x18_fast_I144_Y_0\, \I2.N235\, 
        \I2.ADD_18x18_fast_I143_Y_0\, \I2.N232\, 
        \I2.ADD_18x18_fast_I142_Y_0\, 
        \I2.ADD_18x18_fast_I141_Y_0\, \I2.N225\, \I2.SUB9_1l3r\, 
        \I2.N_4401\, \I2.un21_pipe5_dt_3_net_1\, 
        \I2.un78_pipe5_dt_3_net_1\, \I2.STATE3_0_sqmuxa_1_0\, 
        \I2.N_3016\, \I2.N_4551\, \I2.N_2327_tz\, 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1\, \I2.TOKINBi_326_net_1\, 
        \I2.MIC_REG3_319_net_1\, \I2.MIC_REG2_311_net_1\, 
        \I2.MIC_REG1_303_net_1\, \I2.BNCID_VECTrff_0_265_0_net_1\, 
        \I2.BNCID_VECTrff_1_264_0_net_1\, 
        \I2.BNCID_VECTrff_2_263_0_net_1\, 
        \I2.BNCID_VECTrff_3_262_0_net_1\, 
        \I2.BNCID_VECTrff_4_261_0_net_1\, 
        \I2.BNCID_VECTrff_5_260_0_net_1\, 
        \I2.BNCID_VECTrff_6_259_0_net_1\, 
        \I2.BNCID_VECTrff_7_258_0_net_1\, 
        \I2.BNCID_VECTrff_8_257_0_net_1\, 
        \I2.BNCID_VECTrff_9_256_0_net_1\, 
        \I2.BNCID_VECTrff_10_255_0_net_1\, 
        \I2.BNCID_VECTrff_11_254_0_net_1\, 
        \I2.BNCID_VECTrff_12_253_0_net_1\, 
        \I2.BNCID_VECTrff_13_252_0_net_1\, 
        \I2.BNCID_VECTrff_14_251_0_net_1\, 
        \I2.BNCID_VECTrff_15_250_0_net_1\, \I2.N_121\, 
        \I2.REG_1_n0_0_net_1\, \I2.N_3858\, \I2.N_177\, 
        \I2.TRGARR_3l2r\, \I2.TRGARR_3l3r\, \I2.TRGARR_3l1r\, 
        \I3.N_1910_0\, NOEAD_c_i_0, \I3.TCNT2_394_net_1\, 
        \I3.TCNT2_n3_net_1\, \I3.TCNT4_387_net_1\, 
        \I3.TCNT4_n2_net_1\, \I3.TCNT4_c2_net_1\, 
        \I3.TCNT3_378_net_1\, \I3.TCNT3_377_net_1\, 
        \I3.TCNT3_n3_net_1\, REGl6r, REG_i_il5r, REGl2r, REGl1r, 
        REGl0r, REGl18r, \I3.N_1904\, \I3.N_1912\, \I3.N_268\, 
        \I3.un22_bltcyc\, \I3.TCNT1_c2_net_1\, 
        \I3.TCNT1_n2_net_1\, \I3.un231_reg_ads_1\, 
        \I3.un41_reg_ads_0_a2_3_a3_0\, \I3.un47_reg_ads_1\, 
        \I3.N_634\, \I3.un60_reg_ads_3\, \I3.N_562\, \I3.N_578\, 
        \I3.N_581\, \I3.N_544\, \I3.un6_tcnt1_net_1\, 
        \I2.N_3_0_adt_net_1070__net_1\, 
        \I2.N_118_i_1_adt_net_1122__net_1\, 
        \I2.N_3877_adt_net_4723_\, \I2.N_3877_adt_net_4725_\, 
        \I2.N_3876_adt_net_4861_\, \I5.N_71_adt_net_9287_\, 
        \I4.STATE1_nsl2r_adt_net_15265_\, 
        \I2.N_4524_adt_net_16596_\, \I2.N_4524_adt_net_16740_\, 
        \I2.N_4646_1_adt_net_19637_Ra1__net_1\, 
        \I2.N_4431_adt_net_22416_\, \I2.N_4424_adt_net_22594_\, 
        \REGl29r_adt_net_35602_\, \REGl28r_adt_net_36082_\, 
        \I2.N_108_adt_net_54237_\, \I2.N_74_i_0_i_adt_net_54331_\, 
        \I2.N_70_adt_net_54406__net_1\, 
        \I2.N_128_0_adt_net_55238_\, \I2.N_29_i_0_adt_net_59529_\, 
        \I2.N531_0_adt_net_60100_\, \I2.N_3866_adt_net_61361_\, 
        \I2.N_3824_adt_net_90281_\, \I2.N_3830_adt_net_101622_\, 
        \reg_il0r_adt_net_105174_\, \I3.TCNT_n3_adt_net_137329_\, 
        \I3.un1_STATE1_13_1_adt_net_137896__net_1\, 
        \I3.un7_ronly_0_a2_0_a3_adt_net_165588_\, 
        \I3.un221_reg_ads_0_a2_0_a3_adt_net_165933_\, 
        \I3.un68_reg_ads_0_a2_3_a3_adt_net_166224_\, 
        \I2.N_70_adt_net_255801__net_1\, 
        \I2.N_70_adt_net_255802__net_1\, 
        \I2.N_114_adt_net_275711_\, \I2.N_114_adt_net_275800_\, 
        \I2.N_107_adt_net_256839_\, \I2.N_107_0_adt_net_320361_\, 
        \I2.N_107_0_adt_net_320362_\, \I2.N_107_0\, 
        \I2.N525_adt_net_336000_\, \I3.TCNT3_c3\, \I3.TCNT2_c3\, 
        \I5.N_100\, \I5.N_98\, \I5.N_96\, \I5.N_95\, 
        \I5.sstate1se_12_i_net_1\, \I5.sstate1_ns_el9r\, 
        \I5.sstate1_ns_el6r\, \I5.N_77\, \I5.N_70\, 
        \I4.bcnt_5_net_1\, \I4.un1_lead_flag_1\, \I4.I_5\, 
        \I2.N_4329\, \I2.EVNT_NUM_n3_tz_i\, 
        \I2.EVNT_NUM_c3_net_1\, \I2.L2ARR_n3_net_1\, \I2.N_316_i\, 
        \I2.N_4669\, \I2.L2SERV_n3_net_1\, \I2.ROFFSET_n4_tz_i\, 
        \I2.ROFFSET_c4_net_1\, 
        \I2.DTO_16_1_iv_0_a2_4tt_18_m2_0_a2_net_1\, 
        \I2.DTO_16_1_iv_0_o2_2tt_21_N_8\, \I2.N307\, \I2.N_8\, 
        \I2.N_57\, \I2.N_20_i_0\, \I2.N_92_0\, \I2.N_53\, 
        \I2.N_75\, \I2.N_53_0\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_i_1\, \I2.N_70\, 
        \I2.N_59\, \I2.N_66\, 
        \I2.ADD_21x21_fast_I140_Y_0_a2_0_0_0\, \I2.N_16\, 
        \I2.N_13_1\, \I2.N_16_0\, \I2.N_45_0\, \I2.N_128_0\, 
        \I2.ADD_21x21_fast_I121_Y_i_a3_0_i\, \I2.N_2360_tz_tz\, 
        \I2.N_2358_tz_tz\, \I2.un27_pipe5_dt0l2r\, 
        \I2.un27_pipe5_dt1l2r\, \I2.un27_pipe5_dt0l1r\, 
        \I2.un27_pipe5_dt1l1r\, \I2.N_626\, 
        \I2.PIPE10_DT_17_i_0l20r_net_1\, 
        \I2.PIPE10_DT_17_i_0l19r_net_1\, 
        \I2.PIPE10_DT_17_i_0l18r_net_1\, 
        \I2.PIPE10_DT_17_i_0l17r_net_1\, 
        \I2.PIPE10_DT_17_i_0l16r_net_1\, 
        \I2.PIPE10_DT_17_i_0l15r_net_1\, 
        \I2.PIPE10_DT_17_i_0l14r_net_1\, 
        \I2.PIPE10_DT_17_i_0l13r_net_1\, \I2.N_4397\, \I2.N_4402\, 
        \I2.N_4398\, \I2.N_4403\, \I2.un21_pipe5_dt_4_net_1\, 
        \I2.un78_pipe5_dt_4_net_1\, \I2.EVRDYi_496_net_1\, 
        \I2.N_4526\, \I2.TOKINAi_325_net_1\, 
        \I2.BNCID_VECTwa12_1_net_1\, \I2.BNCID_VECTwa13_1_net_1\, 
        \I2.BNCID_VECTwa14_1_net_1\, \I2.BNCID_VECTwa15_1_net_1\, 
        \I2.N_122\, \I2.N_3860\, REGl29r, REGl28r, \I2.N_4431\, 
        \I2.N_4424\, \I2.N_3876\, \I2.N_3877\, reg_il0r, 
        \I3.un10_tcnt2_i_net_1\, NOE16W_c, \I3.TCNT2_396_net_1\, 
        \I3.TCNT2_395_net_1\, \I3.TCNT2_393_net_1\, 
        \I3.TCNT2_n4_net_1\, \I3.TCNT4_386_net_1\, 
        \I3.TCNT4_n3_net_1\, \I3.TCNT3_376_net_1\, 
        \I3.TCNT3_n4_net_1\, \I3.N_1919\, \I3.N_1409\, 
        \I3.TCNT1_c3_net_1\, \I3.TCNT1_n3_net_1\, 
        \I3.un7_ronly_0_a2_0_a3_net_1\, \I3.un10_tcnt2_net_1\, 
        \I3.un227_reg_ads_2\, \I3.N_545\, 
        \I2.N_163_adt_net_1241__net_1\, 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, 
        \I5.sstate1se_12_i_adt_net_8689_\, 
        \I5.sstate1_ns_el8r_adt_net_8886_\, 
        \I5.sstate1_ns_el1r_adt_net_9246_\, 
        \I2.N_4524_adt_net_16701_\, 
        \I2.N_4646_1_adt_net_19635__net_1\, 
        \I2.STATE3_nsl12r_adt_net_24672_\, 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26947_\, 
        \I2.DTO_16_1_iv_0_o2_2tt_21_m3_adt_net_27978_\, 
        \I2.N519_adt_net_54631_\, \I2.N_75_adt_net_54671_\, 
        \I2.N_152_i_adt_net_54710__net_1\, 
        \I2.N_33_adt_net_55020_\, \I2.N_74_adt_net_55281_\, 
        \I2.N_152_i_0_adt_net_55693__net_1\, 
        \I2.N507_adt_net_56251__net_1\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_2_adt_net_56513_\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_N_6_i_adt_net_56543_\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_N_6_i_adt_net_56545_\, 
        \I2.N_100_adt_net_58424_\, 
        \I2.ADD_21x21_fast_I138_Y_0_0_adt_net_58475_\, 
        \I2.N_100_0_adt_net_58633_\, 
        \I2.ADD_21x21_fast_I138_Y_0_0_0_adt_net_58684_\, 
        \I2.un1_NWPIPE7_2_adt_net_73604_\, 
        \I2.un1_NWPIPE7_2_adt_net_73606_\, 
        \I2.N_4397_adt_net_90034_\, \I2.N_4398_adt_net_90118_\, 
        \I2.N_107\, \I2.N507_adt_net_258084__net_1\, 
        \I2.N507_adt_net_56246__net_1\, 
        \I2.N_45_1_adt_net_271427_\, \I2.N_45_1\, 
        \I2.N507_adt_net_283110__net_1\, 
        \I2.N525_0_adt_net_318487_\, \I2.N525_0_adt_net_318530_\, 
        \I2.N525_0_adt_net_58018_\, \I2.N522_0_adt_net_329169_\, 
        \I2.N522_0_adt_net_329219_\, \I2.N525_adt_net_335996_\, 
        \I2.N525_adt_net_57834_\, \I2.N507_adt_net_347769__net_1\, 
        \I2.N507_adt_net_347770__net_1\, 
        \I2.N507_adt_net_347771__net_1\, 
        \I2.N522_0_adt_net_384644_\, \I2.N_96_0_adt_net_469923_\, 
        \I2.N_96_adt_net_481750_\, \I2.N_82_adt_net_496796_\, 
        \I2.N_152_i_0_adt_net_502546_\, 
        \I2.N_40_adt_net_589803__net_1\, 
        \I2.N_40_adt_net_589963__net_1\, 
        \I2.N_40_adt_net_1100__net_1\, 
        \I2.N_147_0_adt_net_604832_\, \I3.TCNT3_c4\, 
        \I3.TCNT2_c4\, \I5.sstate1se_3_i_net_1\, 
        \I5.sstate1_ns_el3r\, \I4.LSRAM_FL_RADDR_0_sqmuxa\, 
        \I4.bcnt_8_net_1\, \I4.N_4_0\, \I4.I_9\, \I2.dataout_0\, 
        \I2.EVNT_NUM_n4_tz_i\, \I2.EVNT_NUM_c4_net_1\, \I2.N_319\, 
        \I2.ROFFSET_n5_tz_i\, \I2.ROFFSET_c5_net_1\, 
        \I2.DTO_16_1_iv_0_o2_2tt_21_m3_net_1\, 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m3_net_1\, 
        \I2.ADD_21x21_fast_I190_Y_0\, 
        \I2.ADD_21x21_fast_I189_Y_0\, \I2.N_63\, \I2.N313\, 
        \I2.ADD_21x21_fast_I188_Y_0\, 
        \I2.ADD_21x21_fast_I187_Y_0\, \I2.N_65\, 
        \I2.ADD_21x21_fast_I186_Y_0\, 
        \I2.ADD_21x21_fast_I185_Y_0\, \I2.N_57_0\, 
        \I2.ADD_21x21_fast_I184_Y_0\, \I2.N_20_i\, \I2.N_92\, 
        \I2.ADD_21x21_fast_I183_Y_0\, 
        \I2.ADD_21x21_fast_I182_Y_0\, \I2.N_91\, 
        \I2.ADD_21x21_fast_I181_Y_0\, \I2.N_74_i_0_i\, \I2.N_74\, 
        \I2.N_70_0\, \I2.N_59_0\, \I2.ADD_21x21_fast_I180_Y_0\, 
        \I2.N_13_0\, \I2.ADD_21x21_fast_I179_Y_0\, \I2.N525\, 
        \I2.ADD_21x21_fast_I178_Y_0\, 
        \I2.ADD_21x21_fast_I177_Y_0\, \I2.N_140\, 
        \I2.ADD_21x21_fast_I176_Y_0\, \I2.N_158_0\, 
        \I2.ADD_21x21_fast_I121_Y_i_a3_0_i_0\, \I2.N_29_i_0\, 
        \I2.ADD_21x21_fast_I175_Y_0\, \I2.N394\, \I2.N_93_0\, 
        \I2.un27_pipe5_dt0l3r\, \I2.un27_pipe5_dt1l3r\, 
        \I2.N_1071\, \I2.N_1070\, \I2.N_1069\, 
        \I2.un28_sram_empty\, \I2.un1_STATE3_8\, \I2.N_124\, 
        \I2.ADE_4l15r_net_1\, \I2.ADE_4l14r_net_1\, 
        \I2.ADE_4l13r_net_1\, \I2.ADE_4l12r_net_1\, 
        \I2.DWACT_ADD_CI_0_partial_sum_1l0r\, \I3.N_57_i_0_0\, 
        NOE32W_c, \I3.TCNT2_392_net_1\, \I3.TCNT2_n5_net_1\, 
        \I3.TCNT4_385_net_1\, \I3.N_263_i\, \I3.TCNT3_375_net_1\, 
        \I3.TCNT3_n5_net_1\, \I3.TCNT1_c4_net_1\, 
        \I3.TCNT1_n4_net_1\, \I3.un12_tcnt3_net_1\, 
        \I3.un68_reg_ads_0_a2_3_a3_net_1\, \I3.N_546\, 
        \I3.un41_reg_ads_2\, \I2.N_140_0_adt_net_947__net_1\, 
        \I2.N_3836_i_0_adt_net_2390__net_1\, 
        \I2.N_152_i_adt_net_4109__net_1\, 
        \I2.N_152_i_0_adt_net_4117__net_1\, 
        \I5.SDAnoe_8_adt_net_9736_\, \I2.N_152_i_adt_net_54890_\, 
        \I2.N_41_adt_net_54991_\, \I2.N_33_adt_net_55021_\, 
        \I2.N_163_0_adt_net_55087_\, \I2.N_139_0_adt_net_55124_\, 
        \I2.N519_0_adt_net_55614_\, \I2.N_152_i_0_adt_net_55873_\, 
        \I2.N498_adt_net_56484_\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_2_adt_net_56515_\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_2_i_adt_net_56602_\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_4_adt_net_56769_\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_adt_net_56806_\, 
        \I2.N_86_i_adt_net_57123_\, \I2.N_40_adt_net_57971_\, 
        \I2.N525_0_adt_net_58015_\, \I2.N_96_0_adt_net_58152_\, 
        \I2.N_40_0_adt_net_58199_\, \I2.N_3_adt_net_59496_\, 
        \I2.N531_adt_net_59960_\, \I2.N531_0_adt_net_60059_\, 
        \I2.un1_NWPIPE7_2_adt_net_73600_\, \I2.N522_0\, \I2.N_96\, 
        \I2.N_82\, \I2.N_152_i_0_adt_net_502321_\, 
        \I2.N_152_i_0_adt_net_502367_\, 
        \I2.N_152_i_0_adt_net_502543_\, 
        \I2.N_152_i_0_adt_net_502544_\, 
        \I2.N_40_0_adt_net_577252_\, \I2.N_40_0_adt_net_577293_\, 
        \I2.N_40_0_adt_net_577295_\, \I2.N_147_0_adt_net_604875_\, 
        \I2.N_152_i_0_adt_net_610537_\, 
        \I2.N_152_i_0_adt_net_610542_\, 
        \I2.N_152_i_0_adt_net_610543_\, \N_1.I3.TCNT3_c5\, 
        \N_1.I3.TCNT2_c5\, \I4.LSRAM_FL_RADDR_0_sqmuxa_1\, 
        \I4.N_48_3\, \I4.bcnt_3l0r_net_1\, \I4.I_13_0\, 
        \I2.DWACT_ADD_CI_0_g_array_1_0l0r\, 
        \I2.DWACT_ADD_CI_0_g_array_12_0l0r\, \I2.NOESRAME_c_i_0\, 
        \I2.EVNT_NUM_n5_tz_i\, \I2.EVNT_NUM_c5_net_1\, 
        \I2.ROFFSET_c6_net_1\, \I2.ADD_21x21_fast_I190_Y_0_0\, 
        \I2.N_103\, \I2.ADD_21x21_fast_I189_Y_0_0\, \I2.N_63_0\, 
        \I2.N_33\, \I2.ADD_21x21_fast_I188_Y_0_0\, \I2.N_163_0\, 
        \I2.N502_i\, \I2.ADD_21x21_fast_I187_Y_0_0\, 
        \I2.un27_pipe5_dt0l16r\, \I2.ADD_21x21_fast_I186_Y_0_0\, 
        \I2.N_32_0\, \I2.N_8_0\, \I2.N507\, 
        \I2.ADD_21x21_fast_I185_Y_0_0\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_1_i\, \I2.N_40\, 
        \I2.ADD_21x21_fast_I184_Y_0_0\, \I2.N_40_0\, 
        \I2.ADD_21x21_fast_I138_Y_0_0\, \I2.N_100\, 
        \I2.ADD_21x21_fast_I183_Y_0_0\, 
        \I2.ADD_21x21_fast_I138_Y_0_0_0\, \I2.N_100_0\, 
        \I2.N_42_0\, \I2.ADD_21x21_fast_I182_Y_0_0\, \I2.N_91_0\, 
        \I2.N519\, \I2.ADD_21x21_fast_I181_Y_0_0\, \I2.N519_0\, 
        \I2.N522\, \I2.ADD_21x21_fast_I180_Y_0_0\, 
        \I2.un27_pipe5_dt0l9r\, \I2.ADD_21x21_fast_I179_Y_0_0\, 
        \I2.N525_0\, \I2.ADD_21x21_fast_I178_Y_0_0\, 
        \I2.ADD_21x21_fast_I177_Y_0_0\, \I2.N_61_0\, \I2.N_29_i\, 
        \I2.ADD_21x21_fast_I176_Y_0_0\, \I2.N_31_0\, \I2.N537_i\, 
        \I2.ADD_21x21_fast_I175_Y_0_0\, \I2.N537_i_0\, 
        \I2.un27_pipe5_dt0l4r\, \I2.N394_0\, \I2.N_1072\, 
        \I2.dataout_1\, \I2.N_126\, \I2.ADO_3l15r_net_1\, 
        \I2.ADO_3l14r_net_1\, \I2.ADO_3l13r_net_1\, 
        \I2.ADO_3l12r_net_1\, \I2.TRGSERV_2l2r\, 
        \I2.TRGSERV_2l3r\, \I2.TRGSERV_2l1r\, 
        \I3.TCNT2_391_net_1\, \I3.TCNT3_374_net_1\, 
        \I3.TCNT1_n5_net_1\, \I3.un15_tcnt4_net_1\, 
        \I3.un224_reg_ads_0_a2_3_a3_net_1\, \I3.N_632\, 
        \I3.un41_reg_ads_0_a2_3_a3_net_1\, \I3.N_573\, 
        \I3.un10_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un2_reg_ads_0_a2_0_a3_net_1\, 
        \I2.PIPE5_DT_6l28r_adt_net_53820_\, 
        \I2.N_152_i_adt_net_54886_\, \I2.N_41_adt_net_54984_\, 
        \I2.N_41_0_adt_net_55921_\, \I2.N_41_0_adt_net_55923_\, 
        \I2.N_33_0_adt_net_55957_\, \I2.N_33_0_adt_net_55958_\, 
        \I2.N498_0_adt_net_56939_\, \I2.N498_0_adt_net_56940_\, 
        \I2.N513_i_adt_net_58503_\, \I2.N513_i_0_adt_net_58712_\, 
        \I2.N_3_0_adt_net_59703_\, \I2.N502_i_0_adt_net_490246_\, 
        \I2.N502_i_0_adt_net_490392_\, 
        \I2.N502_i_0_adt_net_490398_\, 
        \I2.N498_0_adt_net_598283_\, \I2.N498_0_adt_net_598321_\, 
        \N_1.I3.TCNT3_n6\, \N_1.I3.TCNT3_c6\, \N_1.I3.TCNT2_n6\, 
        \N_1.I3.TCNT2_c6\, \I4.LSRAM_FL_RADDR_11\, 
        \I4.LSRAM_FL_RADDR_10\, \I4.LSRAM_FL_RADDR_9\, 
        \I4.bcnt_3l3r_net_1\, \I2.EVNT_NUM_n6_tz_i\, 
        \I2.EVNT_NUM_c6_net_1\, \I2.BNCID_VECTra14_1_net_1\, 
        \I2.BNCID_VECTra15_1_net_1\, \I2.BNCID_VECTra12_1_net_1\, 
        \I2.BNCID_VECTra13_1_net_1\, \I2.N_41\, \I2.N_41_0\, 
        \I2.N498\, \I2.N498_0\, \I2.N_86_i\, \I2.N_33_0\, 
        \I2.N_86_i_0\, \I2.un27_pipe5_dt0l17r\, 
        \I2.un27_pipe5_dt0l15r\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4\, 
        \I2.un27_pipe5_dt0l14r\, \I2.un27_pipe5_dt1l14r\, 
        \I2.N513_i\, \I2.N513_i_0\, \I2.un27_pipe5_dt0l12r\, 
        \I2.N_42_1\, \I2.un27_pipe5_dt0l11r\, 
        \I2.un27_pipe5_dt1l11r\, \I2.un27_pipe5_dt0l10r\, 
        \I2.un27_pipe5_dt1l10r\, \I2.un27_pipe5_dt1l9r\, 
        \I2.N_3_0\, \I2.N531\, \I2.N531_0\, \I2.N_31\, 
        \I2.un27_pipe5_dt1l6r\, \I2.un27_pipe5_dt0l5r\, 
        \I2.un27_pipe5_dt1l5r\, \I2.un27_pipe5_dt1l4r\, 
        \I2.N_4595\, \I3.N_548\, \I2.N502_i_0\, TCNT3_373, 
        \N_1.I3.TCNT3_n7\, TCNT2_390, \N_1.I3.TCNT2_n7\, 
        \I2.EVNT_NUM_n7_tz_i\, \I2.EVNT_NUM_c7_net_1\, \I2.N_1_1\, 
        \I2.N_1_1_0\, \I2.un27_pipe5_dt0l19r\, 
        \I2.un27_pipe5_dt1l19r\, \I2.N_2\, \I2.N_2_0\, 
        \I2.un27_pipe5_dt1l17r\, \I2.N_82_0\, 
        \I2.un27_pipe5_dt1l15r\, \I2.N_1083\, 
        \I2.un27_pipe5_dt0l13r\, \I2.un27_pipe5_dt1l13r\, 
        \I2.un27_pipe5_dt1l12r\, \I2.N_1080\, \I2.N_1079\, 
        \I2.N_1078\, \I2.N_3\, \I2.un27_pipe5_dt1l8r\, 
        \I2.un27_pipe5_dt0l7r\, \I2.un27_pipe5_dt1l7r\, 
        \I2.un27_pipe5_dt0l6r\, \I2.N_1074\, \I2.N_1073\, 
        TCNT3_372, TCNT2_389, \I2.EVNT_NUM_n8_tz_i\, 
        \I2.EVNT_NUM_c8_net_1\, \I2.un27_pipe5_dt0l20r\, 
        \I2.un27_pipe5_dt1l20r\, \I2.un27_pipe5_dt0l18r\, 
        \I2.un27_pipe5_dt1l18r\, \I2.un27_pipe5_dt1l16r\, 
        \I2.N_1084\, \I2.N_1082\, \I2.N_1081\, 
        \I2.un27_pipe5_dt0l8r\, \I2.N_1076\, \I2.N_1075\, 
        \I1.FBOUTl7r_net_1\, \FBOUTl6r\, \FBOUTl5r\, \FBOUTl4r\, 
        \FBOUTl3r\, \FBOUTl2r\, \FBOUTl1r\, 
        \I2.N_3843_adt_net_101094_\, \I2.N_1085\, \I2.N_1077\, 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r_adt_net_107356_\, 
        \I1.un1_sbyte13_i_i_i_1_adt_net_108180_\, 
        \I2.N346_adt_net_69448__net_1\, 
        \I1.N_628_adt_net_107115_\, \I1.N_366\, \I2.N309\, 
        \I2.N307_1\, \I2.SUB9_1l4r\, \I1.N_329\, 
        \I1.SBYTE_58_net_1\, \I2.N311\, \I2.N310\, 
        \I2.ADD_18x18_fast_I146_Y_0\, \I2.N301_1_adt_net_70232_\, 
        \I2.N244\, \I2.N305\, \I2.N_4244\, \I2.N_4245\, 
        \I2.N_4246\, \I2.N_4247\, \I2.N_4248\, \I2.N_4249\, 
        \I2.N_4250\, \I2.N_4251\, \I2.N_4252\, \I2.N_4253\, 
        \I2.N_4254\, \I2.N_4255\, \I2.DTE_2_1_0l4r_net_1\, 
        \I2.DTE_21_1l4r\, \I2.DTE_2_1_0l5r_net_1\, 
        \I2.DTE_2_1_0l6r_net_1\, \I2.DTE_21_1l6r\, 
        \I2.DTE_2_1_0l7r_net_1\, \I2.DTE_21_1l7r\, 
        \I2.DTE_2_1_0l8r_net_1\, \I2.DTE_21_1l8r\, 
        \I2.DTE_2_1_0l9r_net_1\, \I2.DTE_21_1l9r\, 
        \I2.DTE_2_1_0l10r_net_1\, \I2.DTE_21_1l10r\, 
        \I2.DTE_2_1_0l11r_net_1\, \I2.DTE_21_1l12r\, 
        \I2.DTE_21_1l13r\, \I2.DTE_21_1l16r\, \I2.DTE_21_1l19r\, 
        \I2.DTE_21_1l21r\, \I2.DTE_21_1l22r_adt_net_37395_\, 
        \I2.DTE_21_1l23r_adt_net_37285_\, 
        \I2.DTE_21_1l24r_adt_net_37175_\, \I2.N_4644\, 
        \I2.DTE_21_1l26r\, \I2.DTE_21_1l27r\, \I2.DTE_21_1l28r\, 
        \I2.DTE_21_1l17r\, \I2.DTE_21_1_iv_0_18_N_8_i_0\, 
        \I2.DTO_16_1l4r\, \I2.DTO_16_1l6r\, \I2.DTO_16_1l7r\, 
        \I2.DTO_16_1l8r\, \I2.DTO_16_1l9r\, \I2.DTO_16_1l10r\, 
        \I2.DTO_16_1l12r\, \I2.DTO_16_1l13r\, \I2.DTO_16_1l16r\, 
        \I2.DTO_16_1l17r\, \I2.DTO_16_1l18r\, \I2.DTO_16_1l19r\, 
        \I2.DTO_16_1l21r\, \I2.DTO_16_1l22r\, \I2.DTO_16_1l23r\, 
        \I2.DTO_16_1l24r\, \I2.DTO_16_1l25r\, \I2.DTO_16_1l26r\, 
        \I2.DTO_16_1l27r\, \I2.PIPE10_DT_17l29r_adt_net_64809_\, 
        \I1.N_358\, \I2.N_3799\, \I2.N_3800\, \I2.N_3801\, 
        \I2.N_3802\, \I2.N_3803\, \I2.N_3804\, \I2.N_3805\, 
        \I2.N_3806\, \I3.un57_reg_ads_0_a2_3_a3_net_1\, 
        \I3.un60_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un221_reg_ads_0_a2_0_a3_net_1\, 
        \I1.N_77_adt_net_109270_\, 
        \I3.un227_reg_ads_0_a2_3_a3_net_1\, \I2.ROFFSET_n6_tz_i\, 
        \I2.N_4672\, \I1.LOAD_RESi_50_net_1\, 
        \I2.PIPE10_DT_17l29r\, \I5.N_73\, REGl7r, \I2.N_93_i_0\, 
        \I2.N_126_i_0\, \I2.DTE_2_1l15r_net_1\, 
        \I1.ISCK_0_sqmuxa_adt_net_134155_\, 
        \I1.N_1375_adt_net_134070_\, \I1.N_1192_adt_net_133761_\, 
        \I1.N_89_adt_net_128729_\, \I1.N_89_adt_net_128731_\, 
        \I1.N_89_adt_net_128728_\, \I1.N_89_adt_net_128717_\, 
        \I1.N_89_adt_net_128732_\, \I1.N_596_adt_net_124704_\, 
        \I1.REG_74_3_4_il380r_adt_net_123085_\, 
        \I1.REG_74l277r_adt_net_122979_\, 
        \I1.REG_74l278r_adt_net_122893_\, 
        \I1.REG_74l279r_adt_net_122807_\, 
        \I1.REG_74l280r_adt_net_122721_\, 
        \I1.REG_74l281r_adt_net_122635_\, 
        \I1.REG_74l282r_adt_net_122549_\, 
        \I1.REG_74l283r_adt_net_122463_\, 
        \I1.REG_74l284r_adt_net_122377_\, 
        \I1.REG_74l285r_adt_net_122291_\, 
        \I1.REG_74l286r_adt_net_122205_\, 
        \I1.REG_74l287r_adt_net_122119_\, 
        \I1.REG_74l288r_adt_net_122033_\, 
        \I1.REG_74l289r_adt_net_121947_\, 
        \I1.REG_74l290r_adt_net_121861_\, 
        \I1.REG_74l291r_adt_net_121775_\, 
        \I1.REG_74l292r_adt_net_121689_\, 
        \I1.REG_74_12_300_m8_i_0_adt_net_120083_\, 
        \I1.REG_74_12_348_m9_i_adt_net_115429_\, 
        \I1.REG_74_12_348_m9_i_adt_net_115430_\, 
        \I1.REG_74_12_348_m9_i_adt_net_115329_\, 
        \I1.REG_74_2_4_il228r_adt_net_115255_\, 
        \I1.N_273_10_adt_net_114361_\, 
        \I1.N_273_10_adt_net_114360_\, 
        \I1.REG_74_i_o2_0_0_364_m9_i_1_adt_net_114039_\, 
        \I1.N_1370_adt_net_112317_\, 
        \I1.N_50_0_adt_net_109760__net_1\, 
        \I1.N_79_adt_net_109340_\, 
        \I1.sstate_nsl2r_adt_net_107620_\, 
        \I1.N_420_i_adt_net_107486_\, 
        \I2.N_3834_i_0_adt_net_101432_\, 
        \I2.N346_adt_net_4075__net_1\, 
        \I1.N_41_9_adt_net_3739__net_1\, 
        \I1.N_1366_adt_net_112007_\, \I2.N_3_adt_net_940__net_1\, 
        \I3.N_637\, \I3.un13_reg_ads_0_a2_0_a3_net_1\, 
        \I3.N_283_adt_net_143533_\, 
        \I3.un17_reg_ads_0_a2_3_a3_net_1\, 
        \I3.un21_reg_ads_0_a2_0_a3_net_1\, 
        \I3.N_638_adt_net_134637_\, 
        \I3.un25_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un29_reg_ads_0_a2_0_a3_net_1\, 
        \I3.N_638_adt_net_134643_\, 
        \I3.un33_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un37_reg_ads_0_a2_1_a3_net_1\, 
        \I3.un44_reg_ads_0_a2_0_a3_net_1\, 
        \I3.N_638_adt_net_134639_\, 
        \I3.un47_reg_ads_0_a2_0_a3_net_1\, 
        \I3.VDBi_31l1r_adt_net_506111_\, 
        \I3.un51_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un54_reg_ads_0_a2_1_a3_net_1\, 
        \I3.un64_reg_ads_0_a2_3_a3_net_1\, \I3.N_549\, \I3.N_583\, 
        \I3.un71_reg_ads_0_a2_0_a3_net_1\, \I3.N_585\, 
        \I3.un76_reg_ads_0_a2_0_a3_net_1\, \I3.N_582\, 
        \I3.un81_reg_ads_0_a2_0_a3_net_1\, \I3.N_580\, 
        \I3.un86_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un1_REGMAP_30_adt_net_134453_\, 
        \I3.un91_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un96_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un101_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un106_reg_ads_0_a2_0_a3_net_1\, \I3.N_586\, 
        \I3.un111_reg_ads_0_a2_0_a3_net_1\, \I3.N_584\, 
        \I3.un116_reg_ads_0_a2_2_a3_net_1\, \I3.N_639\, 
        \I3.un121_reg_ads_0_a2_0_a3_net_1\, 
        \I3.N_68_adt_net_134367_\, \I3.N_641\, 
        \I3.un126_reg_ads_0_a2_1_a3_net_1\, 
        \I3.un131_reg_ads_0_a2_1_a3_net_1\, 
        \I3.un136_reg_ads_0_a2_2_a3_net_1\, 
        \I3.un141_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un1_REGMAP_30_0_a2_0_adt_net_134424_\, 
        \I3.un146_reg_ads_0_a2_1_a3_net_1\, 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135383_\, 
        \I3.un151_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un156_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un161_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un166_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un171_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un176_reg_ads_0_a2_0_a3_net_1\, 
        \I3.N_560_adt_net_134484_\, 
        \I3.un181_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un186_reg_ads_0_a2_1_a3_net_1\, 
        \I3.un191_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un196_reg_ads_0_a2_2_a3_net_1\, 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1570__net_1\, 
        \I3.un201_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un206_reg_ads_0_a2_1_a3_net_1\, 
        \I3.un211_reg_ads_0_a2_0_a3_net_1\, 
        \I3.un216_reg_ads_0_a2_1_a3_net_1\, 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135385_\, 
        \I3.un231_reg_ads_0_a2_4_a3_net_1\, 
        \I3.un235_reg_ads_0_a2_2_a3_net_1\, \I3.N_68\, 
        \I3.un1_REGMAP_30_0_a2_0_net_1\, \I3.N_58_i_0\, 
        \I3.un1_REGMAP_30_adt_net_134454_\, \I3.un1_REGMAP_30\, 
        \I3.N_560\, \I3.N_2083\, 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135544_\, \I3.N_2086\, 
        \I3.N_177\, \I3.N_178_adt_net_134608__net_1\, 
        \I3.N_178_adt_net_1360__net_1\, \I3.un1_REGMAP_34\, 
        \I3.N_590\, \I3.N_2053\, \I3.N_2042\, 
        \I3.N_638_adt_net_134642_\, \I3.N_2018\, \I3.N_2031\, 
        \I3.N_1641\, \I3.N_638_adt_net_134644_\, 
        \I3.VDBi_52l1r_net_1\, \I3.VDBi_55l1r_net_1\, \I3.N_1907\, 
        \I3.VDBi_20l12r_adt_net_140770_\, 
        \I3.VDBi_20l4r_adt_net_414785_\, 
        \I3.VDBi_29l4r_adt_net_621825_\, 
        \I3.N_638_adt_net_134645_\, \I3.N_638_adt_net_134647_\, 
        \I3.N_2056\, \I3.VDBi_57l7r_adt_net_142960__net_1\, 
        \I3.N_2040\, \I3.N_2033\, \I3.VDBi_52l3r_net_1\, 
        \I3.VDBi_55l3r_net_1\, \I3.VDBi_52l4r_net_1\, 
        \I3.VDBi_55l4r_net_1\, \I3.N_92\, \I3.VDBi_55l10r_net_1\, 
        \I3.VDBi_55l11r_net_1\, \I3.VDBi_55l12r_net_1\, 
        \I3.STATE1_tr24_i_0_a3_28_tz_i\, 
        \I3.STATE1_nsl2r_adt_net_134736__net_1\, 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1577__net_1\, 
        \I3.N_354_0\, \I3.N_2037\, \I3.N_2015\, \I3.N_2016\, 
        \I3.N_2017\, \I3.N_638\, \I3.N_437\, \I3.N_2036\, 
        \I3.N_2044\, \I3.N_2045\, \I3.N_2046\, \I1.N_1384\, 
        \I1.N_1377_adt_net_106750__net_1\, 
        \I1.N_1377_adt_net_1517__net_1\, \I1.N_337\, 
        \I1.N_1193_adt_net_134015_\, \I1.N_1194_adt_net_106064_\, 
        \I1.N_206_adt_net_105994_\, \I1.N_204_adt_net_105924_\, 
        \I1.N_202_adt_net_105770_\, \I1.N_1193\, \I1.N_653\, 
        \I1.N_1375\, \I1.ISI_54_net_1\, \I1.N_1207\, 
        \I1.SBYTE_0_sqmuxa_adt_net_105487_\, \I1.N_371_i\, 
        \I1.SBYTE_0_sqmuxa\, \I1.N_188\, \I1.SBYTE_59_net_1\, 
        \I1.N_190\, \I1.SBYTE_60_net_1\, \I1.N_202\, 
        \I1.SBYTE_61_net_1\, \I1.N_192\, \I1.SBYTE_62_net_1\, 
        \I1.N_204\, \I1.SBYTE_63_net_1\, \I1.N_206\, 
        \I1.SBYTE_64_net_1\, \I1.N_1194\, \I1.SBYTE_65_0\, 
        \I1.N_1366\, \I1.REG_74_4_i_a2_404_N_4_i\, \I1.N_374\, 
        \I1.N_41_8\, \I1.N_273_9\, \I1.N_273_6_i_0\, \I1.N_1370\, 
        \I1.N_41_9\, \I1.REG_74_8_0_o4_372_N_9_i\, 
        \I1.N_113_adt_net_126301__net_1\, 
        \I1.REG_74_8_308_m6_e_net_1\, \I1.REG_74_8_308_N_6_i\, 
        \I1.N_113_adt_net_126306__net_1\, \I1.N_242\, 
        \I1.REG_2_sqmuxa\, \I1.REG_1_sqmuxa\, \I1.REG_29_sqmuxa\, 
        \I1.REG_74l389r_adt_net_111128_\, \I1.REG_30_sqmuxa\, 
        \I1.N_185_9_adt_net_112166_\, 
        \I1.REG_74l397r_adt_net_110358_\, 
        \I1.REG_74l398r_adt_net_110272_\, 
        \I1.REG_74l399r_adt_net_110186_\, \I1.N_97_6\, 
        \I1.REG_74_8_0_N_6_i_i_0\, 
        \I1.N_193_adt_net_118653__net_1\, 
        \I1.N_193_adt_net_118660__net_1\, \I1.N_97_2\, 
        \I1.N_273_10\, \I1.N_57_9_i\, 
        \I1.REG_74_i_o2_i_0l364r_net_1\, \I1.REG_4_sqmuxa\, 
        \I1.REG_3_sqmuxa\, \I1.REG_5_sqmuxa\, \I1.N_179\, 
        \I1.N_396\, \I1.REG_74_12_300_N_15\, 
        \I1.REG_74_12_300_N_11_adt_net_120111_\, 
        \I1.REG_74_13_388_N_11_adt_net_109571_\, 
        \I1.N_395_adt_net_113231_\, \I1.REG_74_2_2_il340r\, 
        \I1.N_73_10_adt_net_117095_\, \I1.N_73_10\, 
        \I1.REG_74_3_4_il380r\, \I1.N_145_12_adt_net_123140_\, 
        \I1.N_145_12\, \I1.REG_6_sqmuxa\, 
        \I1.N_280_adt_net_130103_\, \I1.N_282_adt_net_130017_\, 
        \I1.N_1349_adt_net_129673_\, \I1.N_12233_i\, 
        \I1.REG_74l222r_adt_net_128480_\, 
        \I1.REG_74l224r_adt_net_128308_\, 
        \I1.REG_74l226r_adt_net_128136_\, 
        \I1.REG_74l227r_adt_net_128050_\, 
        \I1.N_89_adt_net_128733_\, \I1.REG_74_12_220_N_13\, 
        \I1.REG_74_12_220_m9_i_adt_net_127882_\, 
        \I1.REG_74_12_220_m9_i_net_1\, \I1.N_89_adt_net_128736_\, 
        \I1.REG_7_sqmuxa\, \I1.REG_74_2_4_il228r\, 
        \I1.REG_74_12_348_m9_i_adt_net_115422_\, \I1.N_240\, 
        \I1.REG_10_sqmuxa\, \I1.REG_9_sqmuxa\, 
        \I1.REG_74_1_404_m7_i_a5_0_net_1\, 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0_adt_net_125522_\, 
        \I1.N_592\, \I1.REG_74_0_iv_0_o2_0_il253r\, \I1.N_4867_i\, 
        \I1.N_395_adt_net_113232_\, \I1.N_395\, 
        \I1.N_658_adt_net_124758_\, 
        \I1.REG_74_i_o2_1_0tt_364_m2_e_net_1\, 
        \I1.REG_74_i_o2_1_0_364_N_5\, 
        \I1.REG_74_i_o2_1_0_364_N_2\, 
        \I1.REG_74_i_o2_1_0_364_N_6\, \I1.N_661_adt_net_114476_\, 
        \I1.REG_14_sqmuxa\, \I1.REG_13_sqmuxa\, 
        \I1.REG_74_12_284_m10_i_o6_net_1\, 
        \I1.REG_74_12_284_m10_i_0_i_adt_net_121593_\, 
        \I1.REG_74_12_284_m10_i_0_i\, 
        \I1.N_161_adt_net_121649__net_1\, \I1.REG_74_12_300_N_11\, 
        \I1.REG_74_1l308r_adt_net_120140_\, \I1.REG_18_sqmuxa\, 
        \I1.REG_17_sqmuxa\, \I1.REG_20_sqmuxa\, 
        \I1.REG_19_sqmuxa\, \I1.REG_22_sqmuxa\, 
        \I1.REG_21_sqmuxa\, \I1.REG_24_sqmuxa\, 
        \I1.REG_74_12_348_m9_i_net_1\, \I1.N_273_11_i\, 
        \I1.REG_23_sqmuxa\, \I1.REG_74_i_o2_0_0_364_m9_i_1_net_1\, 
        \I1.REG_74_1_396_m7_i_a5_0\, 
        \I1.REG_74_i_o2_0_0_364_N_14\, 
        \I1.REG_74_i_o2_0_0_m9_i_0_0_net_1\, 
        \I1.N_661_adt_net_114478_\, \I1.N_584\, 
        \I1.N_257_adt_net_111267_\, \I1.REG_74_1_380_m8_i_0_0\, 
        \I1.REG_74_1_380_N_14\, \I1.REG_74_1_380_N_15_i_i_i\, 
        \I1.N_249_adt_net_112440_\, \I1.REG_27_sqmuxa\, 
        \I1.REG_74_24_404_m3_e_net_1\, \I1.REG_74_2_3_il228r\, 
        \I1.REG_74_24_404_N_6_i_i\, \I1.N_257_adt_net_111276_\, 
        \I1.REG_28_sqmuxa\, \I1.N_265_adt_net_110486_\, 
        \I1.N_273_adt_net_109616_\, \I1.N_363\, \I1.N_413_i_0\, 
        \I1.N_485\, \I1.N_604\, \I1.N_1376_i_0\, \I1.N_415\, 
        \I1.N_68\, \I1.BITCNT_315_net_1\, \I1.N_416\, 
        \I1.BITCNT_316_net_1\, \I1.N_1199\, \I1.BITCNT_317_net_1\, 
        \I1.N_325\, \I1.N_328_i_0\, \I1.N_359\, \I1.N_56\, 
        \I1.N_404_i_i_0_i\, \I1.N_345\, \I1.N_369\, 
        \I1.N_409_i_i_0_i\, \I1.N_403_i_i_0_i\, 
        \I1.N_398_i_i_0_i\, \I1.sstate_nsl6r\, \I1.sstate_nsl9r\, 
        \I1.N_420_i\, \I1.sstate_ns_0_iv_0_il3r_net_1\, 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r\, 
        \I1.N_289_adt_net_107403_\, \I1.sstate_ns_il10r\, 
        \I2.CRC32_804_net_1\, \I2.N_57_i_0\, \I2.N_44_i_0\, 
        \I2.CRC32_798_net_1\, \I2.CRC32_7l3r_net_1\, 
        \I2.CRC32_796_net_1\, \I2.WOFFSET_827_net_1\, 
        \I2.EVNT_WORD_725_net_1\, \I2.EVNT_WORD_724_net_1\, 
        \I2.EVNT_WORD_723_net_1\, \I2.EVNT_WORD_722_net_1\, 
        \I2.EVNT_WORD_721_net_1\, \I2.EVNT_WORD_720_net_1\, 
        \I2.EVNT_WORD_719_net_1\, \I2.EVNT_WORD_718_net_1\, 
        \I2.EVNT_WORD_717_net_1\, \I2.EVNT_WORD_716_net_1\, 
        \I2.EVNT_WORD_715_net_1\, \I2.EVNT_WORD_714_net_1\, 
        \I2.EVNT_WORD_713_net_1\, \I2.SUB8_522_net_1\, 
        \I2.N434_adt_net_69831_\, \I2.SUB8_520_net_1\, 
        \I2.SUB8_519_net_1\, \I2.SUB8_518_net_1\, 
        \I2.N292_adt_net_68955_\, \I2.N291_adt_net_4302__net_1\, 
        \I2.SUB8_516_net_1\, 
        \I2.ADD_18x18_fast_I110_Y_0_adt_net_3684__net_1\, 
        \I2.N296_adt_net_69573_\, \I2.ADD_18x18_fast_I150_Y_0\, 
        \I2.SUB8_515_net_1\, \I2.N299\, \I2.STATE2l1r\, 
        \I2.DTE_21_1l4r_adt_net_39195_\, 
        \I2.DTE_21_1l5r_adt_net_39083_\, 
        \I2.DTE_21_1l6r_adt_net_38967_\, 
        \I2.DTE_21_1l7r_adt_net_38855_\, 
        \I2.DTE_21_1l8r_adt_net_38737_\, 
        \I2.DTE_21_1l9r_adt_net_38621_\, 
        \I2.DTE_21_1l10r_adt_net_38511_\, 
        \I2.DTE_21_1l11r_adt_net_38399_\, 
        \I2.DTE_21_1l12r_adt_net_38281_\, 
        \I2.DTE_21_1l13r_adt_net_38165_\, 
        \I2.DTE_21_1l14r_adt_net_38053_\, 
        \I2.DTE_21_1l15r_adt_net_37935_\, 
        \I2.DTE_21_1l16r_adt_net_37819_\, 
        \I2.DTE_21_1l19r_adt_net_37709_\, 
        \I2.INC_EVNT_NUM_759_net_1\, \I2.REG_1_n1_0_net_1\, 
        \I2.REG_1_n1_net_1\, \I2.N_3844\, \I2.REG_1_n2_0_net_1\, 
        \I2.REG_1_n2_net_1\, \I2.N_3824_adt_net_90291_\, 
        \I2.N_3845\, \I2.N_3831\, \I2.REG_1_n3_net_1\, 
        \I2.N_3832\, \I2.REG_1_n4_net_1\, \I2.N_3847\, 
        \I2.N_3833_i_0\, \I2.REG_1_n5_net_1\, \I2.REG_1_n6_net_1\, 
        \I2.N_3849\, \I2.N_3835_i_0\, \I2.REG_1_n7_net_1\, 
        \I2.N_3836_i_0\, \I2.REG_1_n8_net_1\, \I2.N_129\, 
        \I2.N_3838_adt_net_101306_\, \I2.N_3852\, \I2.N_3837_i_0\, 
        \I2.REG_1_n9_net_1\, \I2.N_3853\, \I2.N_3838\, 
        \I2.REG_1_n10_net_1\, \I2.N_3839_i_0_adt_net_101262_\, 
        \I2.N_3824_adt_net_90285_\, \I2.N_131\, 
        \I2.N_3840_adt_net_101218_\, \I2.N_3839_i_0\, 
        \I2.REG_1_n11_net_1\, \I2.N_3856\, \I2.N_3840\, 
        \I2.REG_1_n12_net_1\, \I2.N_3841_i_0_adt_net_101174_\, 
        \I2.N_136_1\, \I2.N_3841_i_0\, \I2.REG_1_n13_net_1\, 
        \I2.N_3824_adt_net_90287_\, \I2.N_3824_adt_net_90294_\, 
        \I2.N_138\, \I2.N_3859\, \I2.N_3842_i_0\, 
        \I2.REG_1_n14_net_1\, \I2.N_3824_adt_net_90293_\, 
        \I2.N_3843\, \I2.REG_1_n15_net_1\, 
        \I2.N_3824_adt_net_90289_\, \I2.N_3824_adt_net_90295_\, 
        \I2.SUB9_1l5r\, \I2.SUB9_1l6r\, \I2.N344\, \I2.SUB9_1l7r\, 
        \I2.N469\, \I2.SUB9_1l8r\, \I2.N466_adt_net_71184_\, 
        \I2.N340\, \I2.N466\, \I2.SUB9_1l9r\, \I2.N304\, 
        \I2.N463_adt_net_70886_\, \I2.N338\, \I2.N463\, 
        \I2.SUB9_1l10r\, \I2.N302\, \I2.N460_adt_net_70355_\, 
        \I2.N336\, \I2.N460\, \I2.ADD_18x18_fast_I148_Y_0\, 
        \I2.SUB9_1l11r\, \I2.N457_adt_net_69532_\, \I2.N334\, 
        \I2.N457\, \I2.ADD_18x18_fast_I149_Y_0\, \I2.SUB9_1l12r\, 
        \I2.N298\, \I2.N333\, \I2.I114_un1_Y\, \I2.I94_un1_Y\, 
        \I2.N297\, \I2.N332\, \I2.N454_i\, \I2.SUB9_1l13r\, 
        \I2.N296\, \I2.N331\, \I2.I113_un1_Y\, \I2.I92_un1_Y\, 
        \I2.N295\, \I2.N330\, \I2.N451_i\, 
        \I2.ADD_18x18_fast_I151_Y_0\, \I2.SUB9_1l14r\, \I2.N294\, 
        \I2.N328_adt_net_70573_\, \I2.N329\, 
        \I2.I112_un1_Y_adt_net_71518_\, \I2.N328\, 
        \I2.N436_adt_net_70670_\, \I2.N448_i_adt_net_71546_\, 
        \I2.N448_i\, \I2.ADD_18x18_fast_I152_Y_0\, 
        \I2.SUB9_1l15r\, \I2.N292\, \I2.N327\, 
        \I2.I111_un1_Y_adt_net_71419_\, \I2.N291\, \I2.N326\, 
        \I2.N434_adt_net_3677__net_1\, \I2.N445_i_adt_net_71447_\, 
        \I2.N445_i\, \I2.SUB9_1l16r\, \I2.N290\, 
        \I2.I110_un1_Y_adt_net_71212_\, \I2.I110_un1_Y\, 
        \I2.ADD_18x18_fast_I110_Y_0\, \I2.N442_i_adt_net_71348_\, 
        \I2.N442_i\, \I2.SUB9_1l17r\, \I2.N268\, 
        \I2.N436_adt_net_1185__net_1\, \I2.N436_adt_net_70753_\, 
        \I2.N288\, \I2.I109_un1_Y_adt_net_70914_\, 
        \I2.I109_un1_Y\, \I2.N287\, \I2.N434_adt_net_69748_\, 
        \I2.ADD_18x18_fast_I109_Y_0\, \I2.N439_i_adt_net_71055_\, 
        \I2.N439_i\, \I2.ADD_18x18_fast_I155_Y_0\, 
        \I2.SUB9_1l18r\, \I2.N271\, \I2.N321\, \I2.N436\, 
        \I2.ADD_18x18_fast_I156_Y_0\, \I2.SUB9_1l19r\, \I2.N284\, 
        \I2.N434\, \I2.SUB9_1l20r\, \I2.WROi_10_1\, 
        \I2.CRC32_7_il1r\, \I2.N_4293\, \I2.WOFFSETl1r\, 
        \I2.ADE_4l0r_net_1\, \I2.ADO_3l0r_net_1\, \I2.WOFFSETl2r\, 
        \I2.ADE_4l1r_net_1\, \I2.ADO_3l1r_net_1\, \I2.WOFFSETl3r\, 
        \I2.ADE_4l2r_net_1\, \I2.ADO_3l2r_net_1\, \I2.WOFFSETl4r\, 
        \I2.ADE_4l3r_net_1\, \I2.ADO_3l3r_net_1\, \I2.WOFFSETl5r\, 
        \I2.ADE_4l4r_net_1\, \I2.ADO_3l4r_net_1\, \I2.WOFFSETl6r\, 
        \I2.ADE_4l5r_net_1\, \I2.ADO_3l5r_net_1\, \I2.WOFFSETl7r\, 
        \I2.ADE_4l6r_net_1\, \I2.ADO_3l6r_net_1\, \I2.WOFFSETl8r\, 
        \I2.ADE_4l7r_net_1\, \I2.ADO_3l7r_net_1\, \I2.WOFFSETl9r\, 
        \I2.ADE_4l8r_net_1\, \I2.ADO_3l8r_net_1\, 
        \I2.WOFFSETl10r\, \I2.ADE_4l9r_net_1\, 
        \I2.ADO_3l9r_net_1\, \I2.WOFFSETl11r\, 
        \I2.ADE_4l10r_net_1\, \I2.ADO_3l10r_net_1\, 
        \I2.ADO_3l11r_net_1\, \I2.ADE_4l11r_net_1\, 
        \I2.DTE_21_1l11r_Rd1__net_1\, \I2.DTE_1l11r\, 
        \I2.DTE_21_1l14r_Rd1__net_1\, \I2.DTE_1l14r\, 
        \I2.DTE_21_1l15r_Rd1__net_1\, \I2.DTE_1l15r\, 
        \I2.DTE_21_1l20r_Rd1__net_1\, \I2.DTE_1l20r\, 
        \I2.DTE_1l22r\, \I2.DTE_1l23r\, \I2.DTE_1l24r\, 
        \I2.DTO_1l5r_net_1\, \I2.DTO_16_1l11r_Rd1__net_1\, 
        \I2.DTO_1l11r\, \I2.DTO_16_1l14r_Rd1__net_1\, 
        \I2.DTO_1l14r\, \I2.DTO_16_1l15r_Rd1__net_1\, 
        \I2.DTO_1l15r\, \I2.DTO_16_1l20r_Rd1__net_1\, 
        \I2.DTO_1l20r\, \I2.ROFFSET_c7_net_1\, 
        \I2.ROFFSET_c8_net_1\, \I2.ROFFSET_c9_net_1\, 
        \I2.ROFFSET_c10_net_1\, \I2.ROFFSET_n11_tz_i\, 
        \I2.ROFFSET_n10_tz_i\, \I2.ROFFSET_n9_tz_i\, 
        \I2.ROFFSET_n8_tz_i\, \I2.ROFFSET_n7_tz_i\, \I2.N_201\, 
        \I2.N_207\, \I2.G_EVNT_NUM_n9_adt_net_26657_\, \I2.N_218\, 
        \I2.N_287_adt_net_26828_\, \I2.N_282\, \I2.N_281\, 
        \I2.EVNT_NUM_c9_net_1\, \I2.EVNT_NUM_n10_tz_i\, 
        \I2.WPAGEe\, \I2.WPAGE_948_net_1\, \I2.WPAGE_949_net_1\, 
        \I2.WPAGE_950_net_1\, \I2.WPAGE_951_net_1\, 
        \I2.WPAGE_c1_net_1\, \I2.WPAGE_c2_net_1\, 
        \I2.WPAGE_n3_net_1\, \I2.WPAGE_n2_net_1\, 
        \I2.WPAGE_n1_net_1\, \I2.N_28_i_0\, \I5.DATA_12l8r_net_1\, 
        \I5.DATA_12l9r_net_1\, \I5.DATA_12l10r_net_1\, 
        \I5.DATA_12l11r_net_1\, \I5.DATA_12l12r_net_1\, 
        \I5.DATA_12l13r_net_1\, \I5.DATA_12l14r_net_1\, 
        \I5.DATA_12l15r_net_1\, \I5.CHAIN_SELECT_4_net_1\, 
        \I5.COMMAND_4l0r_net_1\, \I5.COMMAND_4l1r_net_1\, 
        \I5.COMMAND_4l2r_net_1\, \I5.COMMAND_4l8r_net_1\, 
        \I5.COMMAND_4l9r_net_1\, \I5.COMMAND_4l10r_net_1\, 
        \I5.COMMAND_4l11r_net_1\, \I5.COMMAND_4l12r_net_1\, 
        \I5.COMMAND_4l13r_net_1\, \I5.COMMAND_4l14r_net_1\, 
        \I5.COMMAND_4l15r_net_1\, \I5.PULSE_I2C_net_1\, 
        \I5.N_464\, \I2.WPAGEl15r_net_1\, \I2.WPAGEl14r_net_1\, 
        \I2.WPAGEl13r_net_1\, \I2.WPAGEl12r_net_1\, 
        \I1.sstatel1r_net_1\, \I1.BITCNTl0r_net_1\, 
        \I1.BITCNTl1r_net_1\, \I1.BITCNTl2r_net_1\, 
        \I1.sstatel7r_net_1\, \I3.RAMDTSl4r_net_1\, 
        \I3.RAMDTSl3r_net_1\, \I3.RAMDTSl1r_net_1\, 
        \I1.sstatel0r_net_1\, \I3.RAMDTSl9r_net_1\, 
        \I3.RAMDTSl10r_net_1\, \I3.RAMDTSl11r_net_1\, 
        \I3.RAMDTSl12r_net_1\, 
        \I2.N_2864_0_adt_net_835284_Rd1__net_1\, 
        \I2.N_4293_Rd1__net_1\, \I2.DTE_1l24r_Rd1__net_1\, 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\, 
        \I2.DTE_1l23r_Rd1__net_1\, \I2.DTE_1l22r_Rd1__net_1\, 
        \PULSEl0r\, \I2.WOFFSETl1r_Rd1__net_1\, 
        \I2.N_4244_Rd1__net_1\, 
        \I2.N_2828_adt_net_1062__adt_net_835312_Rd1__net_1\, 
        \I2.WOFFSETl2r_Rd1__net_1\, \I2.N_4245_Rd1__net_1\, 
        \I2.WOFFSETl3r_Rd1__net_1\, \I2.N_4246_Rd1__net_1\, 
        \I2.WOFFSETl4r_Rd1__net_1\, \I2.N_4247_Rd1__net_1\, 
        \I2.WOFFSETl5r_Rd1__net_1\, \I2.N_4248_Rd1__net_1\, 
        \I2.N_2828_adt_net_1062__adt_net_835308_Rd1__net_1\, 
        \I2.WOFFSETl6r_Rd1__net_1\, \I2.N_4249_Rd1__net_1\, 
        \I2.WOFFSETl7r_Rd1__net_1\, \I2.N_4250_Rd1__net_1\, 
        \I2.WOFFSETl8r_Rd1__net_1\, \I2.N_4251_Rd1__net_1\, 
        \I2.WOFFSETl9r_Rd1__net_1\, \I2.N_4252_Rd1__net_1\, 
        \I2.N_2828_adt_net_1062__adt_net_835304_Rd1__net_1\, 
        \I2.WOFFSETl10r_Rd1__net_1\, \I2.N_4253_Rd1__net_1\, 
        \I2.WOFFSETl11r_Rd1__net_1\, \I2.N_4254_Rd1__net_1\, 
        \I2.DTE_1l11r_Rd1__net_1\, 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, 
        \I2.DTE_1l14r_Rd1__net_1\, 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\, 
        \I2.DTE_1l15r_Rd1__net_1\, \I2.DTE_1l20r_Rd1__net_1\, 
        \I2.DTO_1l11r_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834772_Rd1__net_1\, 
        \I2.DTO_1l14r_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834768_Rd1__net_1\, 
        \I2.DTO_1l15r_Rd1__net_1\, \I2.DTO_1l20r_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834760_Rd1__net_1\, 
        \I1.REG_74_2_2_il340r_adt_net_117067_\, \I2.DTO_16_1l20r\, 
        \I2.DTO_16_1l15r\, \I2.DTO_16_1l14r\, \I2.DTO_16_1l11r\, 
        \I2.DTE_21_1l20r\, \I2.DTE_21_1l15r\, \I2.DTE_21_1l14r\, 
        \I2.DTE_21_1l11r\, \I1.N_50_0_adt_net_109757__net_1\, 
        \I2.N_3836_i_0_adt_net_101388_\, \I2.N288_adt_net_68878_\, 
        \I2.DTE_21_1l22r_Rd1_\, \I2.DTE_21_1l23r_Rd1_\, 
        \I2.DTE_21_1l24r_Rd1_\, \I1.N_1375_adt_net_134063_\, 
        \I1.N_1367_i\, \I1.N_145_12_adt_net_123179_\, \I1.N_347\, 
        \I1.REG_74_11_a0l404r_net_1\, \I2.N_3834_i_0\, 
        \I2.N301_1\, \I2.N300\, \I2.ADD_18x18_fast_I154_Y_0\, 
        \I2.N_4330\, \I2.N_280\, \I2.N_198\, \I2.DTO_1l31r_net_1\, 
        \I2.DTO_1l30r_net_1\, \I2.DTO_1l29r_net_1\, 
        \I2.DTO_1l28r_net_1\, \I2.DTO_1l27r\, \I2.DTO_1l26r\, 
        \I2.DTO_1l25r\, \I2.DTO_1l24r\, \I2.DTO_1l23r\, 
        \I2.DTO_1l22r\, \I2.DTO_1l21r\, \I2.DTO_1l19r\, 
        \I2.DTO_1l18r\, \I2.DTO_1l17r\, \I2.DTO_1l16r\, 
        \I2.DTO_1l13r\, \I2.DTO_1l12r\, \I2.DTO_1l10r\, 
        \I2.DTO_1l9r\, \I2.DTO_1l8r\, \I2.DTO_1l7r\, 
        \I2.DTO_1l6r\, \I2.DTO_1_879_net_1\, \I2.DTO_1l4r\, 
        \I2.DTO_1l3r_net_1\, \I2.DTO_1l2r_net_1\, 
        \I2.DTO_1l1r_net_1\, \I2.DTO_1l0r_net_1\, \I2.DTE_1l27r\, 
        \I2.DTE_1l26r\, \I2.DTE_1l25r\, \I2.DTE_1l21r\, 
        \I2.DTE_2_1l11r_net_1\, \I2.DTE_2_1l10r_net_1\, 
        \I2.DTE_2_1l9r_net_1\, \I2.DTE_2_1l8r_net_1\, 
        \I2.DTE_1l7r\, \I2.DTE_2_1l7r_net_1\, 
        \I2.DTE_2_1l6r_net_1\, \I2.DTE_2_1l5r_net_1\, 
        \I2.DTE_2_1l4r_net_1\, \I2.WOFFSETl12r\, 
        \I2.PIPE10_DT_17l30r\, 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_2_i_adt_net_271662_\, 
        \I1.N_457\, \I2.N306\, \I2.DTE_1l4r\, \I2.DTE_1l6r\, 
        \I2.DTE_1l8r\, \I2.DTE_1l9r\, \I2.DTE_1l10r\, 
        \I2.DTE_1l12r\, \I2.DTE_1l13r\, \I2.DTE_1l16r\, 
        \I2.DTE_1l19r\, \I2.DTE_1l17r\, \I2.DTE_1l18r\, 
        \I2.EVNT_NUM_n9_tz_i\, 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835168_Rd1__net_1\, 
        \I2.DTE_21_1l22r_adt_net_37395_Rd1__net_1\, 
        \I2.DTE_21_1l23r_adt_net_37285_Rd1__net_1\, 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835180_Rd1__net_1\, 
        \I2.DTE_21_1l24r_adt_net_37175_Rd1__net_1\, 
        \I2.DTO_1l27r_Rd1__net_1\, \I2.DTO_16_1l27r_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834756_Rd1__net_1\, 
        \I2.DTO_1l26r_Rd1__net_1\, \I2.DTO_16_1l26r_Rd1__net_1\, 
        \I2.DTO_1l25r_Rd1__net_1\, \I2.DTO_16_1l25r_Rd1__net_1\, 
        \I2.DTO_1l24r_Rd1__net_1\, \I2.DTO_16_1l24r_Rd1__net_1\, 
        \I2.DTO_1l23r_Rd1__net_1\, \I2.DTO_16_1l23r_Rd1__net_1\, 
        \I2.DTO_1l22r_Rd1__net_1\, \I2.DTO_16_1l22r_Rd1__net_1\, 
        \I2.DTO_1l21r_Rd1__net_1\, \I2.DTO_16_1l21r_Rd1__net_1\, 
        \I2.DTO_1l19r_Rd1__net_1\, \I2.DTO_16_1l19r_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834764_Rd1__net_1\, 
        \I2.DTO_1l18r_Rd1__net_1\, \I2.DTO_16_1l18r_Rd1__net_1\, 
        \I2.DTO_1l17r_Rd1__net_1\, \I2.DTO_16_1l17r_Rd1__net_1\, 
        \I2.DTO_1l16r_Rd1__net_1\, \I2.DTO_16_1l16r_Rd1__net_1\, 
        \I2.DTO_1l13r_Rd1__net_1\, \I2.DTO_16_1l13r_Rd1__net_1\, 
        \I2.DTO_1l12r_Rd1__net_1\, \I2.DTO_16_1l12r_Rd1__net_1\, 
        \I2.DTO_1l10r_Rd1__net_1\, \I2.DTO_16_1l10r_Rd1__net_1\, 
        \I2.DTO_1l9r_Rd1__net_1\, \I2.DTO_16_1l9r_Rd1__net_1\, 
        \I2.DTO_1l8r_Rd1__net_1\, \I2.DTO_16_1l8r_Rd1__net_1\, 
        \I2.DTO_1l7r_Rd1__net_1\, \I2.DTO_16_1l7r_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834776_Rd1__net_1\, 
        \I2.DTO_1l6r_Rd1__net_1\, \I2.DTO_16_1l6r_Rd1__net_1\, 
        \I2.DTO_1l4r_Rd1__net_1\, \I2.DTO_16_1l4r_Rd1__net_1\, 
        \I2.DTE_1l27r_Rd1__net_1\, \I2.DTE_21_1l27r_Rd1__net_1\, 
        \I2.DTE_1l26r_Rd1__net_1\, \I2.DTE_21_1l26r_Rd1__net_1\, 
        \I2.DTE_1l25r_Rd1__net_1\, \I2.N_4644_Rd1__net_1\, 
        \I2.DTE_1l21r_Rd1__net_1\, \I2.DTE_21_1l21r_Rd1__net_1\, 
        \I2.DTE_1l7r_Rd1__net_1\, \I2.DTE_21_1l7r_Rd1__net_1\, 
        \I2.WOFFSETl12r_Rd1__net_1\, \I2.N_4255_Rd1__net_1\, 
        \I2.DTE_1l4r_Rd1__net_1\, \I2.DTE_21_1l4r_Rd1__net_1\, 
        \I2.N_2868_1_adt_net_836004_Rd1__net_1\, 
        \I2.DTE_1l6r_Rd1__net_1\, \I2.DTE_21_1l6r_Rd1__net_1\, 
        \I2.DTE_1l8r_Rd1__net_1\, \I2.DTE_21_1l8r_Rd1__net_1\, 
        \I2.DTE_1l9r_Rd1__net_1\, \I2.DTE_21_1l9r_Rd1__net_1\, 
        \I2.DTE_1l10r_Rd1__net_1\, \I2.DTE_21_1l10r_Rd1__net_1\, 
        \I2.DTE_1l12r_Rd1__net_1\, \I2.DTE_21_1l12r_Rd1__net_1\, 
        \I2.DTE_1l13r_Rd1__net_1\, \I2.DTE_21_1l13r_Rd1__net_1\, 
        \I2.DTE_1l16r_Rd1__net_1\, \I2.DTE_21_1l16r_Rd1__net_1\, 
        \I2.DTE_1l19r_Rd1__net_1\, \I2.DTE_21_1l19r_Rd1__net_1\, 
        \I2.DTE_1l17r_Rd1__net_1\, \I2.DTE_21_1l17r_Rd1__net_1\, 
        \I2.N_2868_1_adt_net_835988_Rd1__net_1\, 
        \I2.DTE_1l18r_Rd1__net_1\, 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_Rd1__net_1\, 
        \I1.REG_74l381r_adt_net_111921_\, 
        \I1.REG_74l382r_adt_net_111835_\, 
        \I1.REG_74l383r_adt_net_111749_\, 
        \I1.REG_74l384r_adt_net_111663_\, 
        \I1.REG_74l385r_adt_net_111577_\, 
        \I1.REG_74l386r_adt_net_111491_\, 
        \I1.REG_74l387r_adt_net_111405_\, 
        \I1.REG_74l388r_adt_net_111319_\, \I1.NCS0_net_1\, 
        \I1.sstatel9r_net_1\, \I1.sstatel2r_net_1\, 
        \I1.sstatel10r_net_1\, \I1.LUT_net_1\, 
        \I1.sstatel8r_net_1\, \F_SCK_c\, \REGl205r\, \REGl206r\, 
        \REGl210r\, \REGl213r\, \REGl222r\, \REGl224r\, 
        \REGl226r\, \REGl227r\, \REGl228r\, \REGl245r\, 
        \REGl246r\, \REGl247r\, \REGl248r\, \REGl249r\, 
        \REGl250r\, \REGl251r\, \REGl252r\, \REGl253r\, 
        \REGl254r\, \REGl255r\, \REGl256r\, \REGl257r\, 
        \REGl258r\, \REGl259r\, \REGl260r\, \REGl365r\, 
        \REGl366r\, \REGl367r\, \REGl368r\, \REGl369r\, 
        \REGl370r\, \REGl371r\, \REGl372r\, \REGl373r\, 
        \REGl374r\, \REGl375r\, \REGl376r\, \REGl377r\, 
        \REGl378r\, \REGl379r\, \REGl380r\, \REGl389r\, 
        \REGl390r\, \REGl391r\, \REGl392r\, \REGl393r\, 
        \REGl394r\, \REGl395r\, \REGl396r\, \REGl397r\, 
        \REGl398r\, \REGl399r\, \REGl400r\, \REGl401r\, 
        \REGl402r\, \REGl403r\, \REGl404r\, \I1.BYTECNTl8r_net_1\, 
        \I1.BYTECNTl7r_net_1\, \I1.BYTECNTl6r_net_1\, 
        \I1.BYTECNTl5r_net_1\, \I1.BYTECNT_i_0_il4r_net_1\, 
        \I1.BYTECNTl3r_net_1\, \I1.BYTECNTl2r_net_1\, 
        \I1.BYTECNT_i_0_il1r_net_1\, \I1.BYTECNTl0r_net_1\, 
        \I1.PAGECNTl7r_net_1\, \REGl225r\, \REGl223r\, \REGl221r\, 
        \REGl220r\, \REGl219r\, \REGl218r\, \REGl217r\, 
        \REGl216r\, \REGl215r\, \REGl214r\, \REGl356r\, 
        \REGl355r\, \REGl354r\, \REGl353r\, \REGl352r\, 
        \REGl351r\, \REGl350r\, \REGl349r\, \REGl348r\, 
        \REGl347r\, \REGl346r\, \REGl345r\, \REGl344r\, 
        \REGl343r\, \REGl342r\, \REGl341r\, \REGl381r\, 
        \REGl382r\, \REGl383r\, \REGl384r\, \REGl385r\, 
        \REGl386r\, \REGl387r\, \REGl388r\, \I1.N_304_Rd1__net_1\, 
        \I1.PAGECNTl4r_adt_net_835120_Rd1__net_1\, 
        \I1.PAGECNTl3r_adt_net_835116_Rd1__net_1\, 
        \I1.PAGECNTl2r_adt_net_834908_Rd1__net_1\, 
        \I1.PAGECNTl1r_adt_net_834904_Rd1__net_1\, \REGl364r\, 
        \REGl363r\, \REGl362r\, \REGl361r\, \REGl360r\, 
        \REGl359r\, \REGl358r\, \REGl357r\, \REGl277r\, 
        \REGl278r\, \REGl279r\, \REGl280r\, \REGl281r\, 
        \REGl282r\, \REGl283r\, \REGl284r\, \REGl285r\, 
        \REGl286r\, \REGl287r\, \REGl288r\, \REGl289r\, 
        \REGl290r\, \REGl291r\, \REGl292r\, \REGl293r\, 
        \REGl294r\, \REGl295r\, \REGl296r\, \REGl297r\, 
        \REGl298r\, \REGl299r\, \REGl300r\, \REGl301r\, 
        \REGl302r\, \REGl303r\, \REGl304r\, \REGl305r\, 
        \REGl306r\, \REGl307r\, \REGl308r\, \REGl165r\, 
        \REGl166r\, \REGl167r\, \REGl168r\, \REGl169r\, 
        \REGl170r\, \REGl171r\, \REGl172r\, \REGl173r\, 
        \REGl174r\, \REGl175r\, \REGl176r\, \REGl177r\, 
        \REGl178r\, \REGl179r\, \REGl180r\, \REGl181r\, 
        \REGl182r\, \REGl183r\, \REGl184r\, \REGl185r\, 
        \REGl186r\, \REGl187r\, \REGl188r\, \REGl189r\, 
        \REGl190r\, \REGl191r\, \REGl192r\, \REGl193r\, 
        \REGl194r\, \REGl195r\, \REGl196r\, \REGl197r\, 
        \REGl198r\, \REGl199r\, \REGl200r\, \REGl201r\, 
        \REGl202r\, \REGl203r\, \REGl204r\, \REGl207r\, 
        \REGl208r\, \REGl209r\, \REGl211r\, \REGl212r\, 
        \REGl229r\, \REGl230r\, \REGl231r\, \REGl232r\, 
        \REGl233r\, \REGl234r\, \REGl235r\, \REGl236r\, 
        \REGl237r\, \REGl238r\, \REGl239r\, \REGl240r\, 
        \REGl241r\, \REGl242r\, \REGl243r\, \REGl244r\, 
        \REGl261r\, \REGl262r\, \REGl263r\, \REGl264r\, 
        \REGl265r\, \REGl266r\, \REGl267r\, \REGl268r\, 
        \REGl269r\, \REGl270r\, \REGl271r\, \REGl272r\, 
        \REGl273r\, \REGl274r\, \REGl275r\, \REGl276r\, 
        \REGl309r\, \REGl310r\, \REGl311r\, \REGl312r\, 
        \REGl313r\, \REGl314r\, \REGl315r\, \REGl316r\, 
        \REGl317r\, \REGl318r\, \REGl319r\, \REGl320r\, 
        \REGl321r\, \REGl322r\, \REGl323r\, \REGl324r\, 
        \REGl325r\, \REGl326r\, \REGl327r\, \REGl328r\, 
        \REGl329r\, \REGl330r\, \REGl331r\, \REGl332r\, 
        \REGl333r\, \REGl334r\, \REGl335r\, \REGl336r\, 
        \REGl337r\, \REGl338r\, \REGl339r\, \REGl340r\, 
        \I1.N_299_adt_net_833868_Rd1__net_1\, 
        \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, 
        \I1.N_311_i_i_Rd1__net_1\, \I2.DTO_1_874_net_1\, 
        \I2.DTO_1_875_net_1\, \I2.DTO_1_876_net_1\, 
        \I2.DTO_1_877_net_1\, \I2.DTO_1_902_net_1\, 
        \I2.DTO_1_903_net_1\, \I2.DTO_1_904_net_1\, 
        \I2.DTO_1_905_net_1\, \I2.N_4337\, 
        \I2.ADD_18x18_fast_I153_Y_0\, \I1.N_310_Rd1__net_1\, 
        \I1.N_181\, \I1.N_185_9\, \I1.N_223\, 
        \I1.un1_sbyte13_1_i_1\, \I1.N_161_adt_net_1449__net_1\, 
        \I1.REG_74_13_388_N_11\, \I1.N_656\, \I1.N_596\, 
        \I1.REG_25_sqmuxa\, \I1.N_593\, \I1.N_97\, 
        \I1.N_113_adt_net_3714__net_1\, \I1.N_201_9\, 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, 
        \I1.N_661_adt_net_114485_\, 
        \I1.REG_74l341r_adt_net_116928_\, 
        \I1.REG_74l342r_adt_net_116842_\, 
        \I1.REG_74l343r_adt_net_116756_\, 
        \I1.REG_74l344r_adt_net_116670_\, 
        \I1.REG_74l345r_adt_net_116584_\, 
        \I1.REG_74l346r_adt_net_116498_\, 
        \I1.REG_74l347r_adt_net_116412_\, 
        \I1.REG_74l348r_adt_net_116326_\, \I2.N313_0\, \I2.N308\, 
        \I1.LUT_55_adt_net_133935_\, 
        \I1.REG_74l213r_adt_net_129378_\, 
        \I1.REG_74l214r_adt_net_129292_\, 
        \I1.REG_74l216r_adt_net_129120_\, 
        \I1.REG_74l217r_adt_net_129034_\, 
        \I1.REG_74l218r_adt_net_128948_\, 
        \I1.REG_74l219r_adt_net_128862_\, 
        \I1.REG_74l228r_adt_net_127964_\, 
        \I1.REG_74l261r_adt_net_124629_\, 
        \I1.REG_74l263r_adt_net_124457_\, 
        \I1.REG_74l265r_adt_net_124285_\, 
        \I1.REG_74l266r_adt_net_124199_\, 
        \I1.REG_74l267r_adt_net_124113_\, 
        \I1.REG_74l268r_adt_net_124027_\, 
        \I1.REG_74l270r_adt_net_123818_\, 
        \I1.REG_74l272r_adt_net_123646_\, 
        \I1.REG_74l274r_adt_net_123474_\, 
        \I1.REG_74l275r_adt_net_123388_\, 
        \I1.REG_74l276r_adt_net_123302_\, 
        \I1.N_257_adt_net_111279_\, 
        \I1.REG_74l400r_adt_net_110100_\, 
        \I1.REG_74l401r_adt_net_110014_\, 
        \I1.REG_74l402r_adt_net_109928_\, 
        \I1.REG_74l403r_adt_net_109842_\, 
        \I1.REG_74l404r_adt_net_109656_\, \I1.N_324\, 
        \I1.NCS0_56_net_1\, \I1.N_65_12\, \I1.N_89\, \I1.N_658\, 
        \I1.REG_74_1l308r\, \I1.REG_74_0l348r\, \I1.N_660\, 
        \I1.N_1383\, \I1.PAGECNTe\, \I1.sstate_nsl1r\, \I1.N_289\, 
        \I1.N_43_i_0\, \I1.ISCK_0_sqmuxa\, \I1.N_182_i\, 
        \I1.N_265\, \I1.N_65_adt_net_1433__net_1\, \I1.N_183_i_0\, 
        \I1.N_193_adt_net_1425__net_1\, \I1.REG_74_1l268r\, 
        \I1.N_249\, \I1.N_473\, \I1.N_153\, \I1.N_161\, 
        \I1.N_273\, FCS_c, \I1.LUT_55_net_1\, 
        \I1.REG_74l229r_adt_net_127710_\, 
        \I1.REG_74l230r_adt_net_127624_\, 
        \I1.REG_74l231r_adt_net_127538_\, 
        \I1.REG_74l232r_adt_net_127452_\, 
        \I1.REG_74l233r_adt_net_127366_\, 
        \I1.REG_74l234r_adt_net_127280_\, 
        \I1.REG_74l235r_adt_net_127194_\, 
        \I1.REG_74l236r_adt_net_127108_\, 
        \I1.REG_74l237r_adt_net_126985_\, 
        \I1.REG_74l238r_adt_net_126899_\, 
        \I1.REG_74l239r_adt_net_126813_\, 
        \I1.REG_74l240r_adt_net_126727_\, 
        \I1.REG_74l241r_adt_net_126641_\, 
        \I1.REG_74l242r_adt_net_126555_\, 
        \I1.REG_74l243r_adt_net_126469_\, 
        \I1.REG_74l244r_adt_net_126383_\, 
        \I1.REG_74l349r_adt_net_116203_\, 
        \I1.REG_74l350r_adt_net_116117_\, 
        \I1.REG_74l351r_adt_net_116031_\, 
        \I1.REG_74l352r_adt_net_115945_\, 
        \I1.REG_74l353r_adt_net_115859_\, 
        \I1.REG_74l354r_adt_net_115773_\, 
        \I1.REG_74l355r_adt_net_115687_\, 
        \I1.REG_74l356r_adt_net_115601_\, 
        \I1.REG_74l390r_adt_net_111042_\, 
        \I1.REG_74l391r_adt_net_110956_\, 
        \I1.REG_74l392r_adt_net_110870_\, 
        \I1.REG_74l393r_adt_net_110784_\, 
        \I1.REG_74l395r_adt_net_110612_\, 
        \I1.REG_74l396r_adt_net_110526_\, \I1.N_217\, \I1.N_225\, 
        \I1.REG_74l317r_adt_net_119303_\, 
        \I1.REG_74l318r_adt_net_119217_\, 
        \I1.REG_74l319r_adt_net_119131_\, 
        \I1.REG_74l320r_adt_net_119045_\, 
        \I1.REG_74l321r_adt_net_118959_\, 
        \I1.REG_74l322r_adt_net_118873_\, 
        \I1.REG_74l323r_adt_net_118787_\, 
        \I1.REG_74l324r_adt_net_118701_\, 
        \I1.N_1193_adt_net_133987__net_1\, \I1.N_105\, \I1.N_169\, 
        \I1.N_177\, \I1.N_257\, \I1.REG_74l325r_adt_net_118518_\, 
        \I1.REG_74l326r_adt_net_118432_\, 
        \I1.REG_74l327r_adt_net_118346_\, 
        \I1.REG_74l328r_adt_net_118260_\, 
        \I1.REG_74l329r_adt_net_118174_\, 
        \I1.REG_74l330r_adt_net_118088_\, 
        \I1.REG_74l331r_adt_net_118002_\, 
        \I1.REG_74l332r_adt_net_117916_\, 
        \I1.REG_74l333r_adt_net_117830_\, 
        \I1.REG_74l334r_adt_net_117744_\, 
        \I1.REG_74l335r_adt_net_117658_\, 
        \I1.REG_74l336r_adt_net_117572_\, 
        \I1.REG_74l337r_adt_net_117486_\, 
        \I1.REG_74l338r_adt_net_117400_\, 
        \I1.REG_74l339r_adt_net_117314_\, 
        \I1.REG_74l340r_adt_net_117228_\, \I1.N_602_i\, 
        \I1.N_387_i_0\, \I1.ISCK_53_net_1\, \I1.sstate_nsl2r\, 
        \I1.REG_74l165r_adt_net_133665_\, 
        \I1.REG_74l166r_adt_net_133579_\, 
        \I1.REG_74l167r_adt_net_133493_\, 
        \I1.REG_74l168r_adt_net_133407_\, 
        \I1.REG_74l169r_adt_net_133321_\, 
        \I1.REG_74l170r_adt_net_133235_\, 
        \I1.REG_74l171r_adt_net_133149_\, 
        \I1.REG_74l172r_adt_net_133063_\, 
        \I1.REG_74l174r_adt_net_132854_\, 
        \I1.REG_74l175r_adt_net_132768_\, 
        \I1.REG_74l177r_adt_net_132596_\, 
        \I1.REG_74l178r_adt_net_132510_\, 
        \I1.REG_74l181r_adt_net_132215_\, 
        \I1.REG_74l182r_adt_net_132129_\, 
        \I1.REG_74l183r_adt_net_132043_\, 
        \I1.REG_74l184r_adt_net_131957_\, 
        \I1.REG_74l185r_adt_net_131871_\, 
        \I1.REG_74l186r_adt_net_131785_\, 
        \I1.REG_74l187r_adt_net_131699_\, 
        \I1.REG_74l188r_adt_net_131613_\, 
        \I1.REG_74l189r_adt_net_131527_\, 
        \I1.REG_74l190r_adt_net_131441_\, 
        \I1.REG_74l192r_adt_net_131269_\, 
        \I1.REG_74l193r_adt_net_131183_\, 
        \I1.REG_74l195r_adt_net_131011_\, 
        \I1.REG_74l196r_adt_net_130925_\, 
        \I1.N_129_adt_net_130791_\, \I1.N_1337_adt_net_130705_\, 
        \I1.N_1338_adt_net_130619_\, \I1.N_1339_adt_net_130533_\, 
        \I1.N_1340_adt_net_130447_\, \I1.N_1341_adt_net_130361_\, 
        \I1.N_1342_adt_net_130275_\, \I1.N_1343_adt_net_130189_\, 
        \I1.N_1346_adt_net_129931_\, \I1.N_1347_adt_net_129845_\, 
        \I1.N_1348_adt_net_129759_\, \I1.N_144_adt_net_129587_\, 
        \I1.N_1350_adt_net_129501_\, 
        \I1.REG_74l215r_adt_net_129206_\, 
        \I1.REG_74l220r_adt_net_128776_\, 
        \I1.REG_74l221r_adt_net_128566_\, 
        \I1.REG_74l223r_adt_net_128394_\, 
        \I1.REG_74l225r_adt_net_128222_\, 
        \I1.REG_74l245r_adt_net_126207_\, 
        \I1.REG_74l246r_adt_net_126121_\, 
        \I1.REG_74l247r_adt_net_126035_\, 
        \I1.REG_74l248r_adt_net_125949_\, 
        \I1.REG_74l249r_adt_net_125863_\, 
        \I1.REG_74l250r_adt_net_125777_\, 
        \I1.REG_74l251r_adt_net_125691_\, 
        \I1.REG_74l252r_adt_net_125605_\, 
        \I1.REG_74l253r_adt_net_125400_\, 
        \I1.REG_74l254r_adt_net_125314_\, 
        \I1.REG_74l255r_adt_net_125228_\, 
        \I1.REG_74l256r_adt_net_125142_\, 
        \I1.REG_74l257r_adt_net_125056_\, 
        \I1.REG_74l258r_adt_net_124970_\, 
        \I1.REG_74l259r_adt_net_124884_\, 
        \I1.REG_74l260r_adt_net_124798_\, 
        \I1.REG_74l293r_adt_net_121470_\, 
        \I1.REG_74l294r_adt_net_121384_\, 
        \I1.REG_74l295r_adt_net_121298_\, 
        \I1.REG_74l296r_adt_net_121212_\, 
        \I1.REG_74l297r_adt_net_121126_\, 
        \I1.REG_74l298r_adt_net_121040_\, 
        \I1.REG_74l299r_adt_net_120954_\, 
        \I1.REG_74l300r_adt_net_120868_\, 
        \I1.REG_74l301r_adt_net_120782_\, 
        \I1.REG_74l302r_adt_net_120696_\, 
        \I1.REG_74l303r_adt_net_120610_\, 
        \I1.REG_74l304r_adt_net_120524_\, 
        \I1.REG_74l305r_adt_net_120438_\, 
        \I1.REG_74l306r_adt_net_120352_\, 
        \I1.REG_74l307r_adt_net_120266_\, 
        \I1.REG_74l308r_adt_net_120180_\, 
        \I1.REG_74l309r_adt_net_119991_\, 
        \I1.REG_74l310r_adt_net_119905_\, 
        \I1.REG_74l311r_adt_net_119819_\, 
        \I1.REG_74l312r_adt_net_119733_\, 
        \I1.REG_74l313r_adt_net_119647_\, 
        \I1.REG_74l314r_adt_net_119561_\, 
        \I1.REG_74l315r_adt_net_119475_\, 
        \I1.REG_74l316r_adt_net_119389_\, 
        \I1.REG_74l357r_adt_net_115127_\, 
        \I1.REG_74l358r_adt_net_115041_\, 
        \I1.REG_74l359r_adt_net_114955_\, 
        \I1.REG_74l360r_adt_net_114869_\, 
        \I1.REG_74l361r_adt_net_114783_\, 
        \I1.REG_74l362r_adt_net_114697_\, 
        \I1.REG_74l363r_adt_net_114611_\, 
        \I1.REG_74l364r_adt_net_114525_\, 
        \I1.REG_74l365r_adt_net_113912_\, 
        \I1.REG_74l366r_adt_net_113826_\, 
        \I1.REG_74l367r_adt_net_113740_\, 
        \I1.REG_74l368r_adt_net_113654_\, 
        \I1.REG_74l369r_adt_net_113568_\, 
        \I1.REG_74l370r_adt_net_113482_\, 
        \I1.REG_74l371r_adt_net_113396_\, 
        \I1.REG_74l372r_adt_net_113310_\, 
        \I1.REG_74l373r_adt_net_113087_\, 
        \I1.REG_74l374r_adt_net_113001_\, 
        \I1.REG_74l375r_adt_net_112915_\, 
        \I1.REG_74l376r_adt_net_112829_\, 
        \I1.REG_74l377r_adt_net_112743_\, 
        \I1.REG_74l378r_adt_net_112657_\, 
        \I1.REG_74l379r_adt_net_112571_\, 
        \I1.REG_74l380r_adt_net_112485_\, 
        \I1.REG_74l394r_adt_net_110698_\, \I1.N_628\, \I1.N_368\, 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r_adt_net_107364_\, 
        \I1.N_380\, \I1.N_598\, \I1.N_41\, \I1.N_49\, \I1.N_57\, 
        \I1.N_65\, \I1.N_280\, \I1.N_282\, \I1.N_1349\, 
        \I1.REG_74l213r\, \I1.REG_74l222r\, \I1.REG_74l224r\, 
        \I1.REG_74l226r\, \I1.REG_74l227r\, 
        \I1.REG_74l228r_net_1\, \I1.N_113\, \I1.REG_74l245r\, 
        \I1.REG_74l246r\, \I1.REG_74l247r\, \I1.REG_74l248r\, 
        \I1.REG_74l249r\, \I1.REG_74l250r\, \I1.REG_74l251r\, 
        \I1.REG_74l252r\, \I1.REG_74l253r\, \I1.REG_74l254r\, 
        \I1.REG_74l255r\, \I1.REG_74l256r\, \I1.REG_74l257r\, 
        \I1.REG_74l258r\, \I1.REG_74l259r\, \I1.REG_74l260r\, 
        \I1.N_137\, \I1.N_145\, \I1.N_185\, \I1.N_193\, 
        \I1.REG_74_0l332r\, \I1.N_201\, \I1.N_209\, \I1.N_661\, 
        \I1.REG_74l365r\, \I1.REG_74l366r\, \I1.REG_74l367r\, 
        \I1.REG_74l368r\, \I1.REG_74l369r\, \I1.REG_74l370r\, 
        \I1.REG_74l371r\, \I1.REG_74l372r\, \I1.REG_74l373r\, 
        \I1.REG_74l374r\, \I1.REG_74l375r\, \I1.REG_74l376r\, 
        \I1.REG_74l377r\, \I1.REG_74l378r\, \I1.REG_74l379r\, 
        \I1.REG_74l380r_net_1\, \I1.REG_74l394r\, \I1.N_1162\, 
        \I1.N_79\, \I1.N_77\, \I1.N_75\, \I1.N_1381\, 
        \I1.BYTECNT_n3\, \I1.N_174\, \I1.N_1161\, \I1.BYTECNT_n0\, 
        \I1.N_389_i_i_0\, \I1.N_1378\, \I1.LOAD_RES_i_0\, 
        \I1.REG_74l221r\, \I1.REG_74l223r\, \I1.REG_74l225r\, 
        \I1.REG_74l189r\, \I1.REG_74l191r_adt_net_131355_\, 
        \I1.REG_74l194r_adt_net_131097_\, \I1.REG_74l309r\, 
        \I1.REG_74l310r\, \I1.REG_74l311r\, \I1.REG_74l312r\, 
        \I1.REG_74l313r\, \I1.REG_74l314r\, \I1.REG_74l315r\, 
        \I1.REG_74l316r_net_1\, \I1.REG_74l317r\, 
        \I1.REG_74l318r\, \I1.REG_74l319r\, \I1.REG_74l320r\, 
        \I1.REG_74l321r\, \I1.REG_74l322r\, \I1.REG_74l323r\, 
        \I1.REG_74l324r_net_1\, \I1.REG_74l357r\, 
        \I1.REG_74l358r\, \I1.REG_74l359r\, \I1.REG_74l360r\, 
        \I1.REG_74l361r\, \I1.REG_74l362r\, \I1.REG_74l363r\, 
        \I1.REG_74l364r\, \I1.PAGECNT_320_net_1\, 
        \I1.REG_1_129_net_1\, \I1.REG_1_128_net_1\, 
        \I1.REG_1_127_net_1\, \I1.REG_1_125_net_1\, 
        \I1.REG_1_123_net_1\, \I1.N_463_1\, \I1.N_362\, 
        \I1.N_406\, \I1.N_1385\, \I1.N_603_i\, \I1.N_1386\, 
        \I1.REG_74l173r_adt_net_132940_\, 
        \I1.REG_74l176r_adt_net_132682_\, 
        \I1.REG_74l179r_adt_net_132424_\, 
        \I1.REG_74l180r_adt_net_132338_\, 
        \I1.N_68_adt_net_108395_\, 
        \I1.un1_sbyte13_i_i_i_1_adt_net_108267_\, 
        \I1.N_1193_adt_net_1562__net_1\, \I1.REG_74l165r\, 
        \I1.REG_74l166r\, \I1.REG_74l167r\, \I1.REG_74l168r\, 
        \I1.REG_74l169r\, \I1.REG_74l170r\, \I1.REG_74l171r\, 
        \I1.REG_74l172r_net_1\, \I1.REG_74l174r\, 
        \I1.REG_74l175r\, \I1.REG_74l177r\, \I1.REG_74l178r\, 
        \I1.REG_74l181r\, \I1.REG_74l182r\, \I1.REG_74l183r\, 
        \I1.REG_74l184r\, \I1.REG_74l185r\, \I1.REG_74l186r\, 
        \I1.REG_74l187r\, \I1.REG_74l188r_net_1\, \I1.N_129\, 
        \I1.N_1337\, \I1.N_1338\, \I1.N_1339\, \I1.N_1340\, 
        \I1.N_1341\, \I1.N_1342\, \I1.N_1343\, 
        \I1.REG_1_106_net_1\, \I1.REG_1_107_net_1\, \I1.N_1346\, 
        \I1.N_1347\, \I1.N_1348\, \I1.REG_1_111_net_1\, 
        \I1.N_144\, \I1.N_1350\, \I1.REG_1_114_net_1\, 
        \I1.REG_74l214r\, \I1.REG_74l215r\, \I1.REG_74l216r\, 
        \I1.REG_74l217r\, \I1.REG_74l218r\, \I1.REG_74l219r\, 
        \I1.REG_74l220r_net_1\, \I1.REG_74l229r\, 
        \I1.REG_74l230r\, \I1.REG_74l231r\, \I1.REG_74l232r\, 
        \I1.REG_74l233r\, \I1.REG_74l234r\, \I1.REG_74l235r\, 
        \I1.REG_74l236r_net_1\, \I1.REG_74l237r\, 
        \I1.REG_74l238r\, \I1.REG_74l239r\, \I1.REG_74l240r\, 
        \I1.REG_74l241r\, \I1.REG_74l242r\, \I1.REG_74l243r\, 
        \I1.REG_74l244r_net_1\, \I1.REG_1_146_net_1\, 
        \I1.REG_1_147_net_1\, \I1.REG_1_148_net_1\, 
        \I1.REG_1_149_net_1\, \I1.REG_1_150_net_1\, 
        \I1.REG_1_151_net_1\, \I1.REG_1_152_net_1\, 
        \I1.REG_1_153_net_1\, \I1.REG_1_154_net_1\, 
        \I1.REG_1_155_net_1\, \I1.REG_1_156_net_1\, 
        \I1.REG_1_157_net_1\, \I1.REG_1_158_net_1\, 
        \I1.REG_1_159_net_1\, \I1.REG_1_160_net_1\, 
        \I1.REG_1_161_net_1\, \I1.REG_74l277r\, 
        \I1.REG_1_178_net_1\, \I1.REG_74l278r\, 
        \I1.REG_1_179_net_1\, \I1.REG_74l279r\, 
        \I1.REG_1_180_net_1\, \I1.REG_74l280r\, 
        \I1.REG_1_181_net_1\, \I1.REG_74l281r\, 
        \I1.REG_1_182_net_1\, \I1.REG_74l282r\, 
        \I1.REG_1_183_net_1\, \I1.REG_74l283r\, 
        \I1.REG_1_184_net_1\, \I1.REG_74l284r_net_1\, 
        \I1.REG_1_185_net_1\, \I1.REG_74l285r\, 
        \I1.REG_1_186_net_1\, \I1.REG_74l286r\, 
        \I1.REG_1_187_net_1\, \I1.REG_74l287r\, 
        \I1.REG_1_188_net_1\, \I1.REG_74l288r\, 
        \I1.REG_1_189_net_1\, \I1.REG_74l289r\, 
        \I1.REG_1_190_net_1\, \I1.REG_74l290r\, 
        \I1.REG_1_191_net_1\, \I1.REG_74l291r\, 
        \I1.REG_1_192_net_1\, \I1.REG_74l292r_net_1\, 
        \I1.REG_1_193_net_1\, \I1.REG_74l293r\, \I1.REG_74l294r\, 
        \I1.REG_74l295r\, \I1.REG_74l296r\, \I1.REG_74l297r\, 
        \I1.REG_74l298r\, \I1.REG_74l299r\, 
        \I1.REG_74l300r_net_1\, \I1.REG_74l301r\, 
        \I1.REG_74l302r\, \I1.REG_74l303r\, \I1.REG_74l304r\, 
        \I1.REG_74l305r\, \I1.REG_74l306r\, \I1.REG_74l307r\, 
        \I1.REG_74l308r_net_1\, \I1.REG_74l341r\, 
        \I1.REG_74l342r\, \I1.REG_74l343r\, \I1.REG_74l344r\, 
        \I1.REG_74l345r\, \I1.REG_74l346r\, \I1.REG_74l347r\, 
        \I1.REG_74l348r_net_1\, \I1.REG_74l349r\, 
        \I1.REG_74l350r\, \I1.REG_74l351r\, \I1.REG_74l352r\, 
        \I1.REG_74l353r\, \I1.REG_74l354r\, \I1.REG_74l355r\, 
        \I1.REG_74l356r_net_1\, \I1.REG_1_266_net_1\, 
        \I1.REG_1_267_net_1\, \I1.REG_1_268_net_1\, 
        \I1.REG_1_269_net_1\, \I1.REG_1_270_net_1\, 
        \I1.REG_1_271_net_1\, \I1.REG_1_272_net_1\, 
        \I1.REG_1_273_net_1\, \I1.REG_1_274_net_1\, 
        \I1.REG_1_275_net_1\, \I1.REG_1_276_net_1\, 
        \I1.REG_1_277_net_1\, \I1.REG_1_278_net_1\, 
        \I1.REG_1_279_net_1\, \I1.REG_1_280_net_1\, 
        \I1.REG_1_281_net_1\, \I1.REG_74l381r\, \I1.REG_74l382r\, 
        \I1.REG_74l383r\, \I1.REG_74l384r\, \I1.REG_74l385r\, 
        \I1.REG_74l386r\, \I1.REG_74l387r\, 
        \I1.REG_74l388r_net_1\, \I1.REG_74l389r\, 
        \I1.REG_1_290_net_1\, \I1.REG_74l390r\, 
        \I1.REG_1_291_net_1\, \I1.REG_74l391r\, 
        \I1.REG_1_292_net_1\, \I1.REG_74l392r\, 
        \I1.REG_1_293_net_1\, \I1.REG_74l393r\, 
        \I1.REG_1_294_net_1\, \I1.REG_1_295_net_1\, 
        \I1.REG_74l395r\, \I1.REG_1_296_net_1\, 
        \I1.REG_74l396r_net_1\, \I1.REG_1_297_net_1\, 
        \I1.REG_74l397r\, \I1.REG_1_298_net_1\, \I1.REG_74l398r\, 
        \I1.REG_1_299_net_1\, \I1.REG_74l399r\, 
        \I1.REG_1_300_net_1\, \I1.REG_74l400r\, 
        \I1.REG_1_301_net_1\, \I1.REG_74l401r\, 
        \I1.REG_1_302_net_1\, \I1.REG_74l402r\, 
        \I1.REG_1_303_net_1\, \I1.REG_74l403r\, 
        \I1.REG_1_304_net_1\, \I1.REG_74l404r_net_1\, 
        \I1.REG_1_305_net_1\, \I1.BYTECNT_306_net_1\, 
        \I1.BYTECNT_307_net_1\, \I1.BYTECNT_308_net_1\, 
        \I1.BYTECNT_309_net_1\, \I1.BYTECNT_310_net_1\, 
        \I1.N_304_adt_net_105325_Ra1_\, \I1.BYTECNT_311_net_1\, 
        \I1.BYTECNT_312_net_1\, \I1.BYTECNT_313_net_1\, 
        \I1.BYTECNT_314_net_1\, \I1.un1_sbyte13_i_i_i_1_net_1\, 
        \I1.N_1380\, \I1.PAGECNT_318_net_1\, \I1.N_1379\, 
        \I1.PAGECNT_319_net_1\, \I1.N_1377\, 
        \I1.PAGECNT_321_net_1\, \I1.PAGECNT_n5\, 
        \I1.PAGECNT_322_net_1\, \I1.PAGECNT_n4\, \I1.PAGECNT_n3\, 
        \I1.PAGECNT_n2\, \I1.PAGECNT_n1\, \I1.PAGECNT_n0\, 
        \I1.PAGECNT_327_net_1\, \I1.PAGECNT_326_net_1\, 
        \I1.PAGECNT_325_net_1\, \I1.PAGECNT_324_net_1\, 
        \I1.PAGECNT_323_net_1\, \I1.REG_1_209_net_1\, 
        \I1.REG_1_208_net_1\, \I1.REG_1_207_net_1\, 
        \I1.REG_1_206_net_1\, \I1.REG_1_205_net_1\, 
        \I1.REG_1_204_net_1\, \I1.REG_1_203_net_1\, 
        \I1.REG_1_202_net_1\, \I1.REG_1_201_net_1\, 
        \I1.REG_1_200_net_1\, \I1.REG_1_199_net_1\, 
        \I1.REG_1_198_net_1\, \I1.REG_1_197_net_1\, 
        \I1.REG_1_196_net_1\, \I1.REG_1_195_net_1\, 
        \I1.REG_1_194_net_1\, \I1.N_50_0_adt_net_109756__net_1\, 
        \I1.REG_1_289_net_1\, \I1.REG_1_288_net_1\, 
        \I1.REG_1_287_net_1\, \I1.REG_1_286_net_1\, 
        \I1.REG_1_285_net_1\, \I1.REG_1_284_net_1\, 
        \I1.REG_1_283_net_1\, \I1.REG_1_282_net_1\, 
        \I1.REG_1_242_net_1\, \I1.REG_1_243_net_1\, 
        \I1.REG_1_244_net_1\, \I1.REG_1_245_net_1\, 
        \I1.REG_1_246_net_1\, \I1.REG_1_247_net_1\, 
        \I1.REG_1_248_net_1\, \I1.REG_1_249_net_1\, 
        \I1.REG_1_250_net_1\, \I1.REG_1_251_net_1\, 
        \I1.REG_1_252_net_1\, \I1.REG_1_253_net_1\, 
        \I1.REG_1_254_net_1\, \I1.REG_1_255_net_1\, 
        \I1.REG_1_256_net_1\, \I1.REG_1_257_net_1\, 
        \I1.REG_1_115_net_1\, \I1.REG_1_116_net_1\, 
        \I1.REG_1_117_net_1\, \I1.REG_1_118_net_1\, 
        \I1.REG_1_119_net_1\, \I1.REG_1_120_net_1\, 
        \I1.REG_1_121_net_1\, \I1.REG_1_122_net_1\, 
        \I1.REG_1_124_net_1\, \I1.REG_1_126_net_1\, 
        \I1.REG_74l262r_adt_net_124543_\, 
        \I1.REG_74l264r_adt_net_124371_\, 
        \I1.REG_74l269r_adt_net_123904_\, 
        \I1.REG_74l271r_adt_net_123732_\, 
        \I1.REG_74l273r_adt_net_123560_\, 
        \I1.N_321_adt_net_105403_\, \I1.N_333_Ra1_\, 
        \I1.REG_1_66_net_1\, \I1.REG_1_67_net_1\, 
        \I1.REG_1_68_net_1\, \I1.REG_1_69_net_1\, 
        \I1.REG_1_70_net_1\, \I1.REG_1_71_net_1\, 
        \I1.REG_1_72_net_1\, \I1.REG_1_73_net_1\, 
        \I1.REG_74l173r\, \I1.REG_1_74_net_1\, 
        \I1.REG_1_75_net_1\, \I1.REG_1_76_net_1\, 
        \I1.REG_74l176r\, \I1.REG_1_77_net_1\, 
        \I1.REG_1_78_net_1\, \I1.REG_1_79_net_1\, 
        \I1.REG_74l179r\, \I1.REG_1_80_net_1\, 
        \I1.REG_74l180r_net_1\, \I1.REG_1_81_net_1\, 
        \I1.REG_1_82_net_1\, \I1.REG_1_83_net_1\, 
        \I1.REG_1_84_net_1\, \I1.REG_1_85_net_1\, 
        \I1.REG_1_86_net_1\, \I1.REG_1_87_net_1\, 
        \I1.REG_1_88_net_1\, \I1.REG_1_89_net_1\, 
        \I1.REG_1_90_net_1\, \I1.REG_74l190r\, 
        \I1.REG_1_91_net_1\, \I1.REG_74l191r\, 
        \I1.REG_1_92_net_1\, \I1.REG_74l192r\, 
        \I1.REG_1_93_net_1\, \I1.REG_74l193r\, 
        \I1.REG_1_94_net_1\, \I1.REG_74l194r\, 
        \I1.REG_1_95_net_1\, \I1.REG_74l195r\, 
        \I1.REG_1_96_net_1\, \I1.REG_74l196r_net_1\, 
        \I1.REG_1_97_net_1\, \I1.REG_1_98_net_1\, 
        \I1.REG_1_99_net_1\, \I1.REG_1_100_net_1\, 
        \I1.REG_1_101_net_1\, \I1.REG_1_102_net_1\, 
        \I1.REG_1_103_net_1\, \I1.REG_1_104_net_1\, 
        \I1.REG_1_105_net_1\, \I1.REG_1_108_net_1\, 
        \I1.REG_1_109_net_1\, \I1.REG_1_110_net_1\, 
        \I1.REG_1_112_net_1\, \I1.REG_1_113_net_1\, 
        \I1.REG_1_130_net_1\, \I1.REG_1_131_net_1\, 
        \I1.REG_1_132_net_1\, \I1.REG_1_133_net_1\, 
        \I1.REG_1_134_net_1\, \I1.REG_1_135_net_1\, 
        \I1.REG_1_136_net_1\, \I1.REG_1_137_net_1\, 
        \I1.REG_1_138_net_1\, \I1.REG_1_139_net_1\, 
        \I1.REG_1_140_net_1\, \I1.REG_1_141_net_1\, 
        \I1.REG_1_142_net_1\, \I1.REG_1_143_net_1\, 
        \I1.REG_1_144_net_1\, \I1.REG_1_145_net_1\, 
        \I1.REG_74l261r\, \I1.REG_1_162_net_1\, \I1.REG_74l262r\, 
        \I1.REG_1_163_net_1\, \I1.REG_74l263r\, 
        \I1.REG_1_164_net_1\, \I1.REG_74l264r\, 
        \I1.REG_1_165_net_1\, \I1.REG_74l265r\, 
        \I1.REG_1_166_net_1\, \I1.REG_74l266r\, 
        \I1.REG_1_167_net_1\, \I1.REG_74l267r\, 
        \I1.REG_1_168_net_1\, \I1.REG_74l268r_net_1\, 
        \I1.REG_1_169_net_1\, \I1.REG_74l269r\, 
        \I1.REG_1_170_net_1\, \I1.REG_74l270r\, 
        \I1.REG_1_171_net_1\, \I1.REG_74l271r\, 
        \I1.REG_1_172_net_1\, \I1.REG_74l272r\, 
        \I1.REG_1_173_net_1\, \I1.REG_74l273r\, 
        \I1.REG_1_174_net_1\, \I1.REG_74l274r\, 
        \I1.REG_1_175_net_1\, \I1.REG_74l275r\, 
        \I1.REG_1_176_net_1\, \I1.REG_74l276r_net_1\, 
        \I1.REG_1_177_net_1\, \I1.REG_1_210_net_1\, 
        \I1.REG_1_211_net_1\, \I1.REG_1_212_net_1\, 
        \I1.REG_1_213_net_1\, \I1.REG_1_214_net_1\, 
        \I1.REG_1_215_net_1\, \I1.REG_1_216_net_1\, 
        \I1.REG_1_217_net_1\, \I1.REG_1_218_net_1\, 
        \I1.REG_1_219_net_1\, \I1.REG_1_220_net_1\, 
        \I1.REG_1_221_net_1\, \I1.REG_1_222_net_1\, 
        \I1.REG_1_223_net_1\, \I1.REG_1_224_net_1\, 
        \I1.REG_1_225_net_1\, \I1.REG_74l325r\, \I1.REG_74l326r\, 
        \I1.REG_74l327r\, \I1.REG_74l328r\, \I1.REG_74l329r\, 
        \I1.REG_74l330r\, \I1.REG_74l331r\, 
        \I1.REG_74l332r_net_1\, \I1.REG_74l333r\, 
        \I1.REG_74l334r\, \I1.REG_74l335r\, \I1.REG_74l336r\, 
        \I1.REG_74l337r\, \I1.REG_74l338r\, \I1.REG_74l339r\, 
        \I1.REG_74l340r_net_1\, \I1.REG_1_258_net_1\, 
        \I1.REG_1_259_net_1\, \I1.REG_1_260_net_1\, 
        \I1.REG_1_261_net_1\, \I1.REG_1_262_net_1\, 
        \I1.REG_1_263_net_1\, \I1.REG_1_264_net_1\, 
        \I1.REG_1_265_net_1\, \I1.N_332\, \I1.N_386_i_i_0\, 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\, 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Ra1_\, 
        \I1.N_304_Ra1_\, \I1.N_174_adt_net_108976_\, 
        \I1.N_317_Ra1_\, \I1.N_299_Ra1_\, 
        \I1.REG_74_12_220_m9_i_a6_0\, \I1.N_323\, \I1.N_300_Ra1_\, 
        \I1.N_232_1\, \I1.N_237\, \I1.REG_1_226_net_1\, 
        \I1.REG_1_227_net_1\, \I1.REG_1_228_net_1\, 
        \I1.REG_1_229_net_1\, \I1.REG_1_230_net_1\, 
        \I1.REG_1_231_net_1\, \I1.REG_1_232_net_1\, 
        \I1.REG_1_233_net_1\, \I1.REG_1_234_net_1\, 
        \I1.REG_1_235_net_1\, \I1.REG_1_236_net_1\, 
        \I1.REG_1_237_net_1\, \I1.REG_1_238_net_1\, 
        \I1.REG_1_239_net_1\, \I1.REG_1_240_net_1\, 
        \I1.REG_1_241_net_1\, \I1.N_327\, \I1.REG_74_1_a0_0l228r\, 
        \I1.N_392_i\, \I1.N_1381_adt_net_109130_\, 
        \I1.REG_74_0_iv_0_0_o2_245_m6_i_0_tz_i_adt_net_1555__net_1\, 
        \I1.REG_15_sqmuxa_adt_net_1457__net_1\, \I1.N_305_Ra1_\, 
        \I1.N_321\, \I1.N_223_adt_net_108706_\, \I1.N_1169\, 
        \I1.REG_74_5_404_m1_e_0_net_1\, \I1.N_590\, \I1.N_267\, 
        \I1.N_253\, \I1.REG_74_1_i_a2_a0_2l404r\, \I1.N_127_i\, 
        \I1.REG_74_1_380_N_16\, \I1.N_334\, \I1.N_591_1\, 
        \I1.N_390_i_i_0_i\, \I1.N_388_i_0_i\, \I1.N_308_Ra1_\, 
        \I1.N_393_i_i_0_i\, \I1.N_330_i_0_i\, \I1.N_260\, 
        \I1.REG_74_9_0_o4_a0_2l372r\, \I1.N_346\, 
        \I1.REG_74_13_388_N_16_adt_net_109531_\, 
        \I1.REG_74_3_4_il380r_adt_net_123086_\, 
        \I1.REG_74_8_308_m9_i_1\, 
        \I1.REG_74_2_2_il340r_adt_net_117061_\, 
        \I1.REG_74_2_4_il228r_adt_net_115250_\, 
        \I1.N_1367_i_adt_net_112072_\, \I1.N_75_adt_net_109200_\, 
        \I1.N_223_adt_net_108707_\, 
        \I1.REG_74_12_300_N_15_adt_net_3731__net_1\, 
        \I1.REG_74_4_i_a2_404_N_4_i_adt_net_1465__net_1\, 
        \I1.N_311_i_i_Ra1_\, \I1.N_273_5_i\, \I1.REG_15_sqmuxa\, 
        \I1.REG_16_sqmuxa\, \I1.REG_74_1_396_m7_i_3\, \I1.N_259\, 
        \I1.N_255\, \I1.REG_74_8_0_324_m6_e_net_1\, \I1.N_243\, 
        \I1.REG_74_8_1_tzl340r_net_1\, \I1.REG_74_1_396_N_12\, 
        \I1.N_335\, \I1.N_394_i_i_0_i\, \I1.N_310_Ra1_\, 
        \I2.N303\, \I5.DATA_1_sqmuxa_2\, \I5.sstate1_ns_el11r\, 
        \I2.DTE_1l28r\, \I5.sstate1l2r_net_1\, 
        \I2.DTE_1l28r_Rd1__net_1\, \I2.DTE_21_1l28r_Rd1__net_1\, 
        \I3.TCNT3_i_0_il6r_net_1\, \TICKl1r\, \I3.TCNT3l7r_net_1\, 
        \I3.TCNT3l5r_net_1\, \I3.TCNT2_i_0_il6r_net_1\, 
        \I3.TCNT2l7r_net_1\, \I3.TCNT2l5r_net_1\, 
        \I5.sstate1l4r_net_1\, \I5.sstate1l10r_net_1\, \TICKl3r\, 
        \I5.sstate1l3r_net_1\, \I4.bcnt_i_0_il2r_net_1\, 
        \LSRAM_FL_RADDRl2r\, \I4.bcntl1r_net_1\, 
        \LSRAM_FL_RADDRl1r\, \I4.bcntl0r_net_1\, 
        \LSRAM_FL_RADDRl0r\, \I0.BNC_RESF2_net_1\, 
        \I0.EV_RESF2_net_1\, \I2.TRAIL_MIS7_i_net_1\, 
        \I2.LSRAM_FL_RD7_net_1\, \I2.STATE5l1r_net_1\, 
        \I2.STATE5l2r_net_1\, \I2.EVNT_NUM_c1_net_1\, \I2.N_187\, 
        \I2.TDCDASl30r_net_1\, \I2.TDCDBSl30r_net_1\, 
        \I2.TDCDASl18r_net_1\, \I2.TDCDBSl18r_net_1\, 
        \I2.TDCDASl17r_net_1\, \I2.TDCDBSl17r_net_1\, 
        \I2.TDCDASl16r_net_1\, \I2.TDCDBSl16r_net_1\, 
        \I2.TDCDASl15r_net_1\, \I2.TDCDBSl15r_net_1\, 
        \I2.TDCDASl14r_net_1\, \I2.TDCDBSl14r_net_1\, 
        \I2.TDCDBSl13r_net_1\, \I2.TDCDASl13r_net_1\, 
        \I2.TDCDBSl12r_net_1\, \I2.TDCDASl12r_net_1\, 
        \I2.TDCDBSl11r_net_1\, \I2.TDCDASl11r_net_1\, 
        \I2.TDCDBSl10r_net_1\, \I2.TDCDASl10r_net_1\, 
        \I2.TDCDBSl9r_net_1\, \I2.TDCDASl9r_net_1\, 
        \I2.TDCDBSl8r_net_1\, \I2.TDCDASl8r_net_1\, 
        \I2.STATE2l4r_net_1\, \I2.STATE2l3r_net_1\, 
        \I2.RAMDT4l4r_net_1\, \I2.RAMDT4l11r_net_1\, 
        \I2.RAMDT4l3r_net_1\, \I2.RAMDT4l10r_net_1\, 
        \I2.RAMDT4l2r_net_1\, \I2.RAMDT4l9r_net_1\, 
        \I2.RAMDT4l1r_net_1\, \I2.RAMDT4l8r_net_1\, 
        \I2.RAMDT4l0r_net_1\, \I2.RAMDT4l7r_net_1\, \I2.N_622\, 
        \I2.N_625\, \I2.N_633\, \I2.L2AF2_net_1\, \I2.N247\, 
        \I2.CHAIN_ERRS_net_1\, \I2.MTDIAS_net_1\, 
        \I2.END_TDC5_net_1\, \I2.N_3830\, \I2.N_3829\, 
        \I2.REG_1_n0_net_1\, \I2.TDCDRYBS_net_1\, 
        \I2.TDCDRYAS_net_1\, \I1.N_300_Rd1__net_1\, 
        \I1.N_305_Rd1__net_1\, \I1.N_308_Rd1__net_1\, 
        \I1.PAGECNT_0l9r_adt_net_835132_Rd1__net_1\, 
        \I1.PAGECNTl9r_net_1\, \I3.TCNT1l0r_net_1\, 
        \I3.TCNT2_i_0_il0r_net_1\, \I3.TCNT2l1r_net_1\, 
        \I3.TCNT2_i_0_il2r_net_1\, \I3.TCNT2l3r_net_1\, 
        \I3.TCNT2_i_0_il4r_net_1\, \I3.TCNT4_i_0_il0r_net_1\, 
        \I3.TICKl2r_net_1\, \I3.TCNT4l1r_net_1\, 
        \I3.TCNT4_i_0_il2r_net_1\, \I3.TCNT4l3r_net_1\, 
        \I3.TCNT3_i_0_il0r_net_1\, \I3.TCNT3l1r_net_1\, 
        \I3.TCNT3_i_0_il2r_net_1\, \I3.TCNT3l3r_net_1\, 
        \I3.TCNT3_i_0_il4r_net_1\, \I3.N_311\, \I3.N_277\, 
        \I3.TCNT1l5r_net_1\, \I3.TCNT1l4r_net_1\, 
        \I3.TCNT1_i_0_il3r_net_1\, \I3.TCNT1l2r_net_1\, 
        \I3.TCNT1_i_0_il1r_net_1\, \I3.N_547\, 
        \I1.PAGECNT_0l8r_adt_net_834720__adt_net_835724_Rd1__net_1\, 
        \I5.sstate1l9r_net_1\, \I2.TDCDASl29r_net_1\, 
        \I2.N_3016_adt_net_24530_\, \I2.N295_adt_net_68996_\, 
        \I2.N311_adt_net_69399_\, \I2.N_3832_adt_net_101495_\, 
        \I2.N_3832_adt_net_101536_\, \I1.PAGECNTl5r_net_1\, 
        \I1.PAGECNTl6r_net_1\, \I3.REGMAPl57r_net_1\, 
        \I3.REGMAPl39r_net_1\, \I3.REGMAP_i_0_il38r_net_1\, 
        \I1.PAGECNTl0r_adt_net_833884_Rd1__net_1\, 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__net_1\, 
        \I3.REGMAPl16r_net_1\, \I3.REGMAPl43r_net_1\, 
        \I3.REGMAPl34r_net_1\, \I3.REGMAP_i_il46r_net_1\, 
        \I3.REGMAPl47r_net_1\, \I3.REGMAPl35r_net_1\, 
        \I3.REGMAP_i_0_il36r_net_1\, \I3.REGMAPl37r_net_1\, 
        \I3.REGMAP_i_0_il40r_net_1\, \I3.REGMAPl41r_net_1\, 
        \I3.REGMAP_i_0_il42r_net_1\, \I3.REGMAPl44r_net_1\, 
        \I3.REGMAP_i_0_il45r_net_1\, \I3.REGMAPl29r_net_1\, 
        \I3.REGMAP_i_0_il30r_net_1\, \I3.REGMAPl31r_net_1\, 
        \I3.REGMAP_i_0_il32r_net_1\, \I3.REGMAPl22r_net_1\, 
        \I3.REGMAPl25r_net_1\, \I3.REGMAPl26r_net_1\, 
        \I3.REGMAPl27r_net_1\, \I3.REGMAP_i_0_il19r_net_1\, 
        \I3.REGMAPl28r_net_1\, \I3.REGMAPl23r_net_1\, 
        \I3.REGMAP_i_0_il24r_net_1\, \I3.REGMAPl18r_net_1\, 
        \I3.REGMAPl21r_net_1\, \I3.REGMAPl20r_net_1\, 
        \I3.STATE1_ipl2r_net_1\, \I2.G_EVNT_NUM_i_0_il0r_net_1\, 
        \I3.TCNT2_c1\, \I5.N_65\, \I4.bcntl3r_net_1\, 
        \I2.MIC_REG2l3r_adt_net_834020_Rd1__net_1\, 
        \I2.sram_empty_0_i_0_i\, \I2.sram_empty_1_i_0_i\, 
        \I2.sram_empty_2_i_0_i\, \I2.un21_sram_empty_2_net_1\, 
        \I2.un21_sram_empty_3_net_1\, \I2.L2AF3_net_1\, 
        \I2.RAMDT4l6r_net_1\, \I2.RAMDT4l13r_net_1\, \I2.N_4543\, 
        \I2.N_4544\, \I2.N_215\, \I2.STATE3l0r_net_1\, 
        \I2.STATE3l4r_net_1\, \I2.MIC_REG3l7r_net_1\, 
        \I2.MIC_REG3l6r_net_1\, \I2.MIC_REG3l5r_net_1\, 
        \I2.MIC_REG3l4r_net_1\, \I2.MIC_REG3l1r_net_1\, 
        \I2.MIC_REG3l0r_net_1\, \I2.MIC_REG2l7r_net_1\, 
        \I2.MIC_REG2l6r_net_1\, \I2.MIC_REG2_i_0_il5r_net_1\, 
        \I2.MIC_REG2_i_0_il4r_net_1\, \I2.MIC_REG2l1r_net_1\, 
        \I2.MIC_REG2l0r_net_1\, \I2.MIC_REG1l7r_net_1\, 
        \I2.MIC_REG1_i_il6r_net_1\, \I2.MIC_REG1l5r_net_1\, 
        \I2.MIC_REG1l4r_net_1\, \I2.MIC_REG1l1r_net_1\, 
        \I2.MIC_REG1l0r_net_1\, \I2.G_1\, \I2.N_3545_i_i\, 
        \I2.G_1_0\, \I2.N_3543_i_i\, \I2.G_1_1\, \I2.N_3541_i_i\, 
        \I1.PAGECNTl8r_net_1\, \I1.N_254\, 
        \I3.STATE1_ipl0r_net_1\, \I3.STATE1_ipl3r_net_1\, 
        \I3.REGMAPl55r_net_1\, \I3.REGMAPl17r_net_1\, \I3.N_2014\, 
        \I3.N_203\, \I2.REG_0l3r_adt_net_848__net_1\, 
        \I2.N_3834_i_0_adt_net_1384__net_1\, 
        \I2.MIC_REG1l3r_adt_net_834596_Rd1__net_1\, 
        \I2.N_4551_adt_net_63747_\, \I2.N_4551_adt_net_63757_\, 
        \I2.PIPE7_DTl26r_net_1\, \I1.N_323_adt_net_108906_\, 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__net_1\, 
        \I2.PIPE7_DTl27r_net_1\, 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Rd1__net_1\, 
        \I3.REGMAPl9r_net_1\, \I3.REGMAPl7r_net_1\, 
        \I3.REGMAPl33r_net_1\, \I3.LWORDS_net_1\, 
        \I2.MIC_REG3l2r_net_1\, \I2.MIC_REG2l2r_net_1\, 
        \I2.MIC_REG1l2r_net_1\, \I1.N_355\, \I1.N_317_Rd1__net_1\, 
        \I4.N_48_3_adt_net_14719_\, \I2.PIPE3_DTl8r_net_1\, 
        \I3.N_58_i_0_adt_net_134395_\, 
        \I3.N_2083_adt_net_134513_\, \I3.N_2086_adt_net_134541_\, 
        \I3.N_177_adt_net_134570_\, \I4.N_7\, 
        \I2.TRGSERVl0r_net_1\, \I2.TRGSERVl1r_net_1\, 
        \I2.PIPE4_DTl9r_net_1\, \I2.PIPE4_DT_i_il1r_net_1\, 
        \I2.N_85\, \I2.MIC_REG3_320_net_1\, 
        \I2.MIC_REG2_312_net_1\, \I2.MIC_REG1_304_net_1\, 
        \I2.N357_adt_net_54497_\, \I2.N357_adt_net_54538_\, 
        \I2.N357_0_adt_net_55523_\, 
        \I2.N_2358_tz_tz_adt_net_55567_\, \I2.PIPE4_DTl10r_net_1\, 
        \I2.PIPE4_DTl4r_net_1\, \I2.PIPE4_DTl6r_net_1\, 
        \I2.PIPE4_DTl5r_net_1\, \I2.N_112_1\, 
        \I2.DWACT_ADD_CI_0_TMP_0l0r\, \I2.PIPE4_DTl7r_net_1\, 
        \I2.RAMDT4l5r_net_1\, \I2.N_72_0\, \I2.N_89\, \I2.N_64\, 
        \I2.N_28\, \I2.PIPE4_DTl3r_net_1\, \I2.N_67\, \I2.N_17_0\, 
        \I2.RAMDT4l12r_net_1\, \I3.N_203_adt_net_24461_\, 
        \I2.PIPE4_DTl8r_net_1\, \I3.REGMAP_i_0_il58r_net_1\, 
        \I3.N_545_adt_net_165680_\, \I2.MIC_REG3l3r_net_1\, 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_o2tt_N_8_Rd1__net_1\, 
        \I1.N_349_Rd1__net_1\, 
        \I1.REG_74_1_380_m8_i_0_Rd1__net_1\, 
        \I1.REG_74_2_0l404r_Rd1__net_1\, \I1.N_238_Rd1__net_1\, 
        \I1.N_268_Rd1__net_1\, \I1.REG_74_12_300_N_13_Rd1__net_1\, 
        \I1.N_341_Rd1__net_1\, \I1.N_606_Rd1__net_1\, 
        \I3.N_264_0_adt_net_1653_Rd1__net_1\, 
        \I2.REG_0l3r_adt_net_19771_Rd1__net_1\, 
        \I2.REG_0l3r_adt_net_19773_Rd1__net_1\, 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_adt_net_19883_Rd1__net_1\, 
        \I1.N_591_1_adt_net_106236_Rd1__net_1\, 
        \I1.REG_15_sqmuxa_adt_net_109461_Rd1__net_1\, 
        \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Rd1__net_1\, 
        \PULSE_0l0r_adt_net_834380_Rd1__net_1\, 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__net_1\, 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Ra1_\, 
        \I2.DTE_0_sqmuxa_i_o2tt_N_8_Ra1_\, \I1.N_349_Ra1_\, 
        \I1.REG_74_1_380_m8_i_0_Ra1_\, \I1.REG_74_2_0l404r_Ra1_\, 
        \I1.N_238_Ra1_\, \I1.N_268_Ra1_\, 
        \I1.REG_74_12_300_N_13_Ra1_\, \I1.N_341_Ra1_\, 
        \I1.N_606_Ra1_\, \I3.N_264_0_adt_net_1653_Ra1__net_1\, 
        \I2.REG_0l3r_adt_net_19771_Ra1__net_1\, 
        \I2.REG_0l3r_adt_net_19773_Ra1__net_1\, 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_adt_net_19883_Ra1_\, 
        \I1.N_591_1_adt_net_106236_Ra1_\, 
        \I1.REG_15_sqmuxa_adt_net_109461_Ra1__net_1\, 
        \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Ra1_\, 
        CLEAR_STAT_12, NOEAD_C_I_0_13, NOEDTK_C_14, PULSEL4R_15, 
        PULSEL5R_16, \HWRES_3_ADT_NET_738__17\, \I1.BITCNTL0R_18\, 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__19\, 
        \I1.N_50_0_ADT_NET_1409__20\, 
        \I1.N_50_0_ADT_NET_1409__21\, 
        \I1.N_50_0_ADT_NET_1409__22\, \I1.N_598_23\, 
        \I1.N_324_24\, \I1.N_324_25\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__26\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__27\, 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, 
        \I2.N_4667_1_ADT_NET_1046__31\, 
        \I2.N_4667_1_ADT_NET_1046__32\, 
        \I2.N_4667_1_ADT_NET_1046__33\, 
        \I2.N_4667_1_ADT_NET_1046__34\, 
        \I2.N_4667_1_ADT_NET_1046__35\, 
        \I2.N_199_0_ADT_NET_1054__36\, 
        \I2.N_199_0_ADT_NET_1054__37\, \I2.CRC32_1_SQMUXA_0_38\, 
        \I2.WR_SRAM_2_ADT_NET_748__39\, \I2.N_4283_I_0_40\, 
        \I2.N_4283_I_0_41\, \I2.N_4283_I_0_42\, 
        \I2.N_4283_I_0_43\, \I2.N_4283_I_0_44\, 
        \I2.N_4283_I_0_45\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__46\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__47\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__48\, 
        \I2.REG_0L3R_ADT_NET_848__49\, \I3.REGMAPL57R_50\, 
        \I2.N_196_51\, \I2.N_196_52\, \I2.N_196_53\, 
        \I2.N_223_54\, \I2.N_4641_55\, \I2.N_4641_56\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__57\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__58\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__59\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_60\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_61\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_62\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_63\, 
        \I2.PIPE7_DTL27R_64\, \I2.PIPE7_DTL27R_65\, 
        \I2.PIPE7_DTL27R_66\, \I2.PIPE7_DTL27R_67\, 
        \I2.PIPE7_DTL27R_68\, \I2.PIPE7_DTL27R_69\, 
        \I2.PIPE7_DTL27R_70\, \I2.PIPE7_DTL27R_71\, 
        \I2.PIPE7_DTL27R_72\, \I2.PIPE7_DTL27R_73\, 
        \I2.PIPE7_DTL27R_74\, \I2.PIPE7_DTL27R_75\, 
        \I2.PIPE7_DTL27R_76\, \I2.PIPE7_DTL27R_77\, 
        \I2.PIPE7_DTL27R_78\, \I2.PIPE7_DTL27R_79\, 
        \I2.PIPE7_DTL27R_80\, \I2.PIPE7_DTL27R_81\, 
        \I2.PIPE7_DTL27R_82\, \I2.PIPE7_DTL27R_83\, 
        \I2.PIPE7_DTL27R_84\, \I2.PIPE7_DTL27R_85\, 
        \I2.PIPE7_DTL27R_86\, \I2.PIPE7_DTL27R_87\, 
        \I2.PIPE7_DTL27R_88\, \I2.PIPE7_DTL27R_89\, 
        \I2.PIPE7_DTL27R_90\, \I2.PIPE7_DTL27R_91\, \I1.N_65_92\, 
        \I1.N_41_9_ADT_NET_3739__93\, \I1.REG_16_SQMUXA_94\, 
        \I1.REG_16_SQMUXA_95\, \I1.N_253_96\, \I1.N_253_97\, 
        \I1.N_253_98\, \I1.REG_74_1_A0_0L228R_99\, 
        \I1.REG_74_1_A0_0L228R_100\, \I1.REG_74_1_A0_0L228R_101\, 
        \I1.REG_74_1_A0_0L228R_102\, \I2.N_74_103\, \I2.N_74_104\, 
        \I2.N_45_1_105\, \I2.N_45_1_106\, \I2.N_72_0_107\, 
        \I2.N_72_0_108\, \I2.N_89_0_109\, \I2.N_89_0_110\, 
        \I2.N_89_0_111\, \I3.REGMAPL39R_112\, 
        \I3.REGMAP_I_0_IL38R_113\, 
        \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, 
        \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, 
        \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, \I3.N_638_117\, 
        \I3.N_2017_118\, \I3.N_2017_119\, \I3.N_2015_120\, 
        \I3.N_2014_121\, \I3.N_2014_122\, \I3.UN1_REGMAP_34_123\, 
        \I3.UN1_REGMAP_34_124\, \I3.N_178_ADT_NET_1360__125\, 
        \I3.N_178_ADT_NET_1360__126\, 
        \I3.N_178_ADT_NET_1360__127\, \I3.N_354_0_128\, 
        \I3.N_354_0_129\, \I3.N_354_0_130\, \I2.N519_131\, 
        \I2.N_74_I_0_I_132\, \I2.N_128_133\, \I2.N_128_134\, 
        \I2.N_128_135\, \I2.RAMDT4L5R_136\, \I2.RAMDT4L5R_137\, 
        \I2.RAMDT4L5R_138\, \I2.RAMDT4L5R_139\, 
        \I2.RAMDT4L12R_140\, \I2.RAMDT4L12R_141\, 
        \I2.RAMDT4L12R_142\, \I2.RAMDT4L12R_143\, 
        \I2.RAMDT4L12R_144\, \I2.RAMDT4L12R_145\, 
        \I2.RAMDT4L12R_146\, \I3.N_264_0_ADT_NET_1653_RD1__147\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__148\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__149\, \I2.N_197_150\, 
        \I2.N_197_151\, \I2.N_197_152\, \I2.N_197_153\, 
        \I2.N_197_154\, \I2.N_182_ADT_NET_1007__155\, 
        \I2.N_223_156\, \I2.N_176_I_157\, 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__158\, 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_160\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__161\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__162\, 
        \I2.TOKOUTBS_163\, \I1.N_89_164\, \I1.N_89_165\, 
        \I1.N_12233_I_166\, \I1.N_243_167\, \I1.N_1169_168\, 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__169\, 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__170\, 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__171\, 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__172\, 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__173\, 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\, 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, 
        \I2.PIPE1_DT_2_SQMUXA_1_1_177\, \I2.N_3889_178\, 
        \I2.N_3889_179\, \I2.N_3879_180\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__181\, 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__182\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__183\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__184\, 
        \I2.N_4646_1_ADT_NET_19635__185\, 
        \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__186\, 
        \I1.REG_74_1L268R_187\, \I1.N_201_9_188\, 
        \I1.N_201_9_189\, \I1.N_396_190\, \I1.N_396_191\, 
        \I1.N_396_192\, 
        \I1.REG_74_4_I_A2_404_N_4_I_ADT_NET_1465__193\, 
        \I1.N_254_194\, \I1.N_254_195\, \I1.N_254_196\, 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__197\, 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__198\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__199\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__200\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__201\, 
        \I1.PAGECNT_326_202\, \I1.PAGECNT_327_203\, 
        \I1.N_473_204\, \I1.N_473_205\, \I1.N_473_206\, 
        \I1.UN1_SBYTE13_1_I_1_207\, \I1.UN1_SBYTE13_1_I_1_208\, 
        \I1.UN1_SBYTE13_1_I_1_209\, \I1.UN1_SBYTE13_1_I_1_210\, 
        \I1.N_328_I_0_211\, \I1.N_328_I_0_212\, 
        \I1.BYTECNTL2R_213\, \I1.BYTECNT_I_0_IL1R_214\, 
        \I2.MIC_REG2L3R_ADT_NET_834020_RD1__215\, 
        \I1.N_304_RA1__216\, \I1.N_65_ADT_NET_1433__217\, 
        \I1.N_65_ADT_NET_1433__218\, \I1.REG_29_SQMUXA_219\, 
        \I1.N_260_220\, \I1.N_260_221\, \I1.N_260_222\, 
        \I1.N_1383_223\, \I1.N_1383_224\, \I1.N_1383_225\, 
        \I1.N_223_226\, \I1.N_223_227\, \I1.N_590_228\, 
        \I1.N_590_229\, \I1.N_590_230\, \I1.N_590_231\, 
        \I1.N_321_232\, \I2.N_4038_233\, \I2.N_4283_I_0_234\, 
        \I2.N_4283_I_0_235\, 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__236\, 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_M3_237\, 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_M3_238\, NOESRAME_C_239, 
        NOESRAME_C_240, NOESRAME_C_241, NOESRAME_C_242, 
        NOESRAME_C_243, \I1.PAGECNTL9R_244\, \I1.PAGECNTL9R_245\, 
        \I1.PAGECNTL9R_246\, \I1.PAGECNTL6R_247\, 
        \I1.PAGECNTL6R_248\, \I1.PAGECNTL6R_249\, 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__251\, 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__252\, 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__253\, 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__254\, \I3.N_281_255\, 
        \I1.N_50_0_ADT_NET_109751__256\, 
        \I1.N_50_0_ADT_NET_109751__257\, 
        \I1.N_50_0_ADT_NET_109751__258\, \I3.N_268_259\, 
        \I1.BITCNTL1R_260\, \I3.N_2040_261\, \I3.N_1907_262\, 
        \I3.N_1907_263\, \I3.N_1907_264\, \I3.N_1907_265\, 
        \I3.N_1907_266\, \I1.N_49_267\, \I1.N_57_268\, 
        \I1.N_57_269\, \I1.N_113_ADT_NET_3714__270\, 
        \I1.N_113_ADT_NET_3714__271\, \I1.N_65_12_272\, 
        \I1.N_65_12_273\, \I1.N_273_9_274\, 
        \I1.REG_15_SQMUXA_275\, \I1.N_254_276\, \I1.N_254_277\, 
        \I1.N_1370_278\, \I1.REG_74_5_404_M1_E_0_279\, 
        \I1.REG_74_5_404_M1_E_0_280\, 
        \I1.N_50_0_ADT_NET_1409__281\, 
        \I1.N_50_0_ADT_NET_1409__282\, \I1.N_435_1_283\, 
        \I1.N_435_1_284\, \I1.N_435_1_285\, 
        \I2.DTE_CL_0_SQMUXA_2_0_286\, 
        \I2.DTE_CL_0_SQMUXA_2_0_287\, 
        \I2.DTE_CL_0_SQMUXA_2_0_288\, 
        \I2.DTE_CL_0_SQMUXA_2_0_289\, 
        \I2.DTE_CL_0_SQMUXA_2_0_290\, \I2.STATE2L4R_291\, 
        \I1.N_50_0_ADT_NET_1409__292\, 
        \I1.N_50_0_ADT_NET_1409__293\, 
        \I1.N_50_0_ADT_NET_1409__294\, 
        \I1.N_50_0_ADT_NET_1409__295\, \I1.N_232_1_296\, 
        \I2.UN1_NWPIPE7_2_297\, \I2.UN1_NWPIPE7_2_298\, 
        \I2.PIPE1_DT_2_SQMUXA_ADT_NET_803__299\, 
        \I2.NWPIPE1_4_SQMUXA_1_0_300\, 
        \I2.NWPIPE1_4_SQMUXA_1_0_301\, \I2.N_4261_302\, 
        \I2.N_4261_303\, \I2.N_4261_304\, \I2.NWPIPE5_305\, 
        \I2.G_EVNT_NUML1R_306\, \I1.SSTATEL0R_307\, 
        \I1.PAGECNTL5R_308\, \I1.PAGECNTL5R_309\, 
        \I1.PAGECNTL5R_310\, \I1.PAGECNTL5R_311\, 
        \I2.G_EVNT_NUM_I_0_IL0R_312\, \I1.N_238_RD1__313\, 
        \I1.N_238_RD1__314\, \I2.REG_0L3R_ADT_NET_19773_RD1__315\, 
        \I3.N_2044_316\, \I3.N_2017_317\, \I3.N_2016_318\, 
        \I3.N_2016_319\, \I1.N_50_0_ADT_NET_1409__320\, 
        \I1.N_50_0_ADT_NET_1409__321\, \I1.N_598_322\, 
        \I1.SSTATE_NS_IL5R_ADT_NET_107266__323\, 
        \I2.UN1_NWPIPE7_2_ADT_NET_73606__324\, 
        \I2.N_74_ADT_NET_55281__325\, 
        \I2.N_74_ADT_NET_55281__326\, 
        \I2.N_140_0_ADT_NET_947__327\, 
        \I2.N_140_0_ADT_NET_947__328\, 
        \I2.N_2826_1_ADT_NET_794__329\, 
        \I2.N_2826_1_ADT_NET_794__330\, 
        \I2.N_2826_1_ADT_NET_794__331\, 
        \I2.N_2826_1_ADT_NET_794__332\, \I2.G_EVNT_NUML2R_333\, 
        \I3.SINGCYC_334\, \I1.N_310_RD1__335\, 
        \I1.REG_74_1_380_M8_I_0_RD1__336\, 
        \I2.DWACT_FINC_E_0L0R_337\, \I2.N_2867_1_338\, 
        \I2.PIPE1_DT_42_3_0L28R_339\, 
        \I2.PIPE1_DT_42_3_0L28R_340\, 
        \I2.PIPE1_DT_42_3_0L28R_341\, 
        \I2.PIPE1_DT_42_3_0L28R_342\, \I2.N_3272_343\, 
        \I2.N_3272_344\, \I2.N_3272_345\, \I3.VAS_I_0_IL15R_346\, 
        \I3.VASL8R_347\, \I2.PIPE7_DTL26R_348\, 
        \I2.PIPE7_DTL26R_349\, \I2.PIPE7_DTL26R_350\, 
        \I2.PIPE7_DTL26R_351\, \I2.PIPE7_DTL26R_352\, 
        \I2.PIPE7_DTL26R_353\, \I2.PIPE7_DTL26R_354\, 
        \I2.PIPE7_DTL26R_355\, \I2.PIPE7_DTL26R_356\, 
        \I2.PIPE7_DTL26R_357\, \I2.PIPE7_DTL26R_358\, 
        \I2.PIPE7_DTL26R_359\, \I2.PIPE7_DTL26R_360\, 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__361\, 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__362\, 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__363\, \I3.N_549_364\, 
        \I3.N_549_365\, \I3.N_548_366\, \I3.N_548_367\, 
        \I3.N_548_368\, \I3.N_547_369\, \I3.N_547_370\, 
        \I3.N_547_371\, \I3.N_547_372\, \I3.N_546_373\, 
        \I3.N_546_374\, \I3.UN1_REGMAP_30_375\, 
        \I2.DT_SRAML0R_376\, \I2.N_4193_377\, \I3.STATE2L0R_378\, 
        \I2.N_2828_ADT_NET_1062__ADT_NET_835312_RD1__379\, 
        \I1.SSTATEL10R_380\, 
        \I2.MIC_REG1L3R_ADT_NET_834596_RD1__381\, 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__382\, 
        \I2.N525_383\, \I2.N_107_ADT_NET_256840__384\, 
        \I2.N_182_ADT_NET_1007__385\, 
        \I2.N_182_ADT_NET_1007__386\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854188__net_1\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854192__net_1\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854196__net_1\, 
        \I2.DT_SRAMl30r_adt_net_854200__net_1\, 
        \I2.REG_0l3r_adt_net_848__adt_net_854204__net_1\, 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, 
        \I2.REG_0l3r_adt_net_848__adt_net_854216__net_1\, 
        \I2.REG_0l3r_adt_net_848__adt_net_854220__net_1\, 
        \I2.REG_0l3r_adt_net_848__adt_net_854224__net_1\, 
        \I2.REG_0l3r_adt_net_848__adt_net_854228__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854232__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854236__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854240__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854244__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854248__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854260__net_1\, 
        \I2.N_2864_0_adt_net_854264__net_1\, 
        \I2.N_2864_0_adt_net_854268__net_1\, 
        \I2.N_2864_0_adt_net_854272__net_1\, 
        \I2.N_2864_0_adt_net_854276__net_1\, 
        \I3.REGMAPl17r_adt_net_854280__net_1\, 
        \I3.REGMAPl17r_adt_net_854284__net_1\, 
        \I3.REGMAPl17r_adt_net_854288__net_1\, 
        \I3.REGMAPl17r_adt_net_854292__net_1\, 
        \I3.REGMAPl17r_adt_net_854296__net_1\, 
        \I3.REGMAPl17r_adt_net_854300__net_1\, 
        \I3.REGMAPl9r_adt_net_854304__net_1\, 
        \I3.REGMAPl9r_adt_net_854308__net_1\, 
        \I3.REGMAPl9r_adt_net_854312__net_1\, 
        \I3.REGMAPl9r_adt_net_854316__net_1\, 
        \I3.REGMAPl9r_adt_net_854320__net_1\, 
        \I3.REGMAPl9r_adt_net_854324__net_1\, 
        \I3.REGMAPl9r_adt_net_854328__net_1\, 
        \I3.REGMAPl9r_adt_net_854332__net_1\, 
        \I3.N_1910_0_adt_net_854336__net_1\, 
        \I3.N_1910_0_adt_net_854340__net_1\, 
        \I3.N_1910_0_adt_net_854344__net_1\, 
        \I3.N_1910_0_adt_net_854348__net_1\, 
        \I3.N_1764_adt_net_854352__net_1\, 
        \I3.STATE1_ipl0r_adt_net_854356__net_1\, 
        \I3.STATE1_ipl0r_adt_net_854360__net_1\, 
        \I3.STATE1_ipl3r_adt_net_854364__net_1\, 
        \I3.STATE1_ipl3r_adt_net_854368__net_1\, 
        \I1.REG_30_sqmuxa_adt_net_854372__net_1\, 
        \I1.REG_30_sqmuxa_adt_net_854376__net_1\, 
        \I1.REG_15_sqmuxa_adt_net_1457__adt_net_854380__net_1\, 
        \I1.PAGECNT_322_adt_net_854384__net_1\, 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854396__net_1\, 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854400__net_1\, 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854404__net_1\, 
        \I2.N_128_adt_net_54291__adt_net_854408__net_1\, 
        \I2.PIPE4_DTl5r_adt_net_854412__net_1\, 
        \I2.PIPE4_DTl5r_adt_net_854416__net_1\, 
        \I2.PIPE4_DTl5r_adt_net_854420__net_1\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854424__net_1\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854428__net_1\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854432__net_1\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854436__net_1\, 
        \I2.N_4667_1_adt_net_1046__adt_net_854440__net_1\, 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854444__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854456__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854460__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854464__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854468__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854472__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854476__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854480__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854484__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854488__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854492__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854496__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854500__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854504__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854508__net_1\, 
        \I3.N_243_4_adt_net_1290__adt_net_854512__net_1\, 
        \I1.N_1367_i_adt_net_854516__net_1\, 
        \I1.un1_sbyte13_1_i_1_adt_net_854520__net_1\, 
        \I1.un1_sbyte13_1_i_1_adt_net_854524__net_1\, 
        \I1.un1_sbyte13_1_i_1_adt_net_106369__adt_net_854528__net_1\, 
        \PULSEl0r_adt_net_854532__net_1\, 
        \PULSEl0r_adt_net_854536__net_1\, 
        \I2.PIPE4_DTl3r_adt_net_854544__net_1\, 
        \I2.PIPE4_DTl3r_adt_net_854548__net_1\, 
        \I2.PIPE4_DTl8r_adt_net_854556__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854560__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854564__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854568__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854572__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854576__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854580__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854584__net_1\, 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854588__net_1\, 
        \I2.N_4671_adt_net_854592__net_1\, 
        \I2.N_4671_adt_net_854596__net_1\, 
        \I2.N_4671_adt_net_854600__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854612__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854616__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854624__net_1\, 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854628__net_1\, 
        \I2.N_3883_adt_net_854632__net_1\, 
        \I2.WOFFSETl0r_adt_net_854636__net_1\, 
        \I2.WOFFSETl0r_adt_net_854640__net_1\, 
        \I2.WOFFSETl0r_adt_net_854644__net_1\, 
        \I2.WOFFSETl0r_adt_net_854648__net_1\, EVREAD_387, 
        REGL32R_388, REGL33R_389, REGL117R_390, 
        \I2.STATE3L7R_391\, \I2.FIFO_END_EVNT_392\, 
        \I2.TEMPF_393\, \I2.BNC_IDL1R_394\, \I2.BNC_IDL0R_395\, 
        \I2.EVNT_NUML0R_396\, \I2.EVNT_NUML1R_397\, 
        \I2.FCNT_C0_398\, \I2.G_EVNT_NUML3R_399\, 
        \I2.ROFFSETL2R_400\, \I2.ENDF_401\, \I2.ENDF_402\, 
        \I2.END_EVNT2_403\, \I2.END_EVNT2_404\, 
        \I2.END_EVNT5_405\, \I2.END_EVNT5_406\, 
        \I2.END_EVNT10_407\, \I2.PIPE4_DTL11R_408\, 
        \I2.PIPE4_DTL11R_409\, \I2.PIPE4_DTL11R_410\, 
        \I2.PIPE4_DTL0R_411\, \I2.STATE3L2R_412\, 
        \I2.STATE3L2R_413\, \I2.STATE3L2R_414\, 
        \I2.STATE3L3R_415\, \I2.STATE3L3R_416\, 
        \I1.SSTATEL6R_417\, \I1.SSTATEL4R_418\, 
        \I3.STATE1_IPL9R_419\, \I3.STATE1_IPL8R_420\, 
        \I3.REGMAPL0R_421\, \I3.MBLTCYC_422\, \I3.MBLTCYC_423\, 
        \I3.WRITES_424\, \I3.DSS_425\, \I3.STATE1_IPL8R_426\, 
        \I3.STATE1_IPL9R_427\, \I3.TCNTL0R_428\, \I3.TCNTL1R_429\, 
        \I3.TCNTL2R_430\, \I3.REG3L4R_431\, \I3.REG3L4R_432\, 
        \I1.SSTATEL9R_433\, \I1.BYTECNTL3R_434\, 
        \I1.BYTECNT_I_0_IL1R_435\, \I1.BYTECNTL0R_436\, 
        \I2.STATE2L3R_437\, \I2.STATE2L3R_438\, 
        \I2.STATE2L3R_439\, \I2.STATE2L3R_440\, 
        \I2.RAMDT4L11R_441\, \I2.RAMDT4L10R_442\, 
        \I2.RAMDT4L7R_443\, \I3.REGMAPL16R_444\, 
        \I3.REGMAPL43R_445\, \I3.REGMAPL34R_446\, 
        \I3.REGMAP_I_IL46R_447\, \I3.REGMAPL47R_448\, 
        \I3.REGMAPL37R_449\, \I3.REGMAP_I_0_IL40R_450\, 
        \I3.REGMAPL44R_451\, \I3.REGMAP_I_0_IL45R_452\, 
        \I2.MIC_REG2L3R_ADT_NET_834020_RD1__453\, 
        \I2.MIC_REG3L1R_454\, \I2.MIC_REG1L1R_455\, 
        \I1.PAGECNTL8R_456\, \I1.PAGECNTL8R_457\, 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_1_RD1__458\, 
        \I3.REGMAPL7R_459\, \I3.REGMAPL7R_460\, 
        \I3.REGMAPL33R_461\, \I2.MIC_REG3L2R_462\, 
        \I2.MIC_REG2L2R_463\, \I2.MIC_REG1L2R_464\, 
        \I2.TRGSERVL0R_465\, \I2.TRGSERVL0R_466\, 
        \I2.TRGSERVL0R_467\, \I2.TRGSERVL1R_468\, 
        \I2.TRGSERVL1R_469\, \I2.TRGSERVL1R_470\, 
        \I2.PIPE4_DTL9R_471\, \I2.PIPE4_DTL9R_472\, 
        \I2.PIPE4_DT_I_IL1R_473\, \I2.PIPE4_DT_I_IL1R_474\, 
        \I2.PIPE4_DTL10R_475\, \I2.PIPE4_DTL10R_476\, 
        \I2.PIPE4_DTL4R_477\, \I2.PIPE4_DTL4R_478\, 
        \I2.PIPE4_DTL6R_479\, \I2.PIPE4_DTL6R_480\, 
        \I2.PIPE4_DTL7R_481\, \I2.PIPE4_DTL7R_482\, 
        \I2.PIPE4_DTL8R_483\, \I2.MIC_REG3L3R_484\, 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_N_8_RD1__485\, 
        \I1.N_349_RD1__486\, \I1.N_341_RD1__487\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__488\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__489\, 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__490\, 
        \I2.MIC_REG2L3R_ADT_NET_834020_RD1__491\, 
        \I1.PAGECNTL9R_492\, \I1.PAGECNT_325_493\, \I1.N_656_494\, 
        \I1.N_656_495\, \I1.N_656_496\, \I1.N_328_I_0_497\, 
        \I1.N_328_I_0_498\, \I1.N_325_499\, \I1.N_325_500\, 
        \I1.N_325_501\, \I2.PIPE7_DTL31R_502\, 
        \I2.TDCDBSL31R_503\, \I2.FCNTL1R_504\, 
        \I2.ROFFSETL0R_505\, \I2.ROFFSETL1R_506\, 
        \I2.STATE2L5R_507\, \I2.STATE2L5R_508\, \I2.TOKOUTAS_509\, 
        \I2.PIPE4_DTL12R_510\, \I2.PIPE4_DTL12R_511\, 
        \I2.PIPE4_DTL12R_512\, \I2.PIPE4_DTL2R_513\, 
        \I2.PIPE4_DTL2R_514\, \I2.RPAGEL15R_515\, 
        \I2.RPAGEL15R_516\, \I2.RPAGEL15R_517\, 
        \I2.RPAGEL15R_518\, \I2.RPAGEL15R_519\, 
        \I2.RPAGEL15R_520\, \I2.RPAGEL15R_521\, 
        \I2.RPAGEL15R_522\, \I2.N_4646_1_ADT_NET_19637_RD1__523\, 
        \I1.SSTATEL8R_524\, \I1.PAGECNTL7R_525\, 
        \I1.PAGECNTL7R_526\, \I2.RAMDT4L8R_527\, 
        \I3.REGMAPL35R_528\, \I3.REGMAP_I_0_IL36R_529\, 
        \I3.REGMAPL41R_530\, \I3.REGMAP_I_0_IL42R_531\, 
        \I3.REGMAPL26R_532\, \I3.REGMAPL27R_533\, 
        \I3.REGMAP_I_0_IL19R_534\, \I3.REGMAPL28R_535\, 
        \I2.MIC_REG2L1R_536\, \I3.REGMAP_I_0_IL58R_537\, 
        \I1.REG_74_1_380_M8_I_0_RD1__538\, \I3.REGMAPL57R_539\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__540\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__541\, \I2.N346_0_542\, 
        \I2.N303_0_543\, \I2.N270_0_544\, \I2.N270_0_545\, 
        \I2.N273_546\, \I2.N273_547\, \I2.N_218_548\, 
        \I2.N_207_549\, \I2.N_207_550\, \I2.N_198_551\, 
        \I2.N_4672_552\, \I2.N_4672_553\, \I2.N_189_554\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854652__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854656__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854660__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854664__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854668__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854672__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854676__net_1\, 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854680__net_1\, 
        \I3.N_2034_adt_net_854684__net_1\, 
        \I3.N_57_i_0_0_adt_net_854688__net_1\, 
        \I3.N_57_i_0_0_adt_net_854692__net_1\, 
        \I3.N_57_i_0_0_adt_net_854696__net_1\, 
        \I3.N_57_i_0_0_adt_net_854700__net_1\, 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, 
        \I1.N_97_6_adt_net_854712__net_1\, 
        \I1.REG_10_sqmuxa_adt_net_854716__net_1\, 
        \I1.REG_10_sqmuxa_adt_net_854720__net_1\, 
        \I1.REG_9_sqmuxa_adt_net_854724__net_1\, 
        \I1.REG_9_sqmuxa_adt_net_854728__net_1\, 
        \I3.PULSE_330_adt_net_854732__net_1\, 
        \I3.PULSE_330_adt_net_854736__net_1\, 
        \I3.N_1409_adt_net_854740__net_1\, 
        \I3.N_1409_adt_net_854744__net_1\, 
        \I3.N_311_adt_net_854748__net_1\, 
        \I3.N_311_adt_net_854752__net_1\, 
        \I1.N_592_adt_net_854756__net_1\, 
        \I1.N_137_adt_net_854760__net_1\, 
        \I1.N_137_adt_net_854764__net_1\, 
        \I1.N_145_adt_net_854768__net_1\, 
        \I1.N_145_adt_net_854772__net_1\, 
        \I1.REG_24_sqmuxa_adt_net_854776__net_1\, 
        \I1.REG_24_sqmuxa_adt_net_854780__net_1\, 
        \I1.N_41_9_adt_net_854784__net_1\, 
        \I1.N_347_adt_net_854788__net_1\, 
        \I1.N_347_adt_net_854792__net_1\, 
        \I1.N_273_6_i_0_adt_net_854796__net_1\, 
        \I1.N_268_Rd1__adt_net_854800__net_1\, 
        \I1.N_237_adt_net_854804__net_1\, 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, 
        \I1.N_1169_adt_net_854812__net_1\, 
        \I1.PAGECNTl9r_adt_net_854816__net_1\, 
        \I1.N_1169_adt_net_854820__net_1\, 
        \I1.N_1169_adt_net_854824__net_1\, 
        \I1.N_1169_adt_net_854828__net_1\, 
        \I1.REG_74_1_a0_0l228r_adt_net_854832__net_1\, 
        \I1.REG_74_1_396_m7_i_3_adt_net_854840__net_1\, 
        \I1.N_223_adt_net_854844__net_1\, 
        \I1.N_223_adt_net_854848__net_1\, 
        \I1.PAGECNT_318_adt_net_854852__net_1\, 
        \I1.PAGECNT_318_adt_net_854856__net_1\, 
        \I1.PAGECNT_319_adt_net_854860__net_1\, 
        \I1.PAGECNT_319_adt_net_854864__net_1\, 
        \I1.PAGECNT_320_adt_net_854868__net_1\, 
        \I1.PAGECNT_320_adt_net_854872__net_1\, 
        \I1.PAGECNT_320_adt_net_854876__net_1\, 
        \I1.PAGECNT_321_adt_net_854880__net_1\, 
        \I1.N_238_Rd1__adt_net_854884__net_1\, 
        \I1.N_238_Rd1__adt_net_854888__net_1\, 
        \I1.PAGECNTe_adt_net_854892__net_1\, 
        \I1.PAGECNTe_adt_net_854896__net_1\, 
        \I1.PAGECNTe_adt_net_854900__net_1\, 
        \I1.N_370_adt_net_854904__net_1\, 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854908__net_1\, 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854912__net_1\, 
        \I1.N_311_i_i_Rd1__adt_net_854920__net_1\, 
        \I1.PAGECNTl6r_adt_net_854924__net_1\, 
        \I1.PAGECNTl6r_adt_net_854928__net_1\, 
        \I1.PAGECNTl6r_adt_net_854932__net_1\, 
        \I2.N258_0_adt_net_854936__net_1\, 
        \I2.LSRAM_OUTl13r_adt_net_854940__net_1\, 
        \I2.LSRAM_OUTl14r_adt_net_854944__net_1\, 
        \I2.PIPE4_DTl7r_adt_net_854552__adt_net_854948__net_1\, 
        \I2.N_2358_tz_tz_adt_net_854952__net_1\, 
        \I2.N_2358_tz_tz_adt_net_854956__net_1\, 
        \I2.N_2867_1_adt_net_854960__net_1\, 
        \I2.N_2867_1_adt_net_854964__net_1\, 
        \I2.N_4283_i_0_adt_net_854968__net_1\, 
        \I2.N_4283_i_0_adt_net_854972__net_1\, 
        \I3.N_203_adt_net_854976__net_1\, 
        \I2.WOFFSETl4r_adt_net_854980__net_1\, 
        \I2.WOFFSETl2r_adt_net_854984__net_1\, 
        \I2.WOFFSETl3r_adt_net_854988__net_1\, 
        \I2.WOFFSETl1r_adt_net_854992__net_1\, 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996__net_1\, 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855000__net_1\, 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        \I3.un1_REGMAP_30_adt_net_855008__net_1\, 
        \I3.REGMAPl23r_adt_net_855012__net_1\, 
        \I3.REGMAPl23r_adt_net_855016__net_1\, 
        \I1.BYTECNTl2r_adt_net_855020__net_1\, 
        \I2.PIPE4_DTl8r_adt_net_854556__adt_net_855024__net_1\, 
        \I2.N_64_0_adt_net_855028__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855032__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855036__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044__net_1\, 
        \I2.N_201_adt_net_855048__net_1\, 
        \I2.N_4669_adt_net_855052__net_1\, 
        \I2.WPAGEe_adt_net_855056__net_1\, 
        \I2.WPAGEe_adt_net_855060__net_1\, 
        \I2.N_3283_adt_net_855064__net_1\, 
        \I2.N_3887_adt_net_855068__net_1\, 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855076__net_1\, 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855088__net_1\, 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092__net_1\, 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096__net_1\, 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100__net_1\, 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855104__net_1\, 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, 
        \I2.STATE2l1r_adt_net_855116__net_1\, 
        \I2.STATE2l1r_adt_net_855120__net_1\, 
        \I2.STATE2l1r_adt_net_855124__net_1\, 
        \I2.STATE2l1r_adt_net_855128__net_1\, 
        \I2.STATE2l1r_adt_net_855132__net_1\, 
        \I2.SUB8_1_sqmuxa_0_adt_net_855136__net_1\, 
        \I2.SUB8_1_sqmuxa_0_adt_net_855140__net_1\, 
        \I2.SUB8_1_sqmuxa_0_adt_net_855144__net_1\, 
        \I2.SUB8_1_sqmuxa_0_adt_net_855148__net_1\, 
        \I2.SUB8_1_sqmuxa_0_adt_net_855152__net_1\, 
        \I2.SUB8_1_sqmuxa_0_adt_net_855156__net_1\, 
        \I2.SUB8_1_sqmuxa_0_adt_net_855160__net_1\, 
        \I2.N_587_adt_net_1201__adt_net_855164__net_1\, 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\, 
        \I2.PIPE7_DTl30r_adt_net_855172__net_1\, 
        \I2.STATE1l12r_adt_net_855176__net_1\, 
        \I2.STATE1l12r_adt_net_855180__net_1\, 
        \I2.STATE1l12r_adt_net_855184__net_1\, 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855192__net_1\, 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855196__net_1\, 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855200__net_1\, 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855208__net_1\, 
        \I2.STATE2l2r_adt_net_855212__net_1\, 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855220__net_1\, 
        \I2.N_3279_0_adt_net_855224__net_1\, 
        \I2.N_3279_0_adt_net_855228__net_1\, 
        \I2.N_3279_0_adt_net_855232__net_1\, 
        \I2.N_3279_0_adt_net_855236__net_1\, 
        \I2.CHAINB_EN244_c_0_adt_net_855240__net_1\, 
        \I2.CHAINB_EN244_c_0_adt_net_855244__net_1\, 
        \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\, 
        \I2.N_3876_adt_net_855252__net_1\, 
        \I2.N_3876_adt_net_855256__net_1\, 
        \I2.CHAINA_EN244_i_adt_net_855260__net_1\, 
        \I2.CHAINA_EN244_i_adt_net_855264__net_1\, 
        \I2.N_3877_adt_net_855268__net_1\, TICKL0R_555, 
        TICKL0R_556, TICKL0R_557, TICKL0R_558, END_FLUSH_559, 
        END_FLUSH_560, COM_SERS_561, EVREAD_562, REGL34R_563, 
        REGL35R_564, REGL36R_565, REGL37R_566, EV_RES_C_567, 
        EV_RES_C_568, EV_RES_C_569, TDCTRG_C_570, 
        \I5.SSTATE1L13R_571\, \I5.PULSE_FL_572\, 
        \I5.BITCNT_C0_573\, \I2.STATE1L17R_574\, \I2.NWPIPE4_575\, 
        \I2.NWPIPE4_576\, \I2.NWPIPE5_577\, \I2.NWPIPE2_578\, 
        \I2.FIFO_END_EVNT_579\, \I2.TDCGDB1_580\, 
        \I2.TRGSERVL2R_581\, \I2.TRGSERVL2R_582\, 
        \I2.TRGSERVL2R_583\, \I2.TRGSERVL2R_584\, 
        \I2.BNC_IDL3R_585\, \I2.OFFSETL0R_586\, 
        \I2.STATE2L0R_587\, \I2.STATE2L0R_588\, 
        \I2.STATE2L2R_589\, \I2.STATE1L10R_590\, 
        \I2.STATE1L5R_591\, \I2.FIFO_FULL_592\, 
        \I2.SRAM_FULL_593\, \I2.END_CHAINB1_594\, 
        \I2.STOP_RDSRAM_595\, \I2.EVNT_NUML2R_596\, 
        \I2.EVNT_NUML3R_597\, \I2.EVNT_NUML4R_598\, 
        \I2.FCNTL2R_599\, \I2.FCNTL2R_600\, \I2.STATE1L13R_601\, 
        \I2.L2ARRL0R_602\, \I2.L2ARRL1R_603\, \I2.L2ARRL2R_604\, 
        \I2.L2ARRL3R_605\, \I2.G_EVNT_NUML4R_606\, 
        \I2.RPAGEL12R_607\, \I2.RPAGEL12R_608\, 
        \I2.RPAGEL13R_609\, \I2.RPAGEL13R_610\, 
        \I2.RPAGEL13R_611\, \I2.RPAGEL14R_612\, 
        \I2.RPAGEL14R_613\, \I2.RPAGEL14R_614\, 
        \I2.RPAGEL14R_615\, \I2.RPAGEL14R_616\, 
        \I2.ROFFSETL3R_617\, \I2.ENDF_618\, \I2.END_EVNT2_619\, 
        \I2.PIPE5_DTL31R_620\, \I2.PIPE5_DTL30R_621\, 
        \I2.PIPE5_DTL30R_622\, \I2.PIPE5_DTL23R_623\, 
        \I2.PIPE5_DTL23R_624\, \I2.PIPE5_DTL21R_625\, 
        \I2.PIPE5_DTL21R_626\, \I2.STATE1L18R_627\, 
        \I2.STATE1L18R_628\, \I2.TOKOUTBS_629\, 
        \I2.STATE1L6R_630\, \I2.STATE1L9R_631\, 
        \I2.STATE1L7R_632\, \I2.STATE1L7R_633\, 
        \I2.PIPE4_DTL19R_634\, \I2.PIPE4_DTL17R_635\, 
        \I2.PIPE4_DTL17R_636\, \I2.PIPE4_DTL15R_637\, 
        \I2.PIPE4_DTL14R_638\, \I2.PIPE4_DTL14R_639\, 
        \I2.PIPE4_DTL14R_640\, \I2.PIPE4_DTL13R_641\, 
        \I2.PIPE4_DTL13R_642\, \I2.PIPE4_DTL0R_643\, 
        \I2.TOKOUT_FL_644\, \I2.STATE1L12R_645\, 
        \I2.STATE1L12R_646\, \I2.STATE1L12R_647\, 
        \I2.STATE1L8R_648\, \I2.L2TYPEL0R_649\, 
        \I2.L2TYPEL8R_650\, \I2.L2TYPEL4R_651\, 
        \I2.L2TYPEL12R_652\, \I2.L2TYPEL2R_653\, 
        \I2.L2TYPEL10R_654\, \I2.L2TYPEL6R_655\, 
        \I2.L2TYPEL14R_656\, \I2.L2TYPE_I_0_IL1R_657\, 
        \I2.L2TYPE_I_0_IL9R_658\, \I2.L2TYPE_I_0_IL5R_659\, 
        \I2.L2TYPE_I_0_IL13R_660\, \I2.L2TYPEL3R_661\, 
        \I2.L2TYPEL11R_662\, \I2.L2TYPEL7R_663\, 
        \I2.L2TYPEL15R_664\, \I2.PIPE5_DTL22R_665\, 
        \I2.PIPE5_DTL22R_666\, \I2.PIPE9_DTL31R_667\, 
        \I2.PIPE9_DTL30R_668\, \I2.PIPE9_DTL29R_669\, 
        \I2.OFFSETL7R_670\, \I2.OFFSETL7R_671\, 
        \I2.OFFSETL6R_672\, \I2.OFFSETL6R_673\, 
        \I2.OFFSETL5R_674\, \I2.OFFSETL4R_675\, 
        \I2.OFFSETL4R_676\, \I2.OFFSETL3R_677\, 
        \I2.OFFSETL2R_678\, \I2.OFFSETL1R_679\, 
        \I2.OFFSETL1R_680\, \I2.PIPE7_DTL25R_681\, 
        \I2.PIPE7_DTL25R_682\, \I2.PIPE7_DTL25R_683\, 
        \I2.PIPE7_DTL25R_684\, \I2.PIPE7_DTL25R_685\, 
        \I2.PIPE7_DTL25R_686\, \I2.PIPE7_DTL25R_687\, 
        \I2.NWPIPE7_688\, \I2.NWPIPE7_689\, \I2.PIPE7_DTL15R_690\, 
        \I2.PIPE7_DTL14R_691\, \I2.PIPE7_DTL13R_692\, 
        \I2.PIPE7_DTL12R_693\, \I2.PIPE7_DTL11R_694\, 
        \I2.PIPE7_DTL10R_695\, \I2.PIPE7_DTL9R_696\, 
        \I2.PIPE7_DTL8R_697\, \I2.PIPE7_DTL7R_698\, 
        \I2.PIPE7_DTL6R_699\, \I2.PIPE7_DTL5R_700\, 
        \I2.PIPE7_DTL3R_701\, \I2.PIPE7_DTL2R_702\, 
        \I2.PIPE7_DTL1R_703\, \I2.SUB8L7R_704\, \I2.SUB8L7R_705\, 
        \I2.SUB8L6R_706\, \I2.SUB8L5R_707\, \I2.SUB8L4R_708\, 
        \I2.SUB8L4R_709\, \I2.SUB8L3R_710\, \I2.BNC_IDL2R_711\, 
        \I2.BNC_IDL4R_712\, \I1.SSTATEL3R_713\, 
        \I1.SSTATEL6R_714\, \I1.SSTATEL4R_715\, \I1.COMMAND_716\, 
        \I3.STATE1_IPL9R_717\, \I3.DSS_718\, \I3.REGMAPL10R_719\, 
        \I3.STATE2L0R_720\, \I3.STATE2L2R_721\, 
        \I3.REGMAPL0R_722\, \I3.REGMAPL51R_723\, 
        \I3.REGMAPL1R_724\, \I3.REGMAPL1R_725\, 
        \I3.REGMAPL13R_726\, \I3.ADACKCYC_727\, 
        \I3.STATE1L10R_728\, \I3.EVREAD_DS_729\, 
        \I3.STATE1_IPL6R_730\, \I3.STATE1_IPL9R_731\, 
        \I3.REGMAPL14R_732\, \I3.REGMAPL14R_733\, 
        \I3.REGMAPL14R_734\, \I3.REGMAPL14R_735\, 
        \I3.REGMAPL2R_736\, \I3.REGMAPL2R_737\, 
        \I3.REGMAPL3R_738\, \I3.REGMAPL8R_739\, 
        \I3.REGMAPL8R_740\, \I3.REGMAPL8R_741\, \I3.REG3L2R_742\, 
        \I3.REGMAPL11R_743\, \I3.REG3L1R_744\, \I3.REG3L0R_745\, 
        \I3.REGMAPL12R_746\, \I3.VAS_I_0_IL7R_747\, 
        \I3.VASL6R_748\, \I2.WPAGEL15R_749\, \I2.WPAGEL14R_750\, 
        \I2.WPAGEL13R_751\, \I2.WPAGEL12R_752\, 
        \I1.BITCNTL2R_753\, \I1.SSTATEL7R_754\, 
        \I1.SSTATEL0R_755\, PULSEL0R_756, 
        \I2.N_2828_ADT_NET_1062__ADT_NET_835308_RD1__757\, 
        \I1.SSTATEL2R_758\, \I1.SSTATEL10R_759\, \I1.LUT_760\, 
        \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__761\, 
        \I1.N_311_I_I_RD1__762\, \I2.STATE5L2R_763\, 
        \I2.RAMDT4L4R_764\, \I2.RAMDT4L3R_765\, 
        \I2.RAMDT4L10R_766\, \I2.RAMDT4L2R_767\, 
        \I2.RAMDT4L9R_768\, \I2.RAMDT4L1R_769\, 
        \I2.RAMDT4L0R_770\, \I3.REGMAPL29R_771\, 
        \I3.REGMAP_I_0_IL30R_772\, \I3.REGMAPL31R_773\, 
        \I3.REGMAP_I_0_IL32R_774\, \I3.REGMAPL22R_775\, 
        \I3.REGMAPL25R_776\, \I3.REGMAP_I_0_IL24R_777\, 
        \I3.REGMAPL18R_778\, \I3.REGMAPL21R_779\, 
        \I3.REGMAPL20R_780\, \I3.REGMAPL55R_781\, 
        \I3.REGMAPL55R_782\, \I3.REGMAPL9R_783\, 
        \I3.REGMAPL9R_784\, \I3.REGMAPL9R_785\, 
        \I3.REGMAPL9R_786\, \I3.LWORDS_787\, \I3.LWORDS_788\, 
        \I2.MIC_REG3L2R_789\, \I2.PIPE4_DTL9R_790\, 
        \I2.PIPE4_DTL10R_791\, \I2.PIPE4_DTL10R_792\, 
        \I2.RAMDT4L12R_793\, \I2.RAMDT4L12R_794\, 
        \I2.RAMDT4L12R_795\, \I2.RAMDT4L12R_796\, 
        \I2.RAMDT4L12R_797\, \I2.RAMDT4L12R_798\, 
        \I2.RAMDT4L12R_799\, \I2.RAMDT4L12R_800\, 
        \I2.RAMDT4L12R_801\, \I3.REGMAP_I_0_IL58R_802\, 
        \I3.REGMAP_I_0_IL58R_803\, \I2.MIC_REG3L3R_804\, 
        \I1.BITCNTL0R_805\, \I2.N_4646_1_ADT_NET_1645_RD1__806\, 
        \I3.REGMAPL57R_807\, \I3.REGMAPL57R_808\, 
        \I2.RAMDT4L5R_809\, \I2.RAMDT4L5R_810\, 
        \I2.RAMDT4L5R_811\, \I2.RAMDT4L5R_812\, 
        \I2.RAMDT4L5R_813\, \I2.RAMDT4L5R_814\, 
        \I2.RAMDT4L5R_815\, \I2.RAMDT4L5R_816\, 
        \I2.RAMDT4L5R_817\, \I2.RAMDT4L5R_818\, 
        \I2.RAMDT4L5R_819\, \I2.RAMDT4L5R_820\, 
        \I2.RAMDT4L5R_821\, \I2.RAMDT4L12R_822\, 
        \I2.RAMDT4L12R_823\, \I2.RAMDT4L12R_824\, 
        \I2.RAMDT4L12R_825\, \I2.RAMDT4L12R_826\, 
        \I2.RAMDT4L12R_827\, \I2.RAMDT4L12R_828\, 
        \I2.RAMDT4L12R_829\, \PULSE_0L0R_ADT_NET_834380_RD1__830\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__831\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__832\, NOESRAME_C_833, 
        NOESRAME_C_834, \I1.PAGECNTL9R_835\, \I1.PAGECNTL6R_836\, 
        \I2.ENDF_837\, \I2.ENDF_838\, \I2.END_EVNT5_839\, 
        \I2.END_EVNT5_840\, \I2.PIPE4_DTL11R_841\, 
        \I2.PIPE4_DTL11R_842\, \I2.PIPE4_DTL11R_843\, 
        \I3.MBLTCYC_844\, \I2.PIPE4_DTL9R_845\, 
        \I2.PIPE4_DTL9R_846\, \I2.PIPE4_DTL9R_847\, 
        \I2.PIPE4_DT_I_IL1R_848\, \I2.PIPE4_DT_I_IL1R_849\, 
        \I2.PIPE4_DTL10R_850\, \I2.PIPE4_DTL10R_851\, 
        \I2.PIPE4_DTL4R_852\, \I2.PIPE4_DTL6R_853\, 
        \I2.PIPE4_DTL6R_854\, \I2.PIPE4_DTL12R_855\, 
        \I2.PIPE4_DTL12R_856\, \I2.PIPE4_DTL12R_857\, 
        \I2.PIPE4_DTL12R_858\, \I2.PIPE4_DTL2R_859\, 
        \I2.PIPE4_DTL2R_860\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__861\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__862\, 
        \PULSE_0L0R_ADT_NET_834380_RD1__863\, \I2.N350_864\, 
        \I2.N307_2_865\, \I2.N264_0_866\, \I2.N264_0_867\, 
        \I2.N267_0_868\, \I2.N267_0_869\, 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__870\, 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__871\, 
        REGL34R_872, REGL38R_873, \I2.ROFFSETL4R_874\, 
        \I2.STATE1L18R_875\, \I3.REGMAPL0R_876\, 
        \I3.STATE1_IPL9R_877\, \I3.TCNTL3R_878\, \I3.END_PK_879\, 
        \I3.SINGCYC_880\, \I3.SINGCYC_881\, \I1.SSTATEL10R_882\, 
        \I2.RAMDT4L4R_883\, 
        \I1.PAGECNT_0L9R_ADT_NET_835132_RD1__884\, 
        \I3.STATE1_IPL2R_885\, \I3.STATE1_IPL2R_886\, 
        \I2.REG_0L3R_ADT_NET_19771_RD1__887\, 
        \I2.REG_0L3R_ADT_NET_19773_RD1__888\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__889\, 
        \I2.N_4646_1_ADT_NET_1645_RD1__890\, \I2.END_EVNT10_891\, 
        \I2.FCNTL2R_892\, \I2.PIPE5_DTL21R_893\, 
        \I2.PIPE5_DTL21R_894\, 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\, 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\, 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855280__net_1\, 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\, 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\, 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\, 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, 
        \I3.N_127_adt_net_855312__net_1\, 
        \I3.N_1935_adt_net_855316__net_1\, 
        \I3.N_1935_adt_net_855320__net_1\, 
        \I3.N_1935_adt_net_855324__net_1\, 
        \I3.N_1935_adt_net_855328__net_1\, 
        \I3.N_1935_adt_net_855332__net_1\, 
        \I3.N_1917_adt_net_855336__net_1\, 
        \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, 
        \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344__net_1\, 
        \I3.N_1463_i_1_adt_net_855348__net_1\, 
        \I3.N_1463_i_1_adt_net_855352__net_1\, 
        \I3.N_1463_i_1_adt_net_855356__net_1\, 
        \I3.N_1463_i_1_adt_net_855360__net_1\, 
        \I3.N_1463_i_1_adt_net_855364__net_1\, 
        \I3.N_354_0_adt_net_855368__net_1\, 
        \I3.N_354_0_adt_net_855372__net_1\, 
        \I3.N_1905_1_adt_net_855376__net_1\, 
        \I3.N_1905_1_adt_net_855380__net_1\, 
        \I3.N_1905_1_adt_net_855384__net_1\, 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\, 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\, 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__adt_net_855516__net_1\, 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536__net_1\, 
        \I1.N_321_adt_net_855540__net_1\, 
        \PULSEl0r_adt_net_854532__adt_net_855544__net_1\, 
        \I1.PAGECNTl5r_adt_net_855548__net_1\, 
        \REG_i_il5r_adt_net_855552__net_1\, 
        \REG_i_il5r_adt_net_855556__net_1\, 
        \REG_i_il5r_adt_net_855560__net_1\, 
        \I2.SUB8l13r_adt_net_855564__net_1\, 
        \I2.SUB8l14r_adt_net_855568__net_1\, 
        \I2.SUB8l15r_adt_net_855572__net_1\, 
        \I2.SUB8l12r_adt_net_855576__net_1\, 
        \I2.SUB8l11r_adt_net_855580__net_1\, 
        \I2.N_3558_i_adt_net_855584__net_1\, 
        \I2.N_3822_adt_net_855588__net_1\, 
        \I2.N_22_i_0_adt_net_855592__net_1\, 
        \I2.N_22_i_0_adt_net_855596__net_1\, 
        \I2.PIPE4_DTl5r_adt_net_854412__adt_net_855600__net_1\, 
        \I2.N_3_0_adt_net_1070__adt_net_855604__net_1\, 
        \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\, 
        \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\, 
        \I2.N_4547_1_adt_net_1209__adt_net_855616__net_1\, 
        \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, 
        \I3.REG3_0_sqmuxa_adt_net_855624__net_1\, 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, 
        \I3.N_1906_i_0_0_adt_net_855636__net_1\, 
        \I3.N_1906_i_0_0_adt_net_855640__net_1\, 
        \I2.MIC_REG2_312_adt_net_855644__net_1\, 
        \I2.N_3234_adt_net_855648__net_1\, 
        \I2.N_3234_adt_net_855652__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668__net_1\, 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672__net_1\, 
        \I2.STATE2l4r_adt_net_855676__net_1\, 
        \I2.STATE2l4r_adt_net_855680__net_1\, 
        \I2.STATE2l4r_adt_net_855684__net_1\, 
        \I2.STATE2l4r_adt_net_855688__net_1\, 
        \I2.STATE2l4r_adt_net_855692__net_1\, 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\, 
        \I2.N_1170_adt_net_1217__adt_net_855700__net_1\, 
        \I2.N_1170_adt_net_1217__adt_net_855704__net_1\, 
        \I2.N_176_i_adt_net_855708__net_1\, 
        \I2.WOFFSETl0r_adt_net_854636__adt_net_855712__net_1\, 
        \I2.L2AS_adt_net_855716__net_1\, 
        \I2.L2AS_adt_net_855720__net_1\, 
        \I2.L2AS_adt_net_855724__net_1\, 
        \I2.N_565_0_adt_net_855728__net_1\, 
        \I2.N_565_0_adt_net_855732__net_1\, 
        \I2.N_565_0_adt_net_855736__net_1\, 
        \I2.TEMPF_adt_net_855740__net_1\, 
        \I2.TEMPF_adt_net_855744__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855756__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768__net_1\, 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, 
        \I2.un8_evread_1_adt_net_855780__net_1\, 
        \I2.un8_evread_1_adt_net_855784__net_1\, 
        \I2.un8_evread_1_adt_net_855788__net_1\, 
        \I2.un8_evread_1_adt_net_855792__net_1\, 
        \I2.un8_evread_1_adt_net_855796__net_1\, 
        \I2.dataout_0_adt_net_855800__net_1\, 
        \I2.dataout_0_adt_net_855804__net_1\, 
        \I2.dataout_0_adt_net_855808__net_1\, 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, 
        \I2.STATE1_ns_0l5r_adt_net_855816__net_1\, 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\, 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\, 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\, 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\, 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855860__net_1\, 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, 
        \I5.N_64_adt_net_855868__net_1\, 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\, 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\, 
        \I3.N_318_adt_net_855884__net_1\, 
        \I3.N_318_adt_net_855888__net_1\, 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        \I2.TEMPF_adt_net_855740__adt_net_855896__net_1\
         : std_logic;

begin 


    \I3.VDBi_40l1r\ : MUX2L
      port map(A => \I3.N_339\, B => \I3.N_133\, S => 
        \I3.N_354_0_adt_net_855368__net_1\, Y => 
        \I3.VDBi_40l1r_net_1\);
    
    \I2.DTE_21_1_IV_0L10R_1302\ : AO21
      port map(A => \I2.DT_TEMPl10r_net_1\, B => \I2.N_4038\, C
         => \I2.DTE_21_1l10r_adt_net_38511_\, Y => 
        \I2.DTE_21_1l10r_adt_net_38525_\);
    
    \I2.CHAINB_ERRS_525\ : MUX2L
      port map(A => \I2.CHAINB_ERRS_net_1\, B => 
        \I2.CHAINB_ERRF1_net_1\, S => 
        \I2.N_3876_adt_net_855252__net_1\, Y => 
        \I2.CHAINB_ERRS_525_net_1\);
    
    \I5.un1_SENS_ADDR_1_I_13\ : XOR2
      port map(A => \I5.DWACT_ADD_CI_0_TMPl0r\, B => 
        \I5.SENS_ADDRl1r_net_1\, Y => \I5.I_13\);
    
    \I2.L2TYPE_604\ : MUX2L
      port map(A => \I2.L2TYPEl15r_net_1\, B => \I2.L2TYPE_4l15r\, 
        S => \I2.N_4482_0\, Y => \I2.L2TYPE_604_net_1\);
    
    \I2.TOKENB_CNT_3_0_a3l0r\ : AND2
      port map(A => \I2.N_177\, B => 
        \I2.DWACT_ADD_CI_0_partial_suml0r\, Y => 
        \I2.TOKENB_CNT_3l0r\);
    
    \I2.END_EVNT2_1142\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT1_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT2_404\);
    
    \I2.ADOl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l11r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl11r);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I46_Y_1675\ : AND2FT
      port map(A => \I2.LSRAM_OUTl17r\, B => 
        \I2.PIPE7_DTl17r_net_1\, Y => \I2.N296_0_adt_net_86398_\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2200\ : AO21
      port map(A => \I3.RAMDTSl13r_net_1\, B => \I3.N_2034\, C
         => \I3.VDBi_57l13r_adt_net_140593_\, Y => 
        \I3.VDBi_57l13r_adt_net_140595_\);
    
    \I2.un1_STATE3_0\ : OR2
      port map(A => \I2.STATE3l5r_net_1\, B => 
        \I2.STATE3l6r_net_1\, Y => \I2.un1_STATE3\);
    
    \I1.REG_1_sqmuxa_adt_net_855388_\ : BFR
      port map(A => \I1.REG_1_sqmuxa\, Y => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\);
    
    \I1.REG_1_173\ : MUX2H
      port map(A => \REGl272r\, B => \I1.REG_74l272r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y => 
        \I1.REG_1_173_net_1\);
    
    \I2.PIPE5_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_705_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl29r_net_1\);
    
    \I5.sstate2l4r\ : DFFS
      port map(CLK => CLK_c, D => \I5.sstate2_ns_el0r\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate2l4r_net_1\);
    
    \I2.ROFFSET_915\ : MUX2H
      port map(A => \I2.ROFFSETl3r_net_1\, B => 
        \I2.ROFFSET_n3_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_915_net_1\);
    
    \I2.PHASE_864\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_C_242);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I27_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl6r\, B => \I2.PIPE7_DTL6R_699\, 
        Y => \I2.N249_0\);
    
    REGl326r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_227_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl326r\);
    
    \I3.TCNT3_n4\ : XOR2
      port map(A => \I3.TCNT3_i_0_il4r_net_1\, B => \I3.TCNT3_c3\, 
        Y => \I3.TCNT3_n4_net_1\);
    
    DPR_padl15r : IB33
      port map(PAD => DPR(15), Y => DPR_cl15r);
    
    \I1.REG_74_0_IV_0L223R_2004\ : AND2
      port map(A => \REGl223r\, B => \I1.N_97\, Y => 
        \I1.REG_74l223r_adt_net_128394_\);
    
    \I2.UN1_ERR_WORDS_RDY_0_SQMUXA_0_0_A5_1031\ : AND2
      port map(A => \I2.BITCNT_c0\, B => \I2.BITCNT_i_0_il4r\, Y
         => \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23152_\);
    
    \I2.DT_SRAM_0l1r\ : MUX2L
      port map(A => \I2.PIPE10_DTl1r_net_1\, B => 
        \I2.PIPE5_DTl1r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, Y => 
        \I2.N_869\);
    
    \I2.EVNT_NUM_n0\ : NOR2
      port map(A => EV_RES_C_569, B => \I2.EVNT_NUMl0r_net_1\, Y
         => \I2.EVNT_NUM_n0_net_1\);
    
    \I3.VDBOFFB_30_IV_0L4R_2405\ : AND2
      port map(A => \REGl289r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162326_\);
    
    \I2.STATE3_ns_o3_0l8r\ : OR2
      port map(A => \I2.N_3012_adt_net_24321_\, B => 
        \I2.N_3012_adt_net_24327_\, Y => \I2.N_3012\);
    
    \I3.TCNT4_386\ : MUX2H
      port map(A => \I3.TCNT4_i_0_il2r_net_1\, B => 
        \I3.TCNT4_n2_net_1\, S => \I3.TICKl2r_net_1\, Y => 
        \I3.TCNT4_386_net_1\);
    
    \I3.REG_1_154\ : MUX2L
      port map(A => VDB_inl5r, B => REGl53r, S => 
        \I3.N_1935_adt_net_855332__net_1\, Y => \I3.REG_1_154_0\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_804\ : NOR3
      port map(A => \I2.N_4646_1_ADT_NET_19635__185\, B => 
        \I2.N_4646_1_adt_net_19637_Rd1__net_1\, C => 
        \I2.END_EVNT2_404\, Y => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__182\);
    
    \I1.N_193_adt_net_118653_\ : NOR2
      port map(A => \I1.REG_74_1_396_m7_i_3\, B => 
        \I1.REG_74_8_0_N_6_i_i_0\, Y => 
        \I1.N_193_adt_net_118653__net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I140_Y_0_O2_1_1559\ : 
        OR3FFT
      port map(A => \I2.N_107_0\, B => \I2.N_13_1\, C => 
        \I2.N_95_0\, Y => \I2.N_74_adt_net_55281_\);
    
    \I2.DT_TEMP_776\ : MUX2H
      port map(A => \I2.DT_TEMPl15r_net_1\, B => 
        \I2.DT_TEMP_7l15r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_776_net_1\);
    
    \I2.REG_1_n1_0\ : XOR2
      port map(A => REGl33r, B => \I2.N_3829\, Y => 
        \I2.REG_1_n1_0_net_1\);
    
    \I1.REG_1_119\ : MUX2H
      port map(A => \REGl218r\, B => \I1.REG_74l218r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_119_net_1\);
    
    \I2.DTE_21_1_IV_0L13R_1287\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.N_44_i_0\, C => 
        \I2.DTE_21_1l13r_adt_net_38169_\, Y => 
        \I2.DTE_21_1l13r_adt_net_38180_\);
    
    \I2.BNCID_VECT_tile_0_I_5\ : DFF
      port map(CLK => CLK_c, D => \I2.TDCTRG_c_i_0\, Q => 
        \I2.N_11\);
    
    \I2.MAJORITY_REG_I_0L1R_895\ : NOR2
      port map(A => \I2.MIC_REG3L1R_454\, B => 
        \I2.MIC_REG1L1R_455\, Y => \I2.N_3877_adt_net_4723_\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2526\ : OR3
      port map(A => \I3.N_2070_adt_net_163505_\, B => 
        \I3.N_2070_adt_net_163499_\, C => 
        \I3.N_2070_adt_net_163500_\, Y => 
        \I3.N_2070_adt_net_163509_\);
    
    \I2.PIPE10_DT_17_il14r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l1r_net_1\, C => \I2.PIPE10_DT_17_i_0l14r_net_1\, 
        Y => \I2.N_3800\);
    
    REGl302r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_203_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl302r\);
    
    \I3.VDBOFFA_31_IV_0L0R_2630\ : AO21
      port map(A => \REGl269r\, B => \I3.REGMAPl31r_net_1\, C => 
        \I3.VDBoffa_31l0r_adt_net_164614_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164643_\);
    
    \I2.DT_TEMP_778\ : MUX2H
      port map(A => \I2.DT_TEMPl17r_net_1\, B => 
        \I2.DT_TEMP_7l17r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_778_net_1\);
    
    \I2.END_EVNT2_1512\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT1_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT2_619\);
    
    \I2.L2TYPEl12r_1545\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_601_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL12R_652\);
    
    \I3.VADm_0_a3l2r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl2r_net_1\, Y => \I3.VADml2r\);
    
    \I2.MIC_ERR_REGSl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_341_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl12r_net_1\);
    
    \I2.BNCID_VECTror_adt_net_48223_\ : AND2
      port map(A => \I2.BNCID_VECTra13_1_net_1\, B => 
        \I2.BNCID_VECTro_1\, Y => 
        \I2.BNCID_VECTror_adt_net_48223__net_1\);
    
    \I2.L2TYPEl8r_1543\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_597_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL8R_650\);
    
    \I2.L2ARR_942\ : MUX2L
      port map(A => \I2.L2ARRl2r_net_1\, B => \I2.L2ARR_n2_net_1\, 
        S => \I2.N_4482_0\, Y => \I2.L2ARR_942_net_1\);
    
    \I1.N_349_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_349_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_349_Rd1__net_1\);
    
    \I3.UN15_ANYCYC_2298\ : NOR2
      port map(A => \I3.PIPEAl29r_net_1\, B => 
        \I3.PIPEAl31r_net_1\, Y => 
        \I3.un15_anycyc_adt_net_147616_\);
    
    \I2.DTO_1_899\ : MUX2L
      port map(A => \I2.DTO_1l25r_Rd1__net_1\, B => 
        \I2.DTO_16_1l25r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834756_Rd1__net_1\, Y
         => \I2.DTO_1l25r\);
    
    \I3.VDBi_57_0_iv_0_a3_8_1l15r\ : AND3FFT
      port map(A => \I3.N_1905_1_adt_net_855384__net_1\, B => 
        \I3.N_2015\, C => \I3.REGMAPl9r_adt_net_854324__net_1\, Y
         => \I3.N_402_1\);
    
    \I1.REG_74_7_i_a2_a0_0_1l404r_918\ : NOR2
      port map(A => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__19\, 
        B => \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Rd1__net_1\, Y
         => \I1.N_232_1_296\);
    
    \I1.SBYTE_8_0_a2_i_m2l4r\ : MUX2L
      port map(A => \FBOUTl3r\, B => REGl87r, S => 
        \I1.sstatel2r_net_1\, Y => \I1.N_1386\);
    
    \I2.PIPE1_DT_42_1_ivl19r\ : OR3
      port map(A => \I2.PIPE1_DT_42l19r_adt_net_47249_\, B => 
        \I2.PIPE1_DT_42l19r_adt_net_47261_\, C => 
        \I2.PIPE1_DT_42l19r_adt_net_47262_\, Y => 
        \I2.PIPE1_DT_42l19r\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855400_\ : BFR
      port map(A => \I1.N_50_0_adt_net_1409__net_1\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\);
    
    \I1.REG_1_176\ : MUX2H
      port map(A => \REGl275r\, B => \I1.REG_74l275r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y => 
        \I1.REG_1_176_net_1\);
    
    \I2.STATE2l0r_1480\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.WPAGEe_adt_net_855056__net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.STATE2L0R_587\);
    
    \I2.SRAM_EVNT_c3_i_o2\ : NAND2
      port map(A => \I2.N_3858\, B => \I2.SRAM_EVNTl3r_net_1\, Y
         => \I2.N_3860\);
    
    \I2.FIRST_TDC_675_1589\ : NOR2FT
      port map(A => \I2.FIRST_TDC_i_0_i\, B => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__169\, Y => 
        \I2.FIRST_TDC_675_adt_net_61236_\);
    
    \I2.G_EVNT_NUM_n8_i\ : NOR3
      port map(A => EV_RES_C_569, B => \I2.N_282\, C => 
        \I2.N_207\, Y => \I2.N_4640\);
    
    \I3.PIPEA_8l12r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854476__net_1\, B => 
        \I3.N_221\, Y => \I3.PIPEA_8l12r_net_1\);
    
    \I3.VDBoffal0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_44_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal0r_net_1\);
    
    \I3.SELBASE32\ : LD
      port map(EN => ASB_c, D => \I3.un6_asb_NE_net_1\, Q => 
        \I3.SELBASE32_net_1\);
    
    \I3.PIPEBl11r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_90_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl11r_net_1\);
    
    \I3.PIPEA_8_0l11r\ : MUX2L
      port map(A => DPR_cl11r, B => \I3.PIPEA1l11r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855352__net_1\, Y => \I3.N_220\);
    
    TDCGDB_pad : OB33PH
      port map(PAD => TDCGDB, A => TDCGDB_c);
    
    \I1.ISCK_0_sqmuxa_0_0_a2_1233\ : NAND3FFT
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__861\, B => 
        \I1.N_359\, C => \I1.sstatel4r_net_1\, Y => 
        \I1.N_656_495\);
    
    \I2.G_EVNT_NUMl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_924_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl10r_net_1\);
    
    \I2.MIC_ERR_REGSl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_331_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl2r_net_1\);
    
    \I3.UN10_TCNT2_2107\ : OR3
      port map(A => \I3.TCNT2_i_0_il6r_net_1\, B => 
        \I3.TCNT2l5r_net_1\, C => \I3.un10_tcnt2_adt_net_135286_\, 
        Y => \I3.un10_tcnt2_adt_net_135290_\);
    
    \I2.LSRAM_RDi\ : DFFS
      port map(CLK => CLK_c, D => \I2.LSRAM_RDi_486_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_RDi_net_1\);
    
    \I2.PIPE6_DTl33r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_487_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl33r_net_1\);
    
    \I1.REG_74_1l276r\ : NOR3FFT
      port map(A => \I1.N_273_5_i\, B => 
        \I1.N_273_6_i_0_adt_net_854796__net_1\, C => 
        \I1.N_201_9_188\, Y => \I1.REG_74_1l268r\);
    
    \I2.N_182_adt_net_1007_\ : OR2
      port map(A => \I2.STATE2l0r_net_1\, B => 
        \I2.STATE2_nsl2r_adt_net_24911_\, Y => 
        \I2.N_182_adt_net_1007__net_1\);
    
    \I2.PIPE5_DTl21r_1519\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_697_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL21R_626\);
    
    \I1.PAGECNTl7r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_320_adt_net_854876__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTl7r_net_1\);
    
    \I3.VDBoff_4_i_il1r\ : MUX2L
      port map(A => \I3.VDBoffbl1r_net_1\, B => 
        \I3.VDBoffal1r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_2065\);
    
    \I3.STATE1_ns_0_iv_0_0_o2l6r\ : AO21FTT
      port map(A => \I3.ASBS_net_1\, B => \I3.STATE1_ipl5r\, C
         => \I3.STATE1_ipl4r\, Y => \I3.N_1920\);
    
    TDCDB_padl4r : IB33
      port map(PAD => TDCDB(4), Y => TDCDB_cl4r);
    
    \I3.PIPEA_235\ : MUX2L
      port map(A => \I3.PIPEAl4r_net_1\, B => 
        \I3.PIPEA_8l4r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854676__net_1\, Y
         => \I3.PIPEA_235_net_1\);
    
    \I1.REG_74_12l268r\ : AO21FTF
      port map(A => \I1.N_73_10_adt_net_117095_\, B => 
        \I1.N_145_12_adt_net_123140_\, C => \I1.N_232_1\, Y => 
        \I1.N_145_12\);
    
    \I3.PIPEAl28r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEA_259_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl28r_net_1\);
    
    \I3.VDBI_57_0_IV_0L19R_2173\ : AO21
      port map(A => REGl67r, B => \I3.N_1839\, C => 
        \I3.VDBi_57l19r_adt_net_139387_\, Y => 
        \I3.VDBi_57l19r_adt_net_139392_\);
    
    \I2.SUB8_508\ : MUX2H
      port map(A => \I2.SUB8l5r_net_1\, B => \I2.SUB8_2l5r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855148__net_1\, Y => 
        \I2.SUB8_508_net_1\);
    
    \I4.un4_bcnt_I_13\ : XOR2
      port map(A => \I4.bcntl3r_net_1\, B => \I4.N_4_0\, Y => 
        \I4.I_13_0\);
    
    \I2.BNCID_VECTror_10_tz_0\ : AO21
      port map(A => \I2.BNCID_VECTra13_1_net_1\, B => 
        \I2.BNCID_VECTro_5\, C => 
        \I2.BNCID_VECTror_10_tz_0_adt_net_48139_\, Y => 
        \I2.BNCID_VECTror_10_tz_0_net_1\);
    
    \I3.majority_5_un102_reg\ : XOR2FT
      port map(A => \I3.REG2l5r_net_1\, B => \I3.REG1l5r_net_1\, 
        Y => \I3.un102_reg\);
    
    \I2.OFFSET_37_8l0r\ : MUX2L
      port map(A => \REGl357r\, B => \REGl293r\, S => 
        \I2.PIPE7_DTL27R_74\, Y => \I2.N_691\);
    
    \I1.REG_74_8_0_o4_0l380r_814\ : NAND2
      port map(A => \I1.N_1366\, B => \I1.N_1367_i\, Y => 
        \I1.N_396_192\);
    
    \I3.un22_bltcyc_0_a3\ : OR2
      port map(A => \I3.MBLTCYC_423\, B => \I3.BLTCYC_net_1\, Y
         => \I3.un22_bltcyc\);
    
    \I2.DTO_16_1l19r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l19r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l19r_Rd1__net_1\);
    
    \I1.BYTECNT_n2_i_o2\ : AND2
      port map(A => \I1.BYTECNTl2r_net_1\, B => 
        \I1.N_323_adt_net_108906_\, Y => \I1.N_323\);
    
    \I2.PIPE5_DT_6_0l7r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l7r\, B => 
        \I2.un27_pipe5_dt0l7r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1076\);
    
    \I2.PIPE8_DT_551\ : MUX2L
      port map(A => \I2.PIPE8_DTl23r_net_1\, B => 
        \I2.PIPE8_DT_21l23r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_551_net_1\);
    
    \I1.REG_74_0_ivl350r\ : AO21
      port map(A => \REGl350r\, B => \I1.N_225\, C => 
        \I1.REG_74l350r_adt_net_116117_\, Y => \I1.REG_74l350r\);
    
    \I2.FID_7_IVL3R_1728\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl3r_net_1\, 
        C => \I2.FID_7l3r_adt_net_93251_\, Y => 
        \I2.FID_7l3r_adt_net_93259_\);
    
    \I2.ADE_4l9r\ : MUX2H
      port map(A => \I2.WOFFSETl10r\, B => \I2.ROFFSETl10r_net_1\, 
        S => NOESRAME_c, Y => \I2.ADE_4l9r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL8R_1472\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl24r_net_1\, Y => 
        \I2.PIPE1_DT_42l8r_adt_net_50426_\);
    
    \I2.FID_7_0_ivl8r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl8r_net_1\, 
        C => \I2.FID_7l8r_adt_net_92747_\, Y => \I2.FID_7l8r\);
    
    \I2.CRC32_12_il2r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_73_i_0_i_0\, Y => 
        \I2.N_3919\);
    
    \I2.CRC32_12_0_0_x2l23r\ : XOR2FT
      port map(A => \I2.CRC32l23r_net_1\, B => \I2.N_4269_i_i\, Y
         => \I2.N_129_i_0_i_0\);
    
    \I3.VDBi_40_sn_m2_0_751\ : NOR2
      port map(A => \I3.REGMAPL57R_50\, B => 
        \I3.REGMAP_i_0_il58r_net_1\, Y => \I3.N_354_0_129\);
    
    \I2.MIC_ERR_REGSl47r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_376_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl47r_net_1\);
    
    VDB_padl9r : IOB33PH
      port map(PAD => VDB(9), A => \I3.VDBml9r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl9r);
    
    \I2.L2TYPE_4_il6r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4446_adt_net_67934_\, C => 
        \I2.N_4446_adt_net_67977_\, Y => \I2.N_4446\);
    
    \I3.TICKil0r_1450\ : DFFC
      port map(CLK => CLK_c, D => \I3.un6_tcnt1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TICKL0R_557);
    
    \I1.BITCNTLDE_I_A2_0_1774\ : AND3FFT
      port map(A => \I1.N_362\, B => \I1.N_349_Rd1__net_1\, C => 
        \I1.N_628_adt_net_107115_\, Y => 
        \I1.N_68_adt_net_108395_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I143_Y_0\ : XOR2
      port map(A => \I2.N_3539_i_i\, B => \I2.G_1_2\, Y => 
        \I2.ADD_18x18_fast_I143_Y_0\);
    
    \I2.un1_END_EVNT1_0_sqmuxa_i_0\ : OR2
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\, 
        B => \I2.N_3234_adt_net_21449_\, Y => \I2.N_3234\);
    
    \I1.REG_74_0_ivl337r\ : AO21
      port map(A => \REGl337r\, B => \I1.N_209\, C => 
        \I1.REG_74l337r_adt_net_117486_\, Y => \I1.REG_74l337r\);
    
    \I2.DTO_16_1_IV_0L31R_1065\ : AND2FT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        B => \I2.DT_TEMPl31r_net_1\, Y => 
        \I2.DTO_16_1l31r_adt_net_28248_\);
    
    \I2.PIPE1_DT_12l1r\ : MUX2H
      port map(A => \I2.TDCDASl20r_net_1\, B => 
        \I2.TDCDASl1r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092__net_1\, Y
         => \I2.PIPE1_DT_12l1r_net_1\);
    
    \I2.STATE1_ns_i_o2l9r_965\ : OR3
      port map(A => FLUSH, B => \I2.FCNT_c1\, C => 
        \I2.FCNTL2R_599\, Y => \I2.N_3272_343\);
    
    \I2.NWPIPE6_449\ : MUX2H
      port map(A => \I2.un1_NWPIPE5_1_i\, B => \I2.NWPIPE6_net_1\, 
        S => END_FLUSH_560, Y => \I2.NWPIPE6_449_net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2460\ : AND2
      port map(A => \REGl318r\, B => \I3.REGMAPl37r_net_1\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162900_\);
    
    \I2.un2_evnt_word_I_73\ : XOR2
      port map(A => \I2.N_4\, B => \I2.WOFFSETl12r\, Y => 
        \I2.I_73\);
    
    \I3.PIPEA1_12l18r\ : AND2
      port map(A => DPR_cl18r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854500__net_1\, Y => 
        \I3.PIPEA1_12l18r_net_1\);
    
    \I3.REG_1_182\ : MUX2L
      port map(A => VDB_inl1r, B => \I3.REGl134r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, Y => 
        \I3.REG_1_182_0\);
    
    \I3.VDBoffbl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_56_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl4r_net_1\);
    
    \I3.VDBi_57_0_ivl28r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l28r_net_1\, C
         => \I3.VDBi_57l28r_adt_net_138311_\, Y => 
        \I3.VDBi_57l28r\);
    
    \I2.NLD_647\ : OAI21FTF
      port map(A => NLD_c, B => \I2.STATE3l13r_net_1\, C => 
        \I2.STATE3l5r_net_1\, Y => \I2.NLD_647_net_1\);
    
    \I2.PIPE10_DT_622\ : MUX2L
      port map(A => \I2.PIPE10_DTl17r_net_1\, B => \I2.N_3803\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_622_net_1\);
    
    \I2.STATEe_nsl3r\ : OR2
      port map(A => \I2.STATEe_nsl3r_adt_net_22965_\, B => 
        \I2.STATEe_nsl3r_adt_net_22967_\, Y => 
        \I2.STATEe_nsl3r_net_1\);
    
    \I2.REG_1l33r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n1_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl33r);
    
    \I3.REG_1_186\ : MUX2L
      port map(A => VDB_inl5r, B => \I3.REGl138r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, Y => 
        \I3.REG_1_186_0\);
    
    \I2.CRC32_12_0_0_m2l23r\ : MUX2H
      port map(A => \I2.DT_SRAMl23r_net_1\, B => 
        \I2.DT_TEMPl23r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854428__net_1\, Y => 
        \I2.N_4269_i_i\);
    
    \I3.VDBi_57_iv_0_0_o2_0_7l0r\ : OR3
      port map(A => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146451_\, B => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146426_\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146450_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r\);
    
    \I2.PIPE1_DT_30l4r\ : MUX2L
      port map(A => \I2.TDCDBSl4r_net_1\, B => 
        \I2.TDCDBSl2r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, Y
         => \I2.PIPE1_DT_30l4r_net_1\);
    
    \I3.REGMAPL9R_3029\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un41_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL9R_783\);
    
    \I2.BNC_IDl10r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_56_0\, CLR => 
        \I2.N_4617_i_0\, SET => \I2.N_4616_i_0\, Q => 
        \I2.BNC_IDl10r_net_1\);
    
    \I3.STATE1_ns_0_iv_0_o2_0_i_a2_0_0_o2l7r\ : AND2
      port map(A => \I3.N_560\, B => \I3.N_2083_adt_net_134513_\, 
        Y => \I3.N_2083\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I207_Y\ : XOR2FT
      port map(A => \I2.N498_1\, B => 
        \I2.SUB_21x21_fast_I207_Y_0\, Y => \I2.SUB8_2l11r\);
    
    \I2.MIC_REG3l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_324_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l7r_net_1\);
    
    \I1.BYTECNT_n7_i_0\ : AND2FT
      port map(A => \I1.N_223_adt_net_854848__net_1\, B => 
        \I1.N_79_adt_net_109340_\, Y => \I1.N_79\);
    
    REGl187r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_88_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl187r\);
    
    \I2.OFFSET_37_1l7r\ : MUX2L
      port map(A => \REGl356r\, B => \REGl292r\, S => 
        \I2.PIPE7_DTL27R_64\, Y => \I2.N_642\);
    
    \I1.N_238_RD1__2882\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_238_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_238_RD1__314\);
    
    \I3.VDBi_57_0_iv_0_0l8r\ : OR3
      port map(A => \I3.VDBi_57l8r_adt_net_142784_\, B => 
        \I3.VDBi_57l8r_adt_net_142792_\, C => 
        \I3.VDBi_57l8r_adt_net_142793_\, Y => \I3.VDBi_57l8r\);
    
    \REG_i_il5r_adt_net_855560_\ : BFR
      port map(A => REG_i_il5r, Y => 
        \REG_i_il5r_adt_net_855560__net_1\);
    
    \I2.N_4667_1_ADT_NET_1046__2757\ : OAI21FTF
      port map(A => \I2.N_4261\, B => \I2.N_4283_I_0_43\, C => 
        \I2.STATE2l2r_adt_net_855212__net_1\, Y => 
        \I2.N_4667_1_ADT_NET_1046__33\);
    
    \I2.UN1_NWPIPE7_2_1669\ : AND2
      port map(A => \I2.PIPE7_DTL27R_64\, B => 
        \I2.PIPE7_DTL26R_348\, Y => 
        \I2.un1_NWPIPE7_2_adt_net_73604_\);
    
    \I3.un29_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.un227_reg_ads_2\, B => \I3.N_573\, Y => 
        \I3.un29_reg_ads_0_a2_0_a3_net_1\);
    
    DTO_padl25r : IOB33PH
      port map(PAD => DTO(25), A => \I2.DTO_1l25r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl25r);
    
    \I1.sstate_tr19_0_a2_0_a4\ : AND2FT
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.sstatel5r_net_1\, Y => \I1.sstate_nsl6r\);
    
    \I3.PIPEA1l3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_301_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l3r_net_1\);
    
    \I3.REGMAPl43r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un196_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAPl43r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I161_Y\ : AND2FT
      port map(A => \I2.I161_un1_Y\, B => 
        \I2.N486_i_adt_net_89208_\, Y => \I2.N486_i\);
    
    \I3.VDBi_57l2r_adt_net_145227_\ : AO21
      port map(A => REGl18r, B => \I3.N_2053\, C => 
        \I3.VDBi_57l2r_adt_net_145226__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145227__net_1\);
    
    \I2.OFFSET_37_17l2r\ : MUX2L
      port map(A => \I2.N_757\, B => \I2.N_749\, S => 
        \I2.PIPE7_DTL26R_354\, Y => \I2.N_765\);
    
    \I5.sstate1se_10_0_0_o4\ : NOR2
      port map(A => \I5.sstate1l6r_net_1\, B => 
        \I5.sstate1l3r_net_1\, Y => \I5.N_77\);
    
    \I2.PIPE5_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_691_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl15r_net_1\);
    
    \I1.SBYTE_62\ : MUX2L
      port map(A => \FBOUTl4r\, B => \I1.N_192\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_62_net_1\);
    
    \I1.LUT_0_sqmuxa_i_0_o2\ : NAND3
      port map(A => \I1.BYTECNTl8r_net_1\, B => 
        \I1.N_341_Rd1__net_1\, C => \I1.N_328_I_0_497\, Y => 
        \I1.N_359\);
    
    \I2.DTE_21_1_0_IVL31R_1227\ : AO21FTT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_289\, B => 
        \I2.DT_SRAMl31r_net_1\, C => 
        \I2.DTE_21_1l31r_adt_net_36411_\, Y => 
        \I2.DTE_21_1l31r_adt_net_36416_\);
    
    \I1.REG_74_13_0_a2l404r\ : NOR2FT
      port map(A => \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, 
        B => \I1.N_240\, Y => \I1.N_584\);
    
    SCLA_pad : OB33PH
      port map(PAD => SCLA, A => \I5.N_107\);
    
    \I2.LSRAM_RADDRl2r\ : MUX2L
      port map(A => \LSRAM_FL_RADDRl2r\, B => 
        \I2.LSRAM_RADDRil2r_net_1\, S => FLUSH, Y => 
        \I2.LSRAM_RADDRl2r_net_1\);
    
    \I2.WOFFSETl11r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl11r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl11r_Rd1__net_1\);
    
    \I3.un81_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_582\, B => \I3.N_553\, Y => 
        \I3.un81_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I41_Y\ : AND2
      port map(A => \I2.N238\, B => \I2.N241\, Y => \I2.N306\);
    
    \I3.VDBI_57_IVL1R_2269\ : AO21
      port map(A => 
        \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344__net_1\, 
        B => \I3.VDBi_52l1r_net_1\, C => 
        \I3.VDBi_57l1r_adt_net_145946_\, Y => 
        \I3.VDBi_57l1r_adt_net_145947_\);
    
    \I2.un1_END_EVNT1_0_sqmuxa_i_0_o2\ : AND2FT
      port map(A => \I2.SRAM_FULL_net_1\, B => \I2.GIROT_net_1\, 
        Y => \I2.N_3882\);
    
    \I2.DTO_16_1_IV_0_0L12R_1161\ : AO21
      port map(A => \I2.DTO_1l12r\, B => \I2.N_196\, C => 
        \I2.DTO_16_1l12r_adt_net_32632_\, Y => 
        \I2.DTO_16_1l12r_adt_net_32634_\);
    
    \I3.REGMAPl51r_1616\ : DFF
      port map(CLK => CLK_c, D => \I3.un7_ronly_0_a2_0_a3_net_1\, 
        Q => \I3.REGMAPL51R_723\);
    
    \I2.PIPE6_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_461_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl7r_net_1\);
    
    \I2.DTO_1_890\ : MUX2L
      port map(A => \I2.DTO_1l16r_Rd1__net_1\, B => 
        \I2.DTO_16_1l16r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834764_Rd1__net_1\, Y
         => \I2.DTO_1l16r\);
    
    \I1.REG_1_93\ : MUX2H
      port map(A => \REGl192r\, B => \I1.REG_74l192r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\, Y => 
        \I1.REG_1_93_net_1\);
    
    ADE_padl6r : OB33PH
      port map(PAD => ADE(6), A => ADE_cl6r);
    
    DTE_padl6r : IOB33PH
      port map(PAD => DTE(6), A => \I2.DTE_1l6r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl6r);
    
    \I2.RAMAD_4_0l17r\ : MUX2H
      port map(A => \I2.RAMAD1l17r_net_1\, B => RAMAD_VMEl17r, S
         => \REG_i_il5r_adt_net_855552__net_1\, Y => \I2.N_544\);
    
    \I3.VADm_0_a3l0r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl0r_net_1\, Y => \I3.VADml0r\);
    
    \I2.MIC_ERR_REGSl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_337_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl8r_net_1\);
    
    VDB_padl18r : IOB33PH
      port map(PAD => VDB(18), A => \I3.VDBml18r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl18r);
    
    \I2.G_EVNT_NUMlde_i_a2\ : NOR2
      port map(A => EV_RES_C_567, B => \I2.INC_EVNT_NUM_net_1\, Y
         => \I2.N_3769\);
    
    \I3.VDBml15r\ : MUX2L
      port map(A => \I3.VDBil15r_net_1\, B => \I3.N_157\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml15r_net_1\);
    
    \I2.PIPE7_DTL26R_2902\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_356\);
    
    \I5.SCL_1_i_a2_0_1\ : NAND3FFT
      port map(A => \I5.sstate1l2r_net_1\, B => 
        \I5.sstate1l10r_net_1\, C => \I5.N_81_i_0_i\, Y => 
        \I5.SCL_1_i_a2_0_1_net_1\);
    
    \I2.N_2358_tz_tz_adt_net_854956_\ : BFR
      port map(A => \I2.N_2358_tz_tz\, Y => 
        \I2.N_2358_tz_tz_adt_net_854956__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I34_P0N_1283\ : OR2FT
      port map(A => \I2.LSRAM_OUTl13r\, B => 
        \I2.PIPE7_DTl13r_net_1\, Y => \I2.N270_0_545\);
    
    \I2.MIC_ERR_REGS_371\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl43r_net_1\, B => 
        \I2.MIC_ERR_REGSl42r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_371_net_1\);
    
    \I3.VDBI_57_0_IV_0L21R_2163\ : AND2FT
      port map(A => \I3.N_1917_adt_net_855336__net_1\, B => 
        \I3.REGl154r\, Y => \I3.VDBi_57l21r_adt_net_139179_\);
    
    \I1.sstate_ns_1_iv_0_il8r\ : AND2FT
      port map(A => 
        \PULSEl0r_adt_net_854532__adt_net_855544__net_1\, B => 
        \I1.N_289_adt_net_107403_\, Y => \I1.N_289\);
    
    \I2.MIC_REG1l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_303_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1l2r_net_1\);
    
    VDB_padl5r : IOB33PH
      port map(PAD => VDB(5), A => VDBm_i_i_m2l5r, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl5r);
    
    \I3.REG_1l91r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_272_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl91r\);
    
    \I2.N_64_0_adt_net_855028_\ : BFR
      port map(A => \I2.N_64_0\, Y => 
        \I2.N_64_0_adt_net_855028__net_1\);
    
    \I2.TDCDASl28r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl28r, Q => 
        \I2.TDCDASl28r_net_1\);
    
    RAMAD_padl9r : OB33PH
      port map(PAD => RAMAD(9), A => RAMAD_cl9r);
    
    \I3.VDBi_40_1l9r\ : MUX2L
      port map(A => REGl126r, B => \I3.VDBi_31l9r_net_1\, S => 
        \I3.REGMAPl16r_net_1\, Y => \I3.N_347\);
    
    \I3.VDBoffl6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_122_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl6r_net_1\);
    
    \I3.STATE1_ILLEGAL_2135\ : XOR2FT
      port map(A => \I3.STATE1_ipl0r_adt_net_854356__net_1\, B
         => \I3.N_1189\, Y => \I3.N_1193_ip_adt_net_136558_\);
    
    \I2.DT_TEMPl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_786_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl25r_net_1\);
    
    \I2.STATE2l0r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.WPAGEe_adt_net_855056__net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.STATE2l0r_net_1\);
    
    \I2.L2TYPEl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_599_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl10r_net_1\);
    
    \I2.PIPE7_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl7r_net_1\);
    
    \I1.N_592_adt_net_854756_\ : BFR
      port map(A => \I1.N_592\, Y => 
        \I1.N_592_adt_net_854756__net_1\);
    
    \I2.DTE_21_1_iv_0l9r\ : OR3
      port map(A => \I2.DTE_21_1l9r_adt_net_38627_\, B => 
        \I2.DTE_21_1l9r_adt_net_38635_\, C => 
        \I2.DTE_21_1l9r_adt_net_38636_\, Y => \I2.DTE_21_1l9r\);
    
    \I2.un1_TOKENB_CNT_I_1\ : AND2
      port map(A => TICKL0R_557, B => \I2.TOKENB_CNTl0r_net_1\, Y
         => \I2.DWACT_ADD_CI_0_TMP_1l0r\);
    
    \I3.VDBOFFB_30_IV_0L7R_2354\ : AND2
      port map(A => \REGl308r\, B => \I3.REGMAPl35r_net_1\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161768_\);
    
    VDB_padl31r : IOB33PH
      port map(PAD => VDB(31), A => \I3.VDBml31r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl31r);
    
    \I2.OFFSET_37_3l4r\ : MUX2L
      port map(A => \I2.N_647\, B => \I2.N_639\, S => 
        \I2.PIPE7_DTL26R_349\, Y => \I2.N_655\);
    
    \I2.SUB9_1_ADD_18x18_fast_I2_P0N\ : OR2
      port map(A => \I2.N_3537_i_i\, B => \I2.G_1_3\, Y => 
        \I2.N232\);
    
    TDCDB_padl25r : IB33
      port map(PAD => TDCDB(25), Y => TDCDB_cl25r);
    
    \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854404_\ : BFR
      port map(A => \I1.PAGECNT_0l8r_adt_net_834720_Rd1__net_1\, 
        Y => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854404__net_1\);
    
    \I2.PIPE1_DT_12l8r\ : MUX2L
      port map(A => \I2.TDCDASl8r_net_1\, B => 
        \I2.TDCDASl6r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, Y
         => \I2.PIPE1_DT_12l8r_net_1\);
    
    \I2.PIPE10_DT_17_i_0l13r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855596__net_1\, B => 
        \I2.PIPE9_DTl13r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l13r_net_1\);
    
    \I1.REG_74_0_ivl234r\ : AO21
      port map(A => \REGl234r\, B => \I1.N_105\, C => 
        \I1.REG_74l234r_adt_net_127280_\, Y => \I1.REG_74l234r\);
    
    \I3.PULSE_332_2294\ : AND2
      port map(A => PULSEl2r, B => 
        \I3.N_1409_adt_net_854744__net_1\, Y => 
        \I3.PULSE_332_adt_net_147433_\);
    
    \I3.VDBi_16_m_i_a2l3r\ : NOR3FTT
      port map(A => \I3.REGMAPL2R_737\, B => \I3.REGMAPL7R_460\, 
        C => \I3.REGMAPl3r_net_1\, Y => \I3.N_2053\);
    
    \I3.RAMAD_VME_32\ : MUX2H
      port map(A => RAMAD_VMEl8r, B => \I3.REGl91r\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_32_net_1\);
    
    \I2.CRC32l21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_816_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l21r_net_1\);
    
    \I2.MAJORITY_REG_I_IL6R_1220\ : OA21
      port map(A => \I2.MIC_REG3l6r_net_1\, B => 
        \I2.MIC_REG1_i_il6r_net_1\, C => \I2.MIC_REG2l6r_net_1\, 
        Y => \REGl28r_adt_net_36082_\);
    
    \I3.VDBOFFB_30_IV_0L7R_2356\ : AO21
      port map(A => \REGl324r\, B => \I3.REGMAPl37r_net_1\, C => 
        \I3.VDBoffb_30l7r_adt_net_161748_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161789_\);
    
    \I2.REG_1l32r_1126\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n0_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL32R_388);
    
    \I2.PIPE1_DT_42_1_IV_2L27R_1366\ : OAI21FTF
      port map(A => \I2.PIPE1_DT_2_SQMUXA_1_1_177\, B => 
        \I2.TDCDBSl27r_net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46027_\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46039_\);
    
    \I1.REG_74_22l404r_810\ : OR3FFT
      port map(A => \I1.REG_74_4_i_a2_404_N_4_i\, B => 
        \I1.N_347_adt_net_854792__net_1\, C => \I1.N_396_191\, Y
         => \I1.N_201_9_188\);
    
    \I2.OFFSET_37_17l5r\ : MUX2L
      port map(A => \I2.N_760\, B => \I2.N_752\, S => 
        \I2.PIPE7_DTL26R_352\, Y => \I2.N_768\);
    
    \I3.REG_1l49r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_150_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl49r);
    
    \I2.resyn_0_I2_TRGCNT_c1_i_a2_0\ : OR3
      port map(A => \I2.N_3794\, B => \I2.TRGCNTl0r_net_1\, C => 
        \I2.TRGCNT_i_0_il1r\, Y => \I2.N_3796\);
    
    \I3.VDBI_57_0_IV_0_0L8R_2226\ : AO21
      port map(A => \I3.VDBil8r_net_1\, B => \I3.N_56\, C => 
        \I3.VDBi_57l8r_adt_net_142786_\, Y => 
        \I3.VDBi_57l8r_adt_net_142793_\);
    
    RAMDT_padl7r : IOB33PH
      port map(PAD => RAMDT(7), A => \I1.RAMDT_SPI_1l0r_net_1\, 
        EN => \I1.RAMDT_SPI_e_net_1\, Y => RAMDT_inl7r);
    
    \I5.sstate1l11r\ : DFFC
      port map(CLK => CLK_c, D => \I5.N_100\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l11r_net_1\);
    
    \I2.STATE2l5r\ : DFFS
      port map(CLK => CLK_c, D => \I2.N_2796_i_0\, SET => 
        CLEAR_STAT_i_0, Q => \I2.STATE2l5r_net_1\);
    
    \I2.STATE1_i_1l8r\ : NOR2
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855244__net_1\, 
        B => \I2.N_3234_adt_net_21449_\, Y => \I2.N_3234_i_0\);
    
    \I2.DTO_16_1_IVL11R_1164\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855680__net_1\, B => 
        \I2.DTO_9l11r\, Y => \I2.DTO_16_1l11r_adt_net_32864_\);
    
    \I3.VDBOFFA_31_IV_0L1R_2602\ : AND2
      port map(A => \REGl230r\, B => \I3.REGMAPl26r_net_1\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164412_\);
    
    \I2.DTO_16_1_IV_0L9R_1175\ : AO21
      port map(A => \I2.N_457\, B => \I2.DTE_2_1l9r_net_1\, C => 
        \I2.DTO_16_1l9r_adt_net_33240_\, Y => 
        \I2.DTO_16_1l9r_adt_net_33251_\);
    
    \I1.REG_1_169\ : MUX2H
      port map(A => \REGl268r\, B => \I1.REG_74l268r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y
         => \I1.REG_1_169_net_1\);
    
    \I3.ADACKCYC\ : DFFC
      port map(CLK => CLK_c, D => \I3.ADACKCYC_112_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.ADACKCYC_net_1\);
    
    \I1.REG_1_125\ : MUX2H
      port map(A => \REGl224r\, B => \I1.REG_74l224r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\, Y => 
        \I1.REG_1_125_net_1\);
    
    \I2.DTO_16_1_IV_0L7R_1188\ : AO21
      port map(A => \I2.N_182_ADT_NET_1007__386\, B => 
        \I2.DT_SRAMl7r_net_1\, C => 
        \I2.DTO_16_1l7r_adt_net_33734_\, Y => 
        \I2.DTO_16_1l7r_adt_net_33735_\);
    
    \I2.FID_7_0_IVL19R_953\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl19r_net_1\, 
        Y => \I2.FID_7l19r_adt_net_17517_\);
    
    REGl382r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_283_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl382r\);
    
    \I3.VDBoffa_51\ : OR3
      port map(A => \I3.VDBoffa_51_adt_net_163358_\, B => 
        \I3.VDBoffa_31l7r_adt_net_163319_\, C => 
        \I3.VDBoffa_31l7r_adt_net_163320_\, Y => 
        \I3.VDBoffa_51_net_1\);
    
    \I2.RAMAD1l11r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_665_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l11r_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2401\ : OR3
      port map(A => \I3.VDBoffb_30l5r_adt_net_162177_\, B => 
        \I3.VDBoffb_30l5r_adt_net_162173_\, C => 
        \I3.VDBoffb_30l5r_adt_net_162174_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162180_\);
    
    \I2.PIPE2_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl29r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl29r_net_1\);
    
    \I1.BYTECNT_n2_i\ : AND2FT
      port map(A => \I1.N_223_adt_net_854844__net_1\, B => 
        \I1.N_174_adt_net_108976_\, Y => \I1.N_174\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2197\ : AO21
      port map(A => REGl130r, B => \I3.N_2058\, C => 
        \I3.VDBi_57l13r_adt_net_140578_\, Y => 
        \I3.VDBi_57l13r_adt_net_140592_\);
    
    \I1.REG_1_74\ : MUX2H
      port map(A => \REGl173r\, B => \I1.REG_74l173r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\, Y => 
        \I1.REG_1_74_net_1\);
    
    \I1.REG_74_i_o2_1_0tt_364_m2_e\ : NOR3
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__net_1\, 
        B => \PULSEl0r_adt_net_854536__net_1\, C => 
        \I1.PAGECNTL7R_526\, Y => 
        \I1.REG_74_i_o2_1_0tt_364_m2_e_net_1\);
    
    \I3.STATE1_ILLEGAL_2126\ : AND2
      port map(A => \I3.STATE1l10r_net_1\, B => 
        \I3.STATE1_IPL8R_10\, Y => \I3.N_1193_ip_adt_net_136530_\);
    
    \I3.STATE1_ILLEGAL_2131\ : AO21
      port map(A => \I3.STATE1_ipl5r\, B => 
        \I3.N_1180_adt_net_1502__net_1\, C => 
        \I3.N_1193_ip_adt_net_136553_\, Y => 
        \I3.N_1193_ip_adt_net_136554_\);
    
    \I2.DT_TEMP_770\ : MUX2H
      port map(A => \I2.DT_TEMPl9r_net_1\, B => 
        \I2.DT_TEMP_7l9r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_770_net_1\);
    
    \I2.FID_7_0_IVL15R_961\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl15r_net_1\, 
        Y => \I2.FID_7l15r_adt_net_17893_\);
    
    \I2.DT_SRAMl7r\ : MUX2L
      port map(A => \I2.N_875\, B => \I2.PIPE2_DTl7r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl7r_net_1\);
    
    \I3.UN7_RONLY_0_A2_0_A2_2637\ : NOR3
      port map(A => \I3.VAS_i_0_il13r\, B => \I3.VASl11r_net_1\, 
        C => \I3.VASl9r_net_1\, Y => \I3.N_544_adt_net_165558_\);
    
    \I2.OFFSET_37_1l5r\ : MUX2L
      port map(A => \REGl354r\, B => \REGl290r\, S => 
        \I2.PIPE7_DTL27R_65\, Y => \I2.N_640\);
    
    \I1.REG_74_0_ivl261r\ : AO21
      port map(A => \REGl261r\, B => 
        \I1.N_137_adt_net_854764__net_1\, C => 
        \I1.REG_74l261r_adt_net_124629_\, Y => \I1.REG_74l261r\);
    
    \I1.REG_1_127\ : MUX2H
      port map(A => \REGl226r\, B => \I1.REG_74l226r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\, Y => 
        \I1.REG_1_127_net_1\);
    
    RAMAD_padl0r : OB33PH
      port map(PAD => RAMAD(0), A => RAMAD_cl0r);
    
    \I3.VDBOFFB_30_IV_0L6R_2378\ : AO21
      port map(A => \REGl387r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l6r_adt_net_161954_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161983_\);
    
    \I3.VDBm_0l26r\ : MUX2L
      port map(A => \I3.PIPEAl26r_net_1\, B => 
        \I3.PIPEBl26r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_168\);
    
    \I2.SUB9_1_ADD_18x18_fast_I141_Y\ : XOR2
      port map(A => \I2.N225\, B => \I2.ADD_18x18_fast_I141_Y_0\, 
        Y => \I2.SUB9_1l4r\);
    
    \I3.VDBOFFB_30_IV_0L4R_2406\ : AND2
      port map(A => \REGl361r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        Y => \I3.VDBoffb_30l4r_adt_net_162330_\);
    
    \I2.PIPE6_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_470_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl16r_net_1\);
    
    TDCDB_padl26r : IB33
      port map(PAD => TDCDB(26), Y => TDCDB_cl26r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I67_Y\ : AND2
      port map(A => \I2.N249_0\, B => \I2.N252_0\, Y => \I2.N317\);
    
    \I2.ADE_4l11r\ : MUX2L
      port map(A => \I2.ROFFSETl12r_net_1\, B => \I2.WOFFSETl12r\, 
        S => NOESRAME_C_243, Y => \I2.ADE_4l11r_net_1\);
    
    \I3.PIPEA1_320\ : MUX2L
      port map(A => \I3.PIPEA1l22r_net_1\, B => 
        \I3.PIPEA1_12l22r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__251\, Y => 
        \I3.PIPEA1_320_net_1\);
    
    \I2.LEAD_FLAG6_643\ : AO21
      port map(A => \I2.N_4529_adt_net_1136__net_1\, B => 
        \I2.N_4529_adt_net_63916_\, C => 
        \I2.LEAD_FLAG6_643_adt_net_63956_\, Y => 
        \I2.LEAD_FLAG6_643_net_1\);
    
    \I5.AIR_WDATAl1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_56_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl1r_net_1\);
    
    \I2.TDCDBSl6r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl6r, Q => 
        \I2.TDCDBSl6r_net_1\);
    
    \I2.PIPE10_DT_17_i_0l16r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855596__net_1\, B => 
        \I2.PIPE9_DTl16r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l16r_net_1\);
    
    VDB_padl24r : IOB33PH
      port map(PAD => VDB(24), A => \I3.VDBml24r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl24r);
    
    \I2.MIC_REG3l6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_323_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l6r_net_1\);
    
    \I2.CHAINA_ERRF1\ : DFFC
      port map(CLK => CLK_c, D => \I2.CHAINA_ERRF1_492_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.CHAINA_ERRF1_net_1\);
    
    \I2.LEAD_FLAG6_7_i_0l6r\ : AOI21
      port map(A => \I2.N_215\, B => \I2.N_484\, C => \I2.N_222\, 
        Y => \I2.N_4529_adt_net_63916_\);
    
    \I2.N_4245_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4245\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4245_Rd1__net_1\);
    
    \I2.SUB8_520_2724\ : AND2FT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855156__net_1\, B
         => \I2.N_3560_i_net_1\, Y => 
        \I2.SUB8_520_adt_net_635605_\);
    
    \I2.DTE_1_868\ : MUX2L
      port map(A => \I2.DTE_1l30r_net_1\, B => 
        \I2.DTE_21_1_0_ivl30r_net_1\, S => \I2.N_2868_1\, Y => 
        \I2.DTE_1_868_net_1\);
    
    \I2.NPRSFIF_328\ : OR3
      port map(A => \I2.STATE3l5r_net_1\, B => 
        \I2.STATE3_i_il10r\, C => \I2.NPRSFIF_328_adt_net_97261_\, 
        Y => \I2.NPRSFIF_328_net_1\);
    
    \I2.STATE5_ns_i_0_a5_1l0r\ : AOI21FTF
      port map(A => COM_SERS, B => \I2.CHAIN_ERRS_net_1\, C => 
        \I2.MSERCLKS_net_1\, Y => \I2.N_4338_1\);
    
    \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_1_RD1__2941\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_1_RD1__458\);
    
    \I1.SSTATE_NS_I_0_A4_0_1_0L0R_1762\ : NOR2
      port map(A => \I1.sstatel10r_net_1\, B => 
        \I1.sstatel5r_net_1\, Y => 
        \I1.sstate_ns_i_0_a4_0_1l0r_adt_net_107171_\);
    
    \I2.PIPE1_DT_42_1_IVL10R_1461\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        B => \I2.PIPE1_DT_12l10r_net_1\, Y => 
        \I2.PIPE1_DT_42l10r_adt_net_49936_\);
    
    \I1.REG_74_0_IVL339R_1877\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l339r_adt_net_117314_\);
    
    \I1.REG_74_0_ivl346r\ : AO21
      port map(A => \REGl346r\, B => \I1.N_217\, C => 
        \I1.REG_74l346r_adt_net_116498_\, Y => \I1.REG_74l346r\);
    
    \I1.REG_74_0_ivl232r\ : AO21
      port map(A => \REGl232r\, B => \I1.N_105\, C => 
        \I1.REG_74l232r_adt_net_127452_\, Y => \I1.REG_74l232r\);
    
    \I3.VDBi_57l2r_adt_net_145305_\ : AO21
      port map(A => \I3.N_2045\, B => \I3.REGl93r\, C => 
        \I3.VDBi_57l2r_adt_net_145304__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145305__net_1\);
    
    \I3.STATE1_ns_1_iv_0l5r\ : OR2
      port map(A => \I3.STATE1_nsl5r_adt_net_136318_\, B => 
        \I3.STATE1_nsl5r_adt_net_136320_\, Y => \I3.STATE1_nsl5r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I2_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L2R_767\, B => \I2.PIPE4_DTL2R_859\, 
        Y => \I2.N_52\);
    
    \I2.RAMDT4L5R_3064\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_818\);
    
    \I1.REG_74_12L268R_1945\ : OR2
      port map(A => \I1.N_145_12_adt_net_123179_\, B => 
        \I1.REG_74_3_4_il380r\, Y => 
        \I1.N_145_12_adt_net_123140_\);
    
    \I3.REG_1l79r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_180_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl79r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I215_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl19r\, B => 
        \I2.PIPE7_DTl19r_net_1\, Y => 
        \I2.SUB_21x21_fast_I215_Y_0\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855396_\ : BFR
      port map(A => \I1.N_50_0_adt_net_1409__net_1\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\);
    
    \I2.DTE_2_1l6r\ : XOR2
      port map(A => \I2.CRC32l26r_net_1\, B => 
        \I2.DTE_2_1_0l6r_net_1\, Y => \I2.DTE_2_1l6r_net_1\);
    
    \I1.REG_1_87\ : MUX2H
      port map(A => \REGl186r\, B => \I1.REG_74l186r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, Y => 
        \I1.REG_1_87_net_1\);
    
    \I2.DTE_1l27r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l27r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l27r_Rd1__net_1\);
    
    \I2.OFFSET_37_27l2r\ : MUX2L
      port map(A => \I2.N_837\, B => \I2.N_821\, S => 
        \I2.PIPE7_DTL25R_687\, Y => \I2.N_845\);
    
    \I3.PIPEA_8l22r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854460__net_1\, B => 
        \I3.N_231\, Y => \I3.PIPEA_8l22r_net_1\);
    
    \I2.DT_TEMPl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_764_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl3r_net_1\);
    
    \I1.PAGECNT_321\ : MUX2H
      port map(A => \I1.PAGECNTl6r_adt_net_854928__net_1\, B => 
        \I1.N_1377\, S => \I1.PAGECNTe_adt_net_854892__net_1\, Y
         => \I1.PAGECNT_321_net_1\);
    
    \I2.DTESl12r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl12r, Q => 
        \I2.DTESl12r_net_1\);
    
    \I1.REG_74l396r\ : AO21FTF
      port map(A => 
        \I1.REG_74_1_396_m7_i_3_adt_net_854840__net_1\, B => 
        \I1.N_265_adt_net_110486_\, C => \I1.REG_74_13_388_N_11\, 
        Y => \I1.N_265\);
    
    \I3.un7_ronly_0_a2_0_a2\ : AND3FFT
      port map(A => \I3.VAS_i_0_il14r\, B => \I3.VAS_i_0_il10r\, 
        C => \I3.N_544_adt_net_165558_\, Y => \I3.N_544\);
    
    \I2.SUB8l7r_1597\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_510_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8L7R_704\);
    
    \I2.DT_TEMP_7l28r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854232__net_1\, B => 
        \I2.DT_SRAMl28r_net_1\, Y => \I2.DT_TEMP_7l28r_net_1\);
    
    \I2.STATEel4r\ : DFFS
      port map(CLK => CLK_c, D => \I2.STATEe_nsl0r_net_1\, SET
         => \I2.STATEe_i_0l0r_net_1\, Q => \I2.STATEel4r_net_1\);
    
    \I2.BNCID_VECTROR_9_TZ_1419\ : AO21
      port map(A => \I2.BNCID_VECTra13_1_net_1\, B => 
        \I2.BNCID_VECTro_13\, C => 
        \I2.BNCID_VECTror_9_tz_adt_net_48087_\, Y => 
        \I2.BNCID_VECTror_9_tz_adt_net_48098_\);
    
    \I1.REG_74_0_IVL399R_1790\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_30_sqmuxa_adt_net_854372__net_1\, Y => 
        \I1.REG_74l399r_adt_net_110186_\);
    
    \I3.VDBi_23l1r_adt_net_145530_\ : AND3FFT
      port map(A => TRM_BUSY_c, B => \I3.REGMAPl3r_net_1\, C => 
        \I3.N_2040_261\, Y => 
        \I3.VDBi_23l1r_adt_net_145530__net_1\);
    
    \I2.PIPE6_DT_0_SQMUXA_I_O4_1594\ : AND2
      port map(A => \I2.N_217\, B => \I2.N_4542\, Y => 
        \I2.N_4551_adt_net_63747_\);
    
    \I2.CRC32_12_il29r\ : NOR2
      port map(A => \I2.N_2867_1_adt_net_854964__net_1\, B => 
        \I2.N_18_i_0_i_0\, Y => \I2.N_3946\);
    
    \I2.DTO_16_1_ivl15r\ : OR2
      port map(A => \I2.DTO_16_1l15r_adt_net_31963_\, B => 
        \I2.DTO_16_1l15r_adt_net_31964_\, Y => \I2.DTO_16_1l15r\);
    
    \I1.REG_74_0_IVL283R_1936\ : NOR2FT
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l283r_adt_net_122463_\);
    
    REGl303r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_204_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl303r\);
    
    \I1.NCS0_56_2071\ : AND2
      port map(A => \I1.NCS0_net_1\, B => \I1.N_436_i_i\, Y => 
        \I1.NCS0_56_adt_net_133847_\);
    
    \I3.VDBI_57_IV_0_0L0R_2287\ : AO21
      port map(A => \I3.PIPEAl0r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l0r_adt_net_146651_\, Y => 
        \I3.VDBi_57l0r_adt_net_146660_\);
    
    \I2.STATE2l4r_adt_net_855676_\ : BFR
      port map(A => \I2.STATE2l4r_adt_net_855684__net_1\, Y => 
        \I2.STATE2l4r_adt_net_855676__net_1\);
    
    \I3.REG_0_sqmuxa_1_0_o2_i_a3\ : AND2
      port map(A => \I3.REGMAPl9r_adt_net_854332__net_1\, B => 
        \I3.N_1906_i_0_0\, Y => \I3.N_1935\);
    
    \I3.VDBOFFB_30_IV_0L6R_2379\ : AO21
      port map(A => \REGl331r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l6r_adt_net_161958_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161984_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I102_Y\ : NAND2
      port map(A => \I2.N313_1\, B => \I2.N317\, Y => \I2.N356\);
    
    \I3.VDBOFFB_30_IV_0L2R_2440\ : AND2
      port map(A => \REGl375r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162702_\);
    
    \I1.REG_18_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_267\, B => \I1.N_242\, Y => 
        \I1.REG_18_sqmuxa\);
    
    \I5.REG_1l423r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_36_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl423r);
    
    \I2.WPAGEL12R_2998\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_951_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEL12R_752\);
    
    \I2.CRC32_7l1r\ : XOR2FT
      port map(A => \I2.CRC32l1r_net_1\, B => 
        \I2.DT_TEMPl1r_net_1\, Y => \I2.CRC32_7_il1r\);
    
    \I2.resyn_0_I2_TRAIL_MIS6_1_sqmuxa_0_a4_i\ : NOR2
      port map(A => \I2.N_4524\, B => \I2.PIPE4_DTl30r_net_1\, Y
         => \I2.N_4643\);
    
    \I2.OFFSET_37_1l3r\ : MUX2L
      port map(A => \REGl352r\, B => \REGl288r\, S => 
        \I2.PIPE7_DTL27R_65\, Y => \I2.N_638\);
    
    \I2.REG_1l32r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n0_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl32r);
    
    \I1.REG_74L220R_2013\ : OR3FFT
      port map(A => \I1.N_1366\, B => 
        \I1.REG_74_12_220_m9_i_net_1\, C => 
        \I1.N_89_adt_net_128733_\, Y => \I1.N_89_adt_net_128736_\);
    
    \I2.PIPE8_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_553_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl25r_net_1\);
    
    \I3.PIPEB_84_2339\ : NOR2FT
      port map(A => \I3.PIPEBl5r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_84_adt_net_160503_\);
    
    \I2.TDCDBSl0r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl0r, Q => 
        \I2.TDCDBSl0r_net_1\);
    
    \I2.un7_bnc_id_1_I_9\ : XOR2
      port map(A => \I2.N_45\, B => \I2.BNC_IDl2r_net_1\, Y => 
        \I2.I_9_1\);
    
    \I1.REG_74_0_ivl376r\ : AO21
      port map(A => \REGl376r\, B => \I1.N_249\, C => 
        \I1.REG_74l376r_adt_net_112829_\, Y => \I1.REG_74l376r\);
    
    \I2.MIC_REG2_311\ : MUX2H
      port map(A => \I2.MIC_REG2l2r_net_1\, B => 
        \I2.MIC_REG2l3r_adt_net_834020_Rd1__net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG2_311_net_1\);
    
    \I2.SRAM_EVNT_n0_0\ : XOR2
      port map(A => \I2.SRAM_EVNTl0r_net_1\, B => \I2.N_132\, Y
         => \I2.SRAM_EVNT_n0_0_net_1\);
    
    \I1.REG_1_123\ : MUX2H
      port map(A => \REGl222r\, B => \I1.REG_74l222r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_123_net_1\);
    
    \I3.TCNT3_n1\ : XOR2
      port map(A => \I3.TCNT3_i_0_il0r_net_1\, B => 
        \I3.TCNT3l1r_net_1\, Y => \I3.TCNT3_n1_net_1\);
    
    SP2_pad : OB33PH
      port map(PAD => SP2, A => \GND\);
    
    \I2.DTESl7r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl7r, Q => 
        \I2.DTESl7r_net_1\);
    
    \I2.PIPE7_DTL26R_2894\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_348\);
    
    \I3.PIPEA_239\ : MUX2L
      port map(A => \I3.PIPEAl8r_net_1\, B => 
        \I3.PIPEA_8l8r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854672__net_1\, Y
         => \I3.PIPEA_239_net_1\);
    
    \I1.REG_74_0_iv_i_a2l209r\ : AO21
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, C => 
        \I1.N_1348_adt_net_129759_\, Y => \I1.N_1348\);
    
    \I2.MIC_REG3L2R_2945\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_319_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3L2R_462\);
    
    \I2.DTO_16_1_IV_0_0L26R_1085\ : AO21
      port map(A => \I2.N_197_150\, B => \I2.DT_SRAMl26r_net_1\, 
        C => \I2.DTO_16_1l26r_adt_net_29428_\, Y => 
        \I2.DTO_16_1l26r_adt_net_29438_\);
    
    \I3.REG_1_275\ : MUX2H
      port map(A => VDB_inl3r, B => \I3.REGl94r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_275_0\);
    
    \I3.REG_1l53r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_154_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl53r);
    
    \I2.LSRAM_INl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_394_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl10r_net_1\);
    
    \I3.PIPEA1_12l12r\ : AND2
      port map(A => DPR_cl12r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854504__net_1\, Y => 
        \I3.PIPEA1_12l12r_net_1\);
    
    \I2.DT_TEMP_7l22r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854236__net_1\, B => 
        \I2.DT_SRAMl22r_net_1\, Y => \I2.DT_TEMP_7l22r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I66_Y\ : AO21
      port map(A => \I2.N300\, B => \I2.N303\, C => \I2.N299\, Y
         => \I2.N334\);
    
    \I2.DT_TEMP_764\ : MUX2H
      port map(A => \I2.DT_TEMPl3r_net_1\, B => 
        \I2.DT_TEMP_7l3r_net_1\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.DT_TEMP_764_net_1\);
    
    \I2.DTO_16_1_IV_0_0L19R_1122\ : AND2
      port map(A => \I2.N_4671_adt_net_854592__net_1\, B => 
        \I2.DT_TEMPl19r_net_1\, Y => 
        \I2.DTO_16_1l19r_adt_net_30968_\);
    
    \I3.un41_reg_ads_0_a2_3_a3_2\ : NAND3FFT
      port map(A => \I3.LWORDS_net_1\, B => \I3.N_553\, C => 
        \I3.N_545\, Y => \I3.un41_reg_ads_2\);
    
    \I2.PIPE10_DT_606\ : MUX2L
      port map(A => \I2.PIPE10_DTl1r_net_1\, B => 
        \I2.PIPE9_DTl1r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_606_net_1\);
    
    \I2.REG_0L3R_ADT_NET_19773_RD1__3102\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.REG_0l3r_adt_net_19773_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.REG_0L3R_ADT_NET_19773_RD1__888\);
    
    \I3.PIPEB_87\ : AO21
      port map(A => DPR_cl8r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_87_adt_net_160377_\, Y => 
        \I3.PIPEB_87_net_1\);
    
    \I2.LSRAM_IN_398\ : MUX2L
      port map(A => \I2.PIPE5_DTl14r_net_1\, B => 
        \I2.LSRAM_INl14r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_398_net_1\);
    
    \I2.PIPE7_DTL27R_2788\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_81\);
    
    \I3.REGMAPl14r_1626\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un57_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL14R_733\);
    
    \I1.REG_74_0_iv_i_a2l197r\ : AO21
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_129_adt_net_130791_\, Y => \I1.N_129\);
    
    \I3.PIPEB_96_2327\ : NOR2FT
      port map(A => \I3.PIPEBl17r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_96_adt_net_159999_\);
    
    \I1.N_1169_adt_net_854820_\ : BFR
      port map(A => \I1.N_1169_adt_net_854824__net_1\, Y => 
        \I1.N_1169_adt_net_854820__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I3_P0N\ : OR2
      port map(A => \I2.N_3539_i_i\, B => \I2.G_1_2\, Y => 
        \I2.N235\);
    
    VAD_padl10r : IOB33PH
      port map(PAD => VAD(10), A => \I3.VADml10r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl10r);
    
    REGl239r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_140_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl239r\);
    
    \I2.OFFSET_37_5l6r\ : MUX2L
      port map(A => \REGl403r\, B => \REGl339r\, S => 
        \I2.PIPE7_DTL27R_76\, Y => \I2.N_673\);
    
    \I1.REG_74_0_ivl299r\ : AO21
      port map(A => \REGl299r\, B => \I1.N_169\, C => 
        \I1.REG_74l299r_adt_net_120954_\, Y => \I1.REG_74l299r\);
    
    \I2.OFFSET_37_27l5r\ : MUX2L
      port map(A => \I2.N_840\, B => \I2.N_824\, S => 
        \I2.PIPE7_DTL25R_687\, Y => \I2.N_848\);
    
    \I2.MIC_ERR_REGS_351\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl23r_net_1\, B => 
        \I2.MIC_ERR_REGSl22r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_351_net_1\);
    
    \I2.MIC_ERR_REGS_359\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl31r_net_1\, B => 
        \I2.MIC_ERR_REGSl30r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_359_net_1\);
    
    \I2.FID_7_ivl4r\ : OR2
      port map(A => \I2.FID_7l4r_adt_net_93158_\, B => 
        \I2.FID_7l4r_adt_net_93159_\, Y => \I2.FID_7l4r\);
    
    \I2.CRC32_825\ : MUX2L
      port map(A => \I2.CRC32l30r_net_1\, B => \I2.N_3947\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_825_net_1\);
    
    \I1.REG_74_7_i_a2_a0_0_1l404r\ : NOR2
      port map(A => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__19\, 
        B => \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_1_RD1__458\, Y => 
        \I1.N_232_1\);
    
    \I3.PULSEl5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_335_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl5r);
    
    \I1.REG_1_126\ : MUX2H
      port map(A => \REGl225r\, B => \I1.REG_74l225r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\, Y => 
        \I1.REG_1_126_net_1\);
    
    \I2.PIPE4_DTL8R_2966\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL8R_483\);
    
    \I2.LSRAM_RADDRl1r\ : MUX2L
      port map(A => \LSRAM_FL_RADDRl1r\, B => 
        \I2.LSRAM_RADDRil1r_net_1\, S => FLUSH, Y => 
        \I2.LSRAM_RADDRl1r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I110_Y_0\ : AND2FT
      port map(A => \I2.N_3560_i_net_1\, B => 
        \I2.ADD_18x18_fast_I110_Y_0_adt_net_3684__net_1\, Y => 
        \I2.ADD_18x18_fast_I110_Y_0\);
    
    \I2.SRAM_EVNT_c0_i\ : OA21FTF
      port map(A => \I2.N_128_1\, B => \I2.N_132\, C => 
        \I2.SRAM_EVNTl0r_net_1\, Y => \I2.N_3825\);
    
    \I3.MYBERRi\ : DFFS
      port map(CLK => CLK_c, D => \I3.MYBERRi_62_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => MYBERR_c);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I32_P0N_1760\ : OR2FT
      port map(A => \I2.LSRAM_OUTl11r\, B => 
        \I2.PIPE7_DTL11R_694\, Y => \I2.N264_0_867\);
    
    \I2.RAMDT4L5R_3063\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_817\);
    
    \I2.DTO_16_1_IVL14R_1149\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854624__net_1\, 
        B => \I2.DT_TEMPl14r_net_1\, C => 
        \I2.DTO_16_1l14r_adt_net_32202_\, Y => 
        \I2.DTO_16_1l14r_adt_net_32208_\);
    
    \I3.PIPEA_8l16r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854468__net_1\, B => 
        \I3.N_225\, Y => \I3.PIPEA_8l16r_net_1\);
    
    \I2.PIPE5_DT_683\ : MUX2L
      port map(A => \I2.PIPE5_DTl7r_net_1\, B => 
        \I2.PIPE5_DT_6l7r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_683_net_1\);
    
    \I1.REG_1_182\ : MUX2H
      port map(A => \REGl281r\, B => \I1.REG_74l281r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\, Y => 
        \I1.REG_1_182_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2612\ : AO21
      port map(A => \REGl262r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        C => \I3.VDBoffa_31l1r_adt_net_164424_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164453_\);
    
    \I2.CRC32_12_IL9R_1349\ : OA21FTF
      port map(A => 
        \I2.N_4667_1_adt_net_1046__adt_net_854424__net_1\, B => 
        \I2.N_57_i_0\, C => \I2.N_2867_1_adt_net_854960__net_1\, 
        Y => \I2.N_3926_adt_net_42578_\);
    
    \I2.PIPE7_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl13r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl13r_net_1\);
    
    REGl172r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_73_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl172r\);
    
    \I1.REG_1_241\ : MUX2H
      port map(A => \REGl340r\, B => \I1.REG_74l340r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\, Y
         => \I1.REG_1_241_net_1\);
    
    \I2.STATE1_ns_o2_0l0r\ : AND2
      port map(A => \I2.N_3287_i_0\, B => \I2.N_3358\, Y => 
        \I2.STATE1_ns_o2_0l0r_net_1\);
    
    \I1.REG_1_sqmuxa_0_a2_0\ : OR3
      port map(A => \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__363\, B
         => \I1.PAGECNTL8R_457\, C => \I1.N_1169_168\, Y => 
        \I1.N_242\);
    
    \I3.REGMAPl10r_1612\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un44_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL10R_719\);
    
    \I3.REG_44_i_a2_0l85r\ : NOR2
      port map(A => VDB_inl2r, B => \I3.N_98\, Y => \I3.N_1665\);
    
    DPR_padl29r : IB33
      port map(PAD => DPR(29), Y => DPR_cl29r);
    
    \I3.un47_reg_ads_0_a2_0_a2\ : OR2FT
      port map(A => \I3.WRITES_8\, B => \I3.N_546_373\, Y => 
        \I3.N_547\);
    
    ADO_padl5r : OB33PH
      port map(PAD => ADO(5), A => ADO_cl5r);
    
    \I5.REG_1_31\ : MUX2L
      port map(A => REGl131r, B => REGl418r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_31_net_1\);
    
    \I5.sstate1l0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1se_12_i_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.sstate1l0r_net_1\);
    
    \I2.EVNT_WORD_713\ : AO21FTT
      port map(A => \I2.N_2864_0_adt_net_854268__net_1\, B => 
        \I2.EVNT_WORDl0r_net_1\, C => 
        \I2.EVNT_WORD_713_adt_net_53148_\, Y => 
        \I2.EVNT_WORD_713_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I137_Y_I_1576\ : OAI21
      port map(A => \I2.PIPE4_DTL12R_858\, B => 
        \I2.PIPE4_DTL13R_642\, C => \I2.RAMDT4L12R_146\, Y => 
        \I2.N_40_0_adt_net_58199_\);
    
    DTE_padl18r : IOB33PH
      port map(PAD => DTE(18), A => \I2.DTE_1l18r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl18r);
    
    \I2.PIPE1_DT_42_1_ivl8r\ : OR3
      port map(A => \I2.PIPE1_DT_42l8r_adt_net_50436_\, B => 
        \I2.PIPE1_DT_42l8r_adt_net_50445_\, C => 
        \I2.PIPE1_DT_42l8r_adt_net_50446_\, Y => 
        \I2.PIPE1_DT_42l8r\);
    
    \I3.un60_reg_ads_0_a2_0_a2\ : OR2
      port map(A => \I3.N_546\, B => \I3.N_554\, Y => \I3.N_632\);
    
    \I2.STATE3_NS_O3L10R_1043\ : NAND2
      port map(A => \I2.DTOSl30r_net_1\, B => \I2.DTOSl28r_net_1\, 
        Y => \I2.N_3016_adt_net_24530_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I62_Y\ : AO21
      port map(A => \I2.N299\, B => \I2.N296\, C => \I2.N295\, Y
         => \I2.N330\);
    
    \I2.EVNT_NUM_n8_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl8r_net_1\, B => 
        \I2.EVNT_NUM_c7_net_1\, Y => \I2.EVNT_NUM_n8_tz_i\);
    
    \I1.PAGECNT_0l8r_adt_net_834720_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_319_adt_net_854860__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__net_1\);
    
    \I2.dataout_0_adt_net_855804_\ : BFR
      port map(A => \I2.dataout_0\, Y => 
        \I2.dataout_0_adt_net_855804__net_1\);
    
    \I1.REG_74_0_IV_I_A2L202R_2032\ : AND2
      port map(A => \REGl202r\, B => \I1.N_182_i\, Y => 
        \I1.N_1341_adt_net_130361_\);
    
    \I1.REG_74_0_IV_0L364R_1843\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.REG_25_sqmuxa\, 
        Y => \I1.REG_74l364r_adt_net_114525_\);
    
    \I3.VDBOFFA_31_IV_0L2R_2590\ : AO21
      port map(A => \REGl191r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.VDBoffa_31l2r_adt_net_164218_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164259_\);
    
    REGl331r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_232_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl331r\);
    
    \I3.EVREAD_DS\ : DFFC
      port map(CLK => CLK_c, D => \I3.EVREAD_DS_124_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I3.EVREAD_DS_net_1\);
    
    REGl312r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_213_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl312r\);
    
    \I3.UN224_REG_ADS_0_A2_3_A2_2_2646\ : NOR2
      port map(A => \I3.VAS_I_0_IL15R_346\, B => \I3.VASL8R_347\, 
        Y => \I3.N_545_adt_net_165680_\);
    
    NOEDTK_pad : OB33PH
      port map(PAD => NOEDTK, A => NOEDTK_C_14);
    
    \I2.STATE2_ns_i_0_1l0r\ : OR3
      port map(A => \I2.STATE2l2r_adt_net_855212__net_1\, B => 
        \I2.STATE2_ns_i_0_1_il0r_adt_net_21493_\, C => 
        \I2.STATE2l1r_adt_net_855116__net_1\, Y => 
        \I2.STATE2_ns_i_0_1_il0r\);
    
    \I2.TDCDASl27r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl27r, Q => 
        \I2.TDCDASl27r_net_1\);
    
    \I2.DTO_9_IV_0L20R_1116\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl20r_net_1\, C => 
        \I2.DTO_9l20r_adt_net_30718_\, Y => 
        \I2.DTO_9l20r_adt_net_30726_\);
    
    \I2.TDCGDA1\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => TDCGDA_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.TDCGDA1_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I144_Y_2658\ : AO21
      port map(A => \I2.N510_adt_net_220872_\, B => 
        \I2.N510_adt_net_220925_\, C => \I2.N510_adt_net_232425_\, 
        Y => \I2.N510\);
    
    \I2.PIPE9_DT_283\ : MUX2L
      port map(A => \I2.PIPE9_DTl14r_net_1\, B => 
        \I2.PIPE8_DTl14r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_283_net_1\);
    
    \I2.DT_TEMP_767\ : MUX2H
      port map(A => \I2.DT_TEMPl6r_net_1\, B => 
        \I2.DT_TEMP_7l6r_net_1\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.DT_TEMP_767_net_1\);
    
    \I3.PIPEA_258\ : MUX2L
      port map(A => \I3.PIPEAl27r_net_1\, B => 
        \I3.PIPEA_8l27r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854656__net_1\, Y
         => \I3.PIPEA_258_net_1\);
    
    \I2.TRGSERVL0R_2950\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.DWACT_ADD_CI_0_partial_sum_1l0r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGSERVL0R_467\);
    
    \I2.L2SERVl3r_1259\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_521\);
    
    \I2.EVNT_NUM_n7_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl7r_net_1\, B => 
        \I2.EVNT_NUM_c6_net_1\, Y => \I2.EVNT_NUM_n7_tz_i\);
    
    \I2.L2TYPE_4_IL4R_1635\ : AND2
      port map(A => \I2.L2TYPEl4r_net_1\, B => 
        \I2.N_4448_adt_net_68212_\, Y => 
        \I2.N_4448_adt_net_68255_\);
    
    \I3.REG_1_178\ : MUX2L
      port map(A => VDB_inl29r, B => REGl77r, S => 
        \I3.N_1935_adt_net_855316__net_1\, Y => \I3.REG_1_178_0\);
    
    \I3.REG_44_il86r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_1632_adt_net_150363_\, Y => \I3.N_1632\);
    
    \I3.PIPEBl14r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_93_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl14r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL15R_1433\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl47r_net_1\, C => 
        \I2.PIPE1_DT_42l15r_adt_net_48697_\, Y => 
        \I2.PIPE1_DT_42l15r_adt_net_48715_\);
    
    \I2.EVNT_NUM_n3_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl3r_net_1\, B => 
        \I2.EVNT_NUM_c2_net_1\, Y => \I2.EVNT_NUM_n3_tz_i\);
    
    \I2.L2TYPEl5r_1552\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_594_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_I_0_IL5R_659\);
    
    \I2.INT_ERRAF1\ : DFFC
      port map(CLK => CLK_c, D => \I2.INT_ERRAF1_494_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.INT_ERRAF1_net_1\);
    
    \I5.SCL_1_i_o4\ : NAND3FFT
      port map(A => \I5.sstate1l13r_net_1\, B => 
        \I5.sstate1l0r_net_1\, C => \I5.SDAnoe_8_adt_net_9736_\, 
        Y => \I5.N_82\);
    
    \I2.END_TDC1_1_SQMUXA_I_O2_1013\ : NOR3FTT
      port map(A => \I2.N_3887_adt_net_21862_\, B => 
        \I2.un6_tdcgdb1_3_net_1\, C => \I2.un6_tdcgdb1_2_net_1\, 
        Y => \I2.N_3887_adt_net_21857_\);
    
    REGl279r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_180_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl279r\);
    
    \I1.REG_1_141\ : MUX2H
      port map(A => \REGl240r\, B => \I1.REG_74l240r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\, Y => 
        \I1.REG_1_141_net_1\);
    
    \I4.un2_end_tdc_1\ : OR3
      port map(A => LEAD_FLAGl7r, B => LEAD_FLAGl6r, C => 
        \I4.un2_end_tdc_1_adt_net_15219_\, Y => 
        \I4.un2_end_tdc_1_net_1\);
    
    \I3.VDBi_40_1l11r\ : MUX2L
      port map(A => REGl128r, B => \I3.VDBi_31l11r_net_1\, S => 
        \I3.REGMAPl16r_net_1\, Y => \I3.N_349\);
    
    \I2.EVNT_NUM_953\ : MUX2L
      port map(A => \I2.EVNT_NUMl10r_net_1\, B => 
        \I2.EVNT_NUM_n10_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_953_net_1\);
    
    \I3.VDBoffa_47\ : OR3
      port map(A => \I3.VDBoffa_47_adt_net_164118_\, B => 
        \I3.VDBoffa_31l3r_adt_net_164079_\, C => 
        \I3.VDBoffa_31l3r_adt_net_164080_\, Y => 
        \I3.VDBoffa_47_net_1\);
    
    \I3.REG2_15_0_a2_0_a3l405r\ : AND3
      port map(A => VDB_inl0r, B => \I3.REGMAPl50r_net_1\, C => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        Y => \I3.REG2_15l405r\);
    
    \I1.REG_74_0_ivl326r\ : AO21
      port map(A => \REGl326r\, B => \I1.N_201\, C => 
        \I1.REG_74l326r_adt_net_118432_\, Y => \I1.REG_74l326r\);
    
    \I2.DTO_16_1_iv_0_o2_0_i_o2l21r_772\ : OAI21FTF
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.N_182_ADT_NET_1007__155\, Y => \I2.N_197_150\);
    
    \I2.PIPE10_DT_17_i_a3_0l13r\ : AND2
      port map(A => \I2.N_22_i_0\, B => \I2.SUB9l20r_net_1\, Y
         => \I2.N_26\);
    
    \I2.FID_7_0_IVL23R_990\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl71r, C => 
        \I2.FID_7l23r_adt_net_19209_\, Y => 
        \I2.FID_7l23r_adt_net_19217_\);
    
    \I2.DTO_cl_64_il31r\ : AOI21FTF
      port map(A => \I2.DTO_cll31r\, B => 
        \I2.un1_DTO_cl_0_sqmuxa\, C => \I2.WROi_10_1\, Y => 
        \I2.DTO_cl_64_il31r_net_1\);
    
    REGl330r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_231_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl330r\);
    
    \I2.ROFFSET_n10_tz\ : XOR2FT
      port map(A => \I2.ROFFSETl10r_net_1\, B => 
        \I2.ROFFSET_c9_net_1\, Y => \I2.ROFFSET_n10_tz_i\);
    
    \I3.VDBoffb_30_iv_0l2r\ : AND2
      port map(A => \REGl367r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162694_\);
    
    \I3.un33_reg_ads_0_a2_0_a2\ : OR3FFT
      port map(A => \I3.VASl4r_net_1\, B => \I3.N_552\, C => 
        \I3.VASl2r_net_1\, Y => \I3.N_634\);
    
    \I2.SUB8_522_2705\ : NOR3FTT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855136__net_1\, B
         => \I2.SUB_21x21_fast_I215_Y_0\, C => 
        \I2.N477_adt_net_438351_\, Y => 
        \I2.SUB8_522_adt_net_552099_\);
    
    \I0.CLEAR_STATi_4\ : OR2
      port map(A => TDC_RES_c_c, B => CLEAR_STAT_12, Y => 
        \I0.CLEAR_STATi_4_net_1\);
    
    \I2.un1_tdc_res_37_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl417r, Y => 
        \I2.N_4618_i_0\);
    
    \I2.OFFSET_37_8l3r\ : MUX2L
      port map(A => \REGl360r\, B => \REGl296r\, S => 
        \I2.PIPE7_DTL27R_71\, Y => \I2.N_694\);
    
    \I3.PIPEA_232\ : MUX2L
      port map(A => \I3.PIPEAl1r_net_1\, B => 
        \I3.PIPEA_8l1r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854680__net_1\, Y
         => \I3.PIPEA_232_net_1\);
    
    \I2.DT_TEMP_7l16r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854244__net_1\, B => 
        \I2.DT_SRAMl16r_net_1\, Y => \I2.DT_TEMP_7l16r_net_1\);
    
    \I2.EVNT_NUMl3r_1490\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_960_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUML3R_597\);
    
    \I2.EVNT_WORD_714\ : MUX2H
      port map(A => \I2.EVNT_WORDl1r_net_1\, B => \I2.I_5_0\, S
         => \I2.N_2864_0_adt_net_854276__net_1\, Y => 
        \I2.EVNT_WORD_714_net_1\);
    
    \I1.BYTECNT_n3_0\ : OAI21
      port map(A => \I1.N_223_adt_net_854844__net_1\, B => 
        \I1.N_392_i\, C => \I1.N_485\, Y => \I1.BYTECNT_n3\);
    
    \I2.G_EVNT_NUM_n1_i\ : NOR3
      port map(A => EV_RES_C_568, B => \I2.N_279\, C => 
        \I2.N_186\, Y => \I2.N_4637\);
    
    \I2.DTO_1l21r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l21r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l21r_Rd1__net_1\);
    
    \I2.CHB_DATA8_2_i\ : OAI21FTF
      port map(A => \I2.CHB_DATA8_net_1\, B => \I2.N_4402\, C => 
        \I2.N_4397_adt_net_90034_\, Y => \I2.N_4397\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I151_Y_i_1\ : OR3FFT
      port map(A => \I2.N_41_0\, B => \I2.N_33_0\, C => 
        \I2.N_63_0\, Y => \I2.N_1_1_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I171_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l1r_net_1\, B => 
        \I2.PIPE4_DT_i_il1r_net_1\, Y => 
        \I2.ADD_21x21_fast_I171_Y_0\);
    
    \I5.AIR_WDATA_62\ : MUX2H
      port map(A => \I5.N_463\, B => \I5.AIR_WDATAl15r_net_1\, S
         => \I5.N_461\, Y => \I5.AIR_WDATA_62_net_1\);
    
    \I3.PIPEB_92\ : AO21
      port map(A => DPR_cl13r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_92_adt_net_160167_\, Y => 
        \I3.PIPEB_92_net_1\);
    
    \I3.VDBOFFA_31_IV_0L3R_2566\ : AND2
      port map(A => \REGl232r\, B => \I3.REGMAPl26r_net_1\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164032_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I141_Y_0_O4_2681\ : 
        AOI21FTT
      port map(A => \I2.N_95_0\, B => \I2.N_45_1_adt_net_271427_\, 
        C => \I2.N_16_0\, Y => \I2.N522_0_adt_net_384644_\);
    
    \I1.REG_74_0_iv_0l271r\ : AO21
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, C => 
        \I1.REG_74l271r_adt_net_123732_\, Y => \I1.REG_74l271r\);
    
    \I2.MAJORITY_REG_IL4R_1020\ : AOI21
      port map(A => \I2.MIC_REG2_i_0_il4r_net_1\, B => 
        \I2.MIC_REG1l4r_net_1\, C => \I2.MIC_REG3l4r_net_1\, Y
         => \I2.N_4424_adt_net_22594_\);
    
    \I3.RAMAD_VMEl12r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_36_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl12r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I177_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_800\, B => 
        \I2.PIPE4_DTl7r_adt_net_854552__adt_net_854948__net_1\, Y
         => \I2.ADD_21x21_fast_I177_Y_0_0\);
    
    \I2.resyn_0_I2_FID_444\ : MUX2H
      port map(A => FID_cl28r, B => \I2.FID_7l28r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\, 
        Y => \I2.FID_444\);
    
    \I2.PIPE6_DT_462\ : MUX2H
      port map(A => \I2.PIPE5_DTl8r_net_1\, B => 
        \I2.PIPE6_DTl8r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_462_net_1\);
    
    \I2.G_EVNT_NUM_n3_i_0_o2_1292\ : AND2FT
      port map(A => \I2.N_187\, B => \I2.G_EVNT_NUML3R_399\, Y
         => \I2.N_189_554\);
    
    \I2.un21_pipe5_dt_4\ : XOR2
      port map(A => \I2.un21_pipe5_dt_3_net_1\, B => 
        \I2.un21_pipe5_dt_2_net_1\, Y => 
        \I2.un21_pipe5_dt_4_net_1\);
    
    \I2.BNCID_VECTrff_14\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_14_251_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_14\);
    
    \I5.SDAnoe_8_0_o4\ : NAND2
      port map(A => \I5.SSTATE1L13R_571\, B => \I5.PULSE_FL_572\, 
        Y => \I5.N_64\);
    
    \I3.VDBi_10l8r\ : AND2FT
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__489\, B => 
        \I3.REGMAPl2r_net_1\, Y => \I3.VDBi_10l8r_net_1\);
    
    \I1.PAGECNT_325\ : MUX2H
      port map(A => \I1.PAGECNTl2r_adt_net_834908_Rd1__net_1\, B
         => \I1.PAGECNT_n2\, S => 
        \I1.PAGECNTe_adt_net_854896__net_1\, Y => 
        \I1.PAGECNT_325_net_1\);
    
    \I2.N_3496_adt_net_926_\ : OR2
      port map(A => \I2.STATEe_ipl2r\, B => \I2.STATEe_ipl3r\, Y
         => \I2.N_3496_adt_net_926__net_1\);
    
    \I3.TCNT1_c2\ : AND2
      port map(A => \I3.TCNT1l2r_net_1\, B => \I3.TCNT1_c1_net_1\, 
        Y => \I3.TCNT1_c2_net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2458\ : AND2
      port map(A => \REGl374r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162892_\);
    
    \I3.PIPEA1l18r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_316_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l18r_net_1\);
    
    \I1.REG_74_0_IV_0L225R_2002\ : AND2
      port map(A => \REGl225r\, B => \I1.N_97\, Y => 
        \I1.REG_74l225r_adt_net_128222_\);
    
    REGl371r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_272_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl371r\);
    
    \I1.REG_74_0_iv_i_a2l201r\ : AO21
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_1340_adt_net_130447_\, Y => \I1.N_1340\);
    
    \I2.DTE_1_873\ : MUX2L
      port map(A => \I2.DTE_1l18r_Rd1__net_1\, B => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835988_Rd1__net_1\, Y => 
        \I2.DTE_1l18r\);
    
    \I2.DT_SRAMl1r\ : MUX2L
      port map(A => \I2.N_869\, B => \I2.PIPE2_DTl1r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl1r_net_1\);
    
    \I2.DTO_9_IV_0L23R_1097\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        B => \I2.G_EVNT_NUMl7r_net_1\, Y => 
        \I2.DTO_9l23r_adt_net_30040_\);
    
    \I3.VDBOFFB_30_IV_0L0R_2482\ : AO21
      port map(A => \REGl317r\, B => \I3.REGMAPl37r_net_1\, C => 
        \I3.VDBoffb_30l0r_adt_net_163078_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163119_\);
    
    \I1.REG_74_22l404r\ : OR3FFT
      port map(A => \I1.REG_74_4_i_a2_404_N_4_i\, B => 
        \I1.N_347_adt_net_854788__net_1\, C => \I1.N_396_190\, Y
         => \I1.N_201_9\);
    
    \I3.VDBi_31l12r\ : MUX2L
      port map(A => \I3.REGl145r\, B => \I3.VDBi_20l12r\, S => 
        \I3.REGMAPl17r_adt_net_854288__net_1\, Y => 
        \I3.VDBi_31l12r_net_1\);
    
    \I2.PIPE1_DT_42_1_IV_2L27R_1365\ : OAI21TTF
      port map(A => REGl447r, B => 
        \I2.N_3234_adt_net_855652__net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46033_\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46038_\);
    
    \I2.MIC_REG3L3R_3050\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_320_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3L3R_804\);
    
    \I1.REG_74_0_IVL377R_1822\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l377r_adt_net_112743_\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_783\ : NOR3
      port map(A => \I2.N_4646_1_adt_net_19635__net_1\, B => 
        \I2.N_4646_1_ADT_NET_19637_RD1__523\, C => 
        \I2.END_EVNT2_403\, Y => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__161\);
    
    \I2.PIPE1_DT_42_1_IVL8R_1475\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl40r_net_1\, C => 
        \I2.PIPE1_DT_42l8r_adt_net_50426_\, Y => 
        \I2.PIPE1_DT_42l8r_adt_net_50444_\);
    
    \I2.BNCID_VECT_tile_I_6_1\ : XOR2
      port map(A => \I2.TRGSERVl1r_net_1\, B => 
        \I2.WADDR_REG1l1r\, Y => \I2.I_6_1_i_0_i\);
    
    \I2.REG_0l3r_adt_net_848__adt_net_854228_\ : BFR
      port map(A => \I2.REG_0l3r_adt_net_848__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__adt_net_854228__net_1\);
    
    \I2.N_565_0_adt_net_855728_\ : BFR
      port map(A => \I2.N_565_0\, Y => 
        \I2.N_565_0_adt_net_855728__net_1\);
    
    \I3.PIPEAl16r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_247_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl16r_net_1\);
    
    \I3.VDBi_57l6r_adt_net_143314_\ : AND2
      port map(A => REGl54r, B => \I3.N_2044\, Y => 
        \I3.VDBi_57l6r_adt_net_143314__net_1\);
    
    REGl383r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_284_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl383r\);
    
    \I3.REGMAPl9r_adt_net_854332_\ : BFR
      port map(A => \I3.REGMAPL9R_783\, Y => 
        \I3.REGMAPl9r_adt_net_854332__net_1\);
    
    \I3.STATE1_ns_1_iv_0l3r\ : OR3
      port map(A => \I3.STATE1_ipl8r\, B => 
        \I3.STATE1_nsl3r_adt_net_136441_\, C => 
        \I3.STATE1_nsl3r_adt_net_136439_\, Y => \I3.STATE1_nsl3r\);
    
    \I2.DTO_16_1_IV_0_0L29R_1074\ : AO21
      port map(A => \I2.DTO_1l29r_net_1\, B => \I2.N_196_52\, C
         => \I2.DTO_16_1l29r_adt_net_28730_\, Y => 
        \I2.DTO_16_1l29r_adt_net_28740_\);
    
    \I2.PIPE8_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_555_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl27r_net_1\);
    
    \I3.un51_reg_ads_0_a2_0_a2\ : NOR2
      port map(A => \I3.VASl12r_net_1\, B => \I3.VASl1r_net_1\, Y
         => \I3.N_552\);
    
    \I2.N_2868_1_adt_net_835988_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2868_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.N_2868_1_adt_net_835988_Rd1__net_1\);
    
    RAMAD_padl5r : OB33PH
      port map(PAD => RAMAD(5), A => RAMAD_cl5r);
    
    \I2.N_4254_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4254\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4254_Rd1__net_1\);
    
    \I3.un206_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_641\, Y => 
        \I3.un206_reg_ads_0_a2_1_a3_net_1\);
    
    \I2.L2SERV_919\ : MUX2H
      port map(A => \I2.RPAGEL15R_522\, B => \I2.L2SERV_n3_net_1\, 
        S => \I2.L2SERVe\, Y => \I2.L2SERV_919_net_1\);
    
    \I5.COMMAND_46\ : MUX2H
      port map(A => \I5.COMMANDl9r_net_1\, B => 
        \I5.COMMAND_4l9r_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.COMMAND_46_net_1\);
    
    \I2.un1_end_flush_9_0_0_o2\ : OAI21FTF
      port map(A => \I2.PIPE5_DTL31R_620\, B => 
        \I2.PIPE5_DTL30R_621\, C => \I2.NWPIPE5_net_1\, Y => 
        \I2.un1_NWPIPE5_1_i\);
    
    \I1.REG_74_8_0_324_m9_i_2\ : NAND2FT
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__net_1\, 
        B => \I1.REG_74_8_308_m9_i_1\, Y => 
        \I1.REG_74_1_396_m7_i_3\);
    
    \I2.EVNT_NUM_82\ : NAND2FT
      port map(A => EV_RES_C_569, B => \I2.EVNT_NUMl1r_net_1\, Y
         => \I2.N_1213\);
    
    ADO_padl12r : OB33PH
      port map(PAD => ADO(12), A => ADO_cl12r);
    
    TDCDB_padl12r : IB33
      port map(PAD => TDCDB(12), Y => TDCDB_cl12r);
    
    \I3.VDBi_23l1r_adt_net_145528_\ : NOR3FFT
      port map(A => REGl1r, B => \I3.N_2056\, C => \I3.N_2031\, Y
         => \I3.VDBi_23l1r_adt_net_145528__net_1\);
    
    \I3.RAMAD_VME_26\ : MUX2H
      port map(A => RAMAD_VMEl2r, B => \I3.VASl3r_net_1\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_26_net_1\);
    
    \I2.DT_SRAM_0l8r\ : MUX2L
      port map(A => \I2.PIPE10_DTl8r_net_1\, B => 
        \I2.PIPE5_DTl8r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, Y => 
        \I2.N_876\);
    
    \I2.RAMAD1l1r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_655_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l1r_net_1\);
    
    \I2.un7_bnc_id_1_I_45\ : XOR2
      port map(A => \I2.BNC_IDl8r_net_1\, B => 
        \I2.DWACT_FINC_El4r\, Y => \I2.I_45_0\);
    
    \I3.REG3l2r_1635\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_127_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3L2R_742\);
    
    \I1.REG_74_0_IVL227R_2000\ : AND2
      port map(A => \FBOUTl6r\, B => \I1.N_12233_i\, Y => 
        \I1.REG_74l227r_adt_net_128050_\);
    
    \I3.N_1463_i_1_adt_net_855356_\ : BFR
      port map(A => \I3.N_1463_i_1\, Y => 
        \I3.N_1463_i_1_adt_net_855356__net_1\);
    
    \I2.G_EVNT_NUM_n1_i_o2\ : AND2
      port map(A => \I2.G_EVNT_NUM_i_0_il0r_net_1\, B => 
        \I2.G_EVNT_NUMl1r_net_1\, Y => \I2.N_186\);
    
    \I1.REG_74_0_iv_0l194r\ : AO21
      port map(A => \FBOUTl5r\, B => \I1.REG_4_sqmuxa\, C => 
        \I1.REG_74l194r_adt_net_131097_\, Y => \I1.REG_74l194r\);
    
    \I1.PAGECNTlde_0_o2_2_1237\ : NAND2FT
      port map(A => \I1.N_310_RD1__335\, B => 
        \I1.N_311_i_i_Rd1__adt_net_854920__net_1\, Y => 
        \I1.N_325_499\);
    
    \I1.REG_74_0_IVL183R_2051\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l183r_adt_net_132043_\);
    
    \I2.PIPE10_DT_610\ : MUX2L
      port map(A => \I2.PIPE10_DTl5r_net_1\, B => 
        \I2.PIPE9_DTl5r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_610_net_1\);
    
    REGl370r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_271_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl370r\);
    
    \I3.STATE1_ns_0_iv_0_0l8r\ : AO21
      port map(A => \I3.un1_REGMAP_34\, B => \I3.TCNT_0_sqmuxa_0\, 
        C => \I3.STATE1_nsl8r_adt_net_136092_\, Y => 
        \I3.STATE1_nsl8r\);
    
    \I1.REG_74_i_o2_0_0_364_m9_i_o7\ : NOR2FT
      port map(A => \I1.PAGECNTl6r_adt_net_854924__net_1\, B => 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__net_1\, Y => 
        \I1.REG_74_i_o2_0_0_364_N_14\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I178_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl8r_adt_net_854556__adt_net_855024__net_1\, Y
         => \I2.ADD_21x21_fast_I178_Y_0\);
    
    \I3.REG_1l52r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_153_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl52r);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I154_Y_0_2691\ : AOI21
      port map(A => \I2.PIPE4_DTl15r_net_1\, B => 
        \I2.PIPE4_DTl16r_net_1\, C => \I2.RAMDT4L12R_794\, Y => 
        \I2.N502_i_0_adt_net_490392_\);
    
    \I2.un7_bnc_id_1_I_19\ : AND2
      port map(A => \I2.BNC_IDL3R_585\, B => \I2.DWACT_FINC_El0r\, 
        Y => \I2.N_37\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I25_G0N\ : AND2FT
      port map(A => \I2.LSRAM_OUTl4r\, B => 
        \I2.PIPE7_DTl4r_net_1\, Y => \I2.N242\);
    
    NWRSRAMO_pad : OB33PH
      port map(PAD => NWRSRAMO, A => NWRSRAMO_c);
    
    \I3.PIPEAl13r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_244_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl13r_net_1\);
    
    \I2.L2AS_adt_net_855724_\ : BFR
      port map(A => \I2.L2AS_net_1\, Y => 
        \I2.L2AS_adt_net_855724__net_1\);
    
    \I2.FID_7_0_ivl26r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl26r_net_1\, 
        C => \I2.FID_7l26r_adt_net_18935_\, Y => \I2.FID_7l26r\);
    
    \I2.un1_STATE2_4_i_0_o2_i_a2_i\ : NOR2
      port map(A => \I2.STATE2L4R_291\, B => \I2.STATE2L0R_587\, 
        Y => \I2.N_4182\);
    
    \I2.DT_TEMP_774\ : MUX2H
      port map(A => \I2.DT_TEMPl13r_net_1\, B => 
        \I2.DT_TEMP_7l13r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_774_net_1\);
    
    \I3.PIPEB_110\ : AO21
      port map(A => DPR_cl31r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\, 
        C => \I3.PIPEB_110_adt_net_159411_\, Y => 
        \I3.PIPEB_110_net_1\);
    
    \I2.PIPE5_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_689_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl13r_net_1\);
    
    \I2.MIC_REG3_322\ : MUX2H
      port map(A => \I2.MIC_REG3l5r_net_1\, B => 
        \I2.MIC_REG3l6r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768__net_1\, Y => 
        \I2.MIC_REG3_322_net_1\);
    
    \I2.ROFFSET_c5\ : NAND2
      port map(A => \I2.ROFFSETl5r_net_1\, B => 
        \I2.ROFFSET_c4_net_1\, Y => \I2.ROFFSET_c5_net_1\);
    
    \I1.REG_74_12_300_m8_i\ : OA21FTT
      port map(A => \I1.N_127_i\, B => 
        \I1.REG_74_12_300_m8_i_0_adt_net_120083_\, C => 
        \I1.REG_74_12_300_N_11_adt_net_120111_\, Y => 
        \I1.REG_74_12_300_N_11\);
    
    \I3.PULSEl7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_337_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl7r);
    
    \I2.TRGSERVl2r_1476\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l2r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVL2R_583\);
    
    \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288_\ : BFR
      port map(A => \I3.un1_STATE2_7_1_adt_net_1473__net_1\, Y
         => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\);
    
    \I3.STATE1_ILLEGAL_2127\ : AO21
      port map(A => \I3.STATE1_IPL9R_11\, B => 
        \I3.N_1168_adt_net_1509__net_1\, C => 
        \I3.N_1193_ip_adt_net_136530_\, Y => 
        \I3.N_1193_ip_adt_net_136550_\);
    
    \I2.CRC32_1_sqmuxa_1_i_o2\ : OR2
      port map(A => \I2.STATE2L4R_291\, B => \I2.STATE2L3R_439\, 
        Y => \I2.N_4261\);
    
    \I2.FCNTl2r_1492\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_945_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.FCNTL2R_599\);
    
    \I2.DT_SRAMl5r\ : MUX2L
      port map(A => \I2.N_873\, B => \I2.PIPE2_DTl5r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__489\, Y => 
        \I2.DT_SRAMl5r_net_1\);
    
    \I2.PIPE5_DT_6_0l4r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l4r\, B => 
        \I2.un27_pipe5_dt0l4r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1073\);
    
    \I2.FIFO_FULL\ : DFFC
      port map(CLK => CLK_c, D => PAF_c_i_0, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.FIFO_FULL_net_1\);
    
    \I3.REG_1l6r\ : AO21
      port map(A => \I3.REG1l6r_net_1\, B => \I3.REG2l6r_net_1\, 
        C => \REGl6r_adt_net_14043_\, Y => REGl6r);
    
    \I5.AIR_PULSE_64\ : MUX2H
      port map(A => \I5.AIR_PULSE_net_1\, B => 
        \I5.AIR_PULSE_3_net_1\, S => TICKL0R_3, Y => 
        \I5.AIR_PULSE_64_net_1\);
    
    \I3.UN6_TCNT1_2099\ : NOR2
      port map(A => \I3.TCNT1l4r_net_1\, B => 
        \I3.TCNT1_i_0_il1r_net_1\, Y => 
        \I3.un6_tcnt1_adt_net_134941_\);
    
    \I2.LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_45_TZ_943\ : NOR2
      port map(A => LEAD_FLAGl2r, B => \I2.PIPE4_DTl21r_net_1\, Y
         => \I2.N_2327_tz_adt_net_16395_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I100_Y\ : AO21
      port map(A => \I2.N313_0\, B => \I2.N466_adt_net_71184_\, C
         => \I2.N340\, Y => \I2.N466\);
    
    \I2.PIPE1_DT_42_1_IVL29R_1355\ : OAI21TTF
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100__net_1\, B
         => \I2.TDCDASl28r_net_1\, C => \I2.TDCDASl29r_net_1\, Y
         => \I2.PIPE1_DT_42l29r_adt_net_45714_\);
    
    \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084_\ : BFR
      port map(A => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855088__net_1\, Y
         => \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\);
    
    \I2.OFFSET_37_17l0r\ : MUX2L
      port map(A => \I2.N_755\, B => \I2.N_747\, S => 
        \I2.PIPE7_DTL26R_351\, Y => \I2.N_763\);
    
    \I2.CRC32_12_il26r\ : NOR2
      port map(A => \I2.N_2867_1_adt_net_854964__net_1\, B => 
        \I2.N_127_i_0_i_0\, Y => \I2.N_3943\);
    
    \I2.STATEE_ILLEGAL_1030\ : XOR2FT
      port map(A => \I2.STATEe_ipl0r\, B => \I2.N_3453\, Y => 
        \I2.N_3457_ip_adt_net_23081_\);
    
    \I2.PIPE1_DT_42_0_0l27r_961\ : NOR3
      port map(A => \I2.PIPE1_DT_42_0l27r_net_1\, B => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\, C => \I2.N_12169_i\, Y => 
        \I2.PIPE1_DT_42_3_0L28R_339\);
    
    \I2.PIPE8_DT_21l0r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl0r\, B => \I2.N_566\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l0r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I188_Y\ : XOR2FT
      port map(A => \I2.N_2_0\, B => 
        \I2.ADD_21x21_fast_I188_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l18r\);
    
    \I2.SUB8_522_2737\ : AO21
      port map(A => \I2.N477_adt_net_438351_\, B => 
        \I2.SUB8_522_adt_net_551987_\, C => 
        \I2.SUB8_522_adt_net_659162_\, Y => 
        \I2.SUB8_522_adt_net_659169_\);
    
    \I2.STATEE_NSL4R_1023\ : AND3FFT
      port map(A => BNC_RES_E, B => \I2.INT_ERRS_net_1\, C => 
        \I2.STATEe_ipl0r\, Y => \I2.STATEe_nsl4r_adt_net_22922_\);
    
    \I3.PIPEAl6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_237_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl6r_net_1\);
    
    \I2.PIPE8_DT_16_el20r\ : AND2
      port map(A => \I2.N_565_0_adt_net_855728__net_1\, B => 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\, Y => 
        \I2.N_4681_i\);
    
    \I1.N_50_0_ADT_NET_1409__2867\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__863\, B => 
        \I1.N_50_0_ADT_NET_109751__256\, Y => 
        \I1.N_50_0_ADT_NET_1409__281\);
    
    VAD_padl4r : IOB33PH
      port map(PAD => VAD(4), A => \I3.VADml4r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl4r);
    
    \I2.PIPE1_DT_42_0_0l27r_962\ : NOR3
      port map(A => \I2.PIPE1_DT_42_0l27r_net_1\, B => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\, C => \I2.N_12169_i\, Y => 
        \I2.PIPE1_DT_42_3_0L28R_340\);
    
    \I2.MIC_ERR_REGSl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_332_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl3r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I37_Y\ : AND2
      port map(A => \I2.N247\, B => \I2.N244\, Y => \I2.N302\);
    
    \I2.PIPE1_DT_42_1_IVL18R_1403\ : OAI21FTF
      port map(A => REGl438r, B => 
        \I2.N_3234_adt_net_855648__net_1\, C => 
        \I2.PIPE1_DT_42l18r_adt_net_47449_\, Y => 
        \I2.PIPE1_DT_42l18r_adt_net_47455_\);
    
    \I5.BITCNTl0r_1466\ : DFFC
      port map(CLK => CLK_c, D => \I5.BITCNT_86_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.BITCNT_C0_573\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I151_Y_I_A4_0_1553\ : OA21
      port map(A => \I2.PIPE4_DTl16r_net_1\, B => 
        \I2.PIPE4_DTl18r_net_1\, C => \I2.RAMDT4L5R_821\, Y => 
        \I2.N_41_adt_net_54991_\);
    
    \I5.COMMAND_48\ : MUX2H
      port map(A => \I5.COMMANDl11r_net_1\, B => 
        \I5.COMMAND_4l11r_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.COMMAND_48_net_1\);
    
    \I2.ROFFSETl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_918_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl0r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I189_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl19r_net_1\, Y => 
        \I2.ADD_21x21_fast_I189_Y_0\);
    
    \I2.DT_TEMPl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_774_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl13r_net_1\);
    
    \I1.REG_74_0_IVL314R_1902\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l314r_adt_net_119561_\);
    
    N_1_I3_TCNT3_c2 : AND2
      port map(A => \I3.TCNT3_i_0_il2r_net_1\, B => \I3.TCNT3_c1\, 
        Y => \I3.TCNT3_c2\);
    
    \I3.STATE1_TR24_I_0_A3_5_2114\ : AO21FTT
      port map(A => \I3.STATE1_tr24_i_0_o2_1_i\, B => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135544_\, C => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135637_\, Y => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135642_\);
    
    \I1.sstatel7r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.sstate_ns_0_iv_0_il3r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel7r_net_1\);
    
    \I3.VDBI_57_0_IV_0L27R_2150\ : AO21
      port map(A => \I3.VDBil27r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l27r_adt_net_138431_\, Y => 
        \I3.VDBi_57l27r_adt_net_138441_\);
    
    \I3.VDBi_31l25r\ : MUX2L
      port map(A => \I3.REGl158r\, B => \I3.VDBi_20l25r\, S => 
        \I3.REGMAPl17r_adt_net_854284__net_1\, Y => 
        \I3.VDBi_31l25r_net_1\);
    
    \I3.un10_reg_ads_0_a2_0_a3\ : NOR3
      port map(A => \I3.N_546\, B => \I3.N_578\, C => \I3.N_553\, 
        Y => \I3.un10_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.PIPE6_DT_0_sqmuxa_i_m2_2\ : MUX2L
      port map(A => LEAD_FLAGl7r, B => LEAD_FLAGl5r, S => 
        \I2.PIPE5_DTL22R_665\, Y => \I2.N_4545\);
    
    \I3.PIPEA1_12l21r\ : AND2
      port map(A => DPR_cl21r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854496__net_1\, Y => 
        \I3.PIPEA1_12l21r_net_1\);
    
    \I2.DT_SRAM_0l30r\ : MUX2H
      port map(A => \I2.PIPE5_DTL30R_622\, B => 
        \I2.PIPE10_DTl30r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854228__net_1\, Y => 
        \I2.N_898\);
    
    \I2.SUB8l18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_521_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_3562_i\);
    
    \I3.VASl12r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_74_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl12r_net_1\);
    
    \I2.UN1_STATE1_39_6_1529\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855232__net_1\, B => 
        \I2.ERR_WORDS_RDY_net_1\, C => 
        \I2.un1_STATE1_39_6_i_adt_net_52470_\, Y => 
        \I2.un1_STATE1_39_6_i_adt_net_52472_\);
    
    \I2.DTO_1_896\ : MUX2L
      port map(A => \I2.DTO_1l22r_Rd1__net_1\, B => 
        \I2.DTO_16_1l22r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834760_Rd1__net_1\, Y
         => \I2.DTO_1l22r\);
    
    \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080_\ : BFR
      port map(A => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855088__net_1\, Y
         => \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\);
    
    \I2.DTO_16_1_IV_0_0L6R_1190\ : AND2
      port map(A => \I2.N_4671_adt_net_854600__net_1\, B => 
        \I2.DT_TEMPl6r_net_1\, Y => 
        \I2.DTO_16_1l6r_adt_net_33910_\);
    
    \I3.TCNT3_n3\ : XOR2
      port map(A => \I3.TCNT3l3r_net_1\, B => \I3.TCNT3_c2\, Y
         => \I3.TCNT3_n3_net_1\);
    
    \I2.L2TYPEl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_598_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_i_0_il9r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I187_Y\ : XOR2FT
      port map(A => \I2.N502_i\, B => 
        \I2.ADD_21x21_fast_I187_Y_0\, Y => 
        \I2.un27_pipe5_dt0l17r\);
    
    N_1_I3_TCNT2_389 : MUX2H
      port map(A => \I3.TCNT2l7r_net_1\, B => \N_1.I3.TCNT2_n7\, 
        S => TICKL0R_558, Y => TCNT2_389);
    
    \I2.DTE_1_853\ : MUX2L
      port map(A => \I2.DTE_1l13r_Rd1__net_1\, B => 
        \I2.DTE_21_1l13r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, Y => 
        \I2.DTE_1l13r\);
    
    \I3.VDBi_370\ : MUX2L
      port map(A => \I3.VDBil30r_net_1\, B => \I3.VDBi_57l30r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_370_net_1\);
    
    \I3.N_264_0_adt_net_1653_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.N_264_0_adt_net_1653_Ra1__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.N_264_0_adt_net_1653_Rd1__net_1\);
    
    \I3.RAMDTSl2r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl2r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl2r_net_1\);
    
    DTO_padl24r : IOB33PH
      port map(PAD => DTO(24), A => \I2.DTO_1l24r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl24r);
    
    \I2.RAMAD1_12l9r\ : MUX2L
      port map(A => \I2.TDCDASl7r_net_1\, B => 
        \I2.TDCDBSl7r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855180__net_1\, Y => 
        \I2.RAMAD1_12l9r_net_1\);
    
    \I2.N_2868_1_adt_net_836004_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2868_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.N_2868_1_adt_net_836004_Rd1__net_1\);
    
    \I2.CHAINA_EN244_i_adt_net_855260_\ : BFR
      port map(A => \I2.CHAINA_EN244_i_adt_net_855264__net_1\, Y
         => \I2.CHAINA_EN244_i_adt_net_855260__net_1\);
    
    \I1.REG_1_82\ : MUX2H
      port map(A => \REGl181r\, B => \I1.REG_74l181r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\, Y => 
        \I1.REG_1_82_net_1\);
    
    REGl307r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_208_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl307r\);
    
    \I2.FID_7_0_ivl23r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl23r_net_1\, 
        C => \I2.FID_7l23r_adt_net_19217_\, Y => \I2.FID_7l23r\);
    
    \I5.REG_1_36\ : MUX2L
      port map(A => \I5.TEMPDATAl3r_net_1\, B => REGl423r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_36_net_1\);
    
    RAMDT_padl6r : IOB33PH
      port map(PAD => RAMDT(6), A => \I1.RAMDT_SPI_1l6r_net_1\, 
        EN => \I1.RAMDT_SPI_e_net_1\, Y => RAMDT_inl6r);
    
    \I2.SUB8_522_2735\ : AND2FT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855156__net_1\, B
         => \I2.SUB8l19r_net_1\, Y => 
        \I2.SUB8_522_adt_net_659162_\);
    
    VDB_padl30r : IOB33PH
      port map(PAD => VDB(30), A => \I3.VDBml30r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl30r);
    
    \I2.DTE_21_1_IV_0_0_18_M7_1219\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.G_EVNT_NUMl2r_net_1\, 
        C => \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35893_\, Y => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35905_\);
    
    \I3.PIPEA_8l26r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854456__net_1\, B => 
        \I3.N_235\, Y => \I3.PIPEA_8l26r_net_1\);
    
    \I2.PHASE_862\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_C_240);
    
    \I2.PIPE4_DTl17r_1528\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl17r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL17R_635\);
    
    \I3.PIPEA1l8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_306_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l8r_net_1\);
    
    \I3.REG_1l64r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_165_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl64r);
    
    \I2.DT_TEMP_777\ : MUX2H
      port map(A => \I2.DT_TEMPl16r_net_1\, B => 
        \I2.DT_TEMP_7l16r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_777_net_1\);
    
    \I2.RAMDT4L12R_3073\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_827\);
    
    \I3.VDBi_57_0_ivl10r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855380__net_1\, B => 
        \I3.VDBi_43l10r_net_1\, C => 
        \I3.VDBi_57l10r_adt_net_141884_\, Y => \I3.VDBi_57l10r\);
    
    \I3.REG_1_193\ : MUX2L
      port map(A => VDB_inl12r, B => \I3.REGl145r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, Y => 
        \I3.REG_1_193_0\);
    
    \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__2829\ : OAI21TTF
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100__net_1\, B
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        C => \I2.FIRST_TDC_1_sqmuxa_net_1\, Y => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__173\);
    
    \I3.VDBm_0l28r\ : MUX2L
      port map(A => \I3.PIPEAl28r_net_1\, B => 
        \I3.PIPEBl28r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_170\);
    
    \I2.STATE1_ns_i_o3l4r\ : NAND2
      port map(A => \I2.CHAINA_EN244_i\, B => 
        \I2.CHAINB_EN244_c_0\, Y => \I2.N_3283\);
    
    \I2.PIPE8_DT_542\ : MUX2L
      port map(A => \I2.PIPE8_DTl14r_net_1\, B => 
        \I2.PIPE8_DT_21l14r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_542_net_1\);
    
    \I1.REG_74_0_iv_0l364r\ : AO21
      port map(A => \REGl364r\, B => \I1.N_661\, C => 
        \I1.REG_74l364r_adt_net_114525_\, Y => \I1.REG_74l364r\);
    
    \I5.BITCNT_N1_I_913\ : OA21TTF
      port map(A => \I5.BITCNT_c0\, B => \I5.BITCNTl1r_net_1\, C
         => \I5.N_144\, Y => \I5.N_52_adt_net_9528_\);
    
    \I2.PIPE8_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_554_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl26r_net_1\);
    
    \I2.DTO_1l23r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l23r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l23r_Rd1__net_1\);
    
    \I2.CRC32_12_i_m2l20r\ : MUX2H
      port map(A => \I2.DT_SRAMl20r_net_1\, B => 
        \I2.DT_TEMPl20r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854432__net_1\, Y => 
        \I2.N_3962_i_i\);
    
    \I5.sstate1se_3_i\ : MUX2H
      port map(A => \I5.sstate1l9r_net_1\, B => 
        \I5.sstate1l10r_net_1\, S => TICKl0r, Y => 
        \I5.sstate1se_3_i_net_1\);
    
    \I3.VDBil9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_349_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil9r_net_1\);
    
    \I2.PIPE10_DT_17_i_0l20r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855592__net_1\, B => 
        \I2.PIPE9_DTl20r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l20r_net_1\);
    
    \I3.VASl10r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_72_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VAS_i_0_il10r\);
    
    \I2.DT_SRAMl23r\ : MUX2L
      port map(A => \I2.N_891\, B => \I2.PIPE2_DTl23r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668__net_1\, 
        Y => \I2.DT_SRAMl23r_net_1\);
    
    \I2.BNCID_VECTwa12_1\ : NOR2
      port map(A => \I2.TRGARRl0r_net_1\, B => 
        \I2.TRGARRl1r_net_1\, Y => \I2.BNCID_VECTwa12_1_net_1\);
    
    \I3.REG_1l154r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_202_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl154r\);
    
    \I3.STATE1_414\ : OR2
      port map(A => \I3.STATE1_ipl5r\, B => 
        \I3.N_1180_adt_net_1502__net_1\, Y => \I3.N_1180\);
    
    \I1.BYTECNT_N5_I_0_1780\ : XOR2
      port map(A => \I1.BYTECNTl5r_net_1\, B => \I1.N_334\, Y => 
        \I1.N_75_adt_net_109200_\);
    
    DTE_padl12r : IOB33PH
      port map(PAD => DTE(12), A => \I2.DTE_1l12r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl12r);
    
    \I3.RAMDTSl10r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl10r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl10r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I183_Y\ : XOR2FT
      port map(A => \I2.N513_i\, B => 
        \I2.ADD_21x21_fast_I183_Y_0\, Y => 
        \I2.un27_pipe5_dt0l13r\);
    
    \I2.PIPE1_DT_42_1_ivl22r\ : OR3
      port map(A => \I2.PIPE1_DT_42l22r_adt_net_46751_\, B => 
        \I2.PIPE1_DT_42l22r_adt_net_46763_\, C => 
        \I2.PIPE1_DT_42l22r_adt_net_46764_\, Y => 
        \I2.PIPE1_DT_42l22r\);
    
    \I2.UN1_STATE1_38_0_1532\ : NOR3
      port map(A => \I2.STATE1l17r_net_1\, B => \I2.N_3358\, C
         => \I2.STATE1_i_0_il16r\, Y => 
        \I2.un1_STATE1_38_adt_net_52564_\);
    
    \I2.DTO_16_1_IV_0L4R_1201\ : AO21
      port map(A => \I2.N_197_150\, B => \I2.DT_SRAMl4r_net_1\, C
         => \I2.DTO_16_1l4r_adt_net_34374_\, Y => 
        \I2.DTO_16_1l4r_adt_net_34386_\);
    
    \I3.VDBi_57l7r_adt_net_143036_\ : AO21
      port map(A => \I3.REGl98r\, B => \I3.N_2045\, C => 
        \I3.VDBi_57l7r_adt_net_143035__net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_143036__net_1\);
    
    \I2.CRC32_12_il5r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_131_i_0_i_0\, Y => 
        \I2.N_3922\);
    
    \I2.TOKOUT_FL_674_adt_net_61290_\ : AO21
      port map(A => \I2.TOKOUTBS_net_1\, B => 
        \I2.STATE1l5r_net_1\, C => \I2.TOKOUT_FL_net_1\, Y => 
        \I2.TOKOUT_FL_674_adt_net_61290__net_1\);
    
    \I2.un1_STATE1_13_0_a2_0_a2\ : OR2
      port map(A => \I2.STATE1L6R_630\, B => \I2.STATE1L7R_633\, 
        Y => \I2.N_3351\);
    
    \I2.PIPE1_DT_42_1_IVL29R_1356\ : OR2FT
      port map(A => \I2.N_3279_0_adt_net_855236__net_1\, B => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\, Y => 
        \I2.PIPE1_DT_42l29r_adt_net_45835_\);
    
    \I2.PIPE5_DT_6_0l8r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l8r\, B => 
        \I2.un27_pipe5_dt0l8r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1077\);
    
    \I2.END_TDC1_0_sqmuxa_1\ : AND3FFT
      port map(A => \I2.un5_tdcgda1_net_1\, B => 
        \I2.un3_tdcgda1_1_adt_net_821__net_1\, C => 
        \I2.TDCGDA1_net_1\, Y => \I2.END_TDC1_0_sqmuxa_1_net_1\);
    
    \I3.RAMAD_VME_40\ : MUX2H
      port map(A => RAMAD_VMEl16r, B => \I3.REGl99r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_40_net_1\);
    
    \I3.N_311_adt_net_854752_\ : BFR
      port map(A => \I3.N_311\, Y => 
        \I3.N_311_adt_net_854752__net_1\);
    
    \I2.WOFFSET_13_il11r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_66\, Y => \I2.N_4254\);
    
    \I2.BNC_IDl2r_1604\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_9_1\, CLR => 
        \I2.N_4622_i_0\, SET => \I2.N_4610_i_0\, Q => 
        \I2.BNC_IDL2R_711\);
    
    \I1.REG_74_2_2l340r\ : OAI21TTF
      port map(A => \I1.PAGECNTL8R_457\, B => 
        \I1.REG_74_8_1_tzl340r_net_1\, C => 
        \I1.REG_74_2_2_il340r_adt_net_117067_\, Y => 
        \I1.REG_74_2_2_il340r\);
    
    \I3.REG_1l140r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_188_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl140r\);
    
    \I2.SUB9l20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_588_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l20r_net_1\);
    
    \I3.N_1174_adt_net_1495_\ : OR2
      port map(A => \I3.STATE1_IPL6R_730\, B => \I3.N_1168\, Y
         => \I3.N_1174_adt_net_1495__net_1\);
    
    \I2.N_4667_1_ADT_NET_1046__2758\ : OAI21FTF
      port map(A => \I2.N_4261\, B => \I2.N_4283_I_0_44\, C => 
        \I2.STATE2L2R_589\, Y => \I2.N_4667_1_ADT_NET_1046__34\);
    
    \I2.OFFSET_37_17l1r\ : MUX2L
      port map(A => \I2.N_756\, B => \I2.N_748\, S => 
        \I2.PIPE7_DTL26R_355\, Y => \I2.N_764\);
    
    \I2.MEM_FULL_i_a3\ : NOR2
      port map(A => \I2.FIFO_FULL_592\, B => \I2.SRAM_FULL_593\, 
        Y => TRM_BUSY_c);
    
    \I3.VDBOFFB_30_IV_0L1R_2473\ : OR3
      port map(A => \I3.VDBoffb_30l1r_adt_net_162937_\, B => 
        \I3.VDBoffb_30l1r_adt_net_162933_\, C => 
        \I3.VDBoffb_30l1r_adt_net_162934_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162940_\);
    
    \I3.VDBOFFA_31_IV_0L2R_2586\ : AND2
      port map(A => \REGl255r\, B => \I3.REGMAPl29r_net_1\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164230_\);
    
    \I3.VDBoffl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_118_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl2r_net_1\);
    
    DPR_padl7r : IB33
      port map(PAD => DPR(7), Y => DPR_cl7r);
    
    \I2.RAMAD1l4r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_658_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l4r_net_1\);
    
    \I2.LSRAM_INl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_404_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl20r_net_1\);
    
    \I2.DTO_16_1_IV_0L20R_1121\ : AO21
      port map(A => \I2.DTO_1l20r\, B => \I2.N_196\, C => 
        \I2.DTO_16_1l20r_adt_net_30778_\, Y => 
        \I2.DTO_16_1l20r_adt_net_30794_\);
    
    \I4.END_FLUSH_2\ : OAI21TTF
      port map(A => \I4.STATE1l1r_net_1\, B => 
        \I4.STATE1l2r_net_1\, C => 
        \I4.END_FLUSH_2_adt_net_15635_\, Y => 
        \I4.END_FLUSH_2_net_1\);
    
    \I3.PIPEA1l7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_305_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l7r_net_1\);
    
    \I2.MTDIAS\ : DFFC
      port map(CLK => CLK_c, D => \I2.MTDIAF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.MTDIAS_net_1\);
    
    REGl313r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_214_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl313r\);
    
    \I3.DSSF1_2_i_i_o3_i_a3\ : AO21
      port map(A => DS0B_c, B => DS1B_c, C => \I3.ASBS_net_1\, Y
         => \I3.N_306\);
    
    \I2.RAMAD1l7r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_661_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l7r_net_1\);
    
    \I5.COMMAND_4l14r\ : AND2FT
      port map(A => REGl7r, B => REGl115r, Y => 
        \I5.COMMAND_4l14r_net_1\);
    
    \I3.VDBi_57_iv_0_0_a2_10l7r\ : OR2FT
      port map(A => \I3.N_2016_318\, B => \I3.REGMAPL14R_733\, Y
         => \I3.N_2017\);
    
    \I1.REG_1_110\ : MUX2H
      port map(A => \REGl209r\, B => \I1.N_1348\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_110_net_1\);
    
    \I3.PIPEA_8l0r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854464__net_1\, B => 
        \I3.N_209\, Y => \I3.PIPEA_8l0r_net_1\);
    
    \I3.REGMAPl5r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un25_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il5r\);
    
    \I2.LEAD_FLAG6l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_639_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl2r);
    
    \I3.TCNTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_382_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTl2r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L7R_2493\ : AND2
      port map(A => \REGl244r\, B => \I3.REGMAPl27r_net_1\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163268_\);
    
    \I3.VDBOFFA_31_IV_0L2R_2587\ : AND2
      port map(A => \REGl215r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.VDBoffa_31l2r_adt_net_164234_\);
    
    \I2.L2TYPE_4_il4r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4448_adt_net_68212_\, C => 
        \I2.N_4448_adt_net_68255_\, Y => \I2.N_4448\);
    
    \I2.PIPE8_DT_16_0l5r\ : MUX2H
      port map(A => \I2.PIPE8_DTl5r_net_1\, B => 
        \I2.PIPE7_DTl5r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_571\);
    
    \I2.DTE_21_1_IV_0L8R_1313\ : AO21FTT
      port map(A => \I2.DTE_cl_0_sqmuxa_2_0\, B => 
        \I2.DT_SRAMl8r_net_1\, C => 
        \I2.DTE_21_1l8r_adt_net_38752_\, Y => 
        \I2.DTE_21_1l8r_adt_net_38753_\);
    
    \I2.L2ARRl0r_1495\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_944_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRL0R_602\);
    
    \I2.PIPE7_DTL27R_2791\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_84\);
    
    \I2.OFFSET_37_27l0r\ : MUX2L
      port map(A => \I2.N_835\, B => \I2.N_819\, S => 
        \I2.PIPE7_DTl25r_net_1\, Y => \I2.N_843\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I139_Y\ : NOR2
      port map(A => \I2.N321_0\, B => \I2.N325_0\, Y => 
        \I2.N400_adt_net_88380_\);
    
    \I3.STATE1_402\ : OR2
      port map(A => \I3.STATE1_IPL9R_731\, B => 
        \I3.N_1168_adt_net_1509__net_1\, Y => \I3.N_1168\);
    
    \I3.PULSEl6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_336_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl6r);
    
    \I2.N_1170_adt_net_1217_\ : OAI21FTF
      port map(A => \I2.STATE3_0_sqmuxa_1_0\, B => \I2.N_3019\, C
         => \I2.ROFFSET_0_sqmuxa_1\, Y => 
        \I2.N_1170_adt_net_1217__net_1\);
    
    \I1.REG_74_1_380_M8_I_0_RD1__2991\ : DFFC
      port map(CLK => CLK_c, D => \I1.REG_74_1_380_m8_i_0_Ra1_\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.REG_74_1_380_M8_I_0_RD1__538\);
    
    \I2.SUB8l13r_adt_net_855564_\ : BFR
      port map(A => \I2.SUB8l13r_net_1\, Y => 
        \I2.SUB8l13r_adt_net_855564__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I11_P0N_i_a4\ : OR2
      port map(A => \I2.RAMDT4L12R_799\, B => 
        \I2.PIPE4_DTl11r_net_1\, Y => \I2.N_91_0\);
    
    \I3.un71_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_583\, B => \I3.N_553\, Y => 
        \I3.un71_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.RESYN_0_I2_LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_47_TZ_944\ : 
        NOR2
      port map(A => LEAD_FLAGl6r, B => \I2.PIPE4_DTl21r_net_1\, Y
         => \I2.N_2329_tz_adt_net_16479_\);
    
    \I2.PIPE1_DT_42_1_ivl5r\ : OR3
      port map(A => \I2.PIPE1_DT_42l5r_adt_net_51177_\, B => 
        \I2.PIPE1_DT_42l5r_adt_net_51186_\, C => 
        \I2.PIPE1_DT_42l5r_adt_net_51187_\, Y => 
        \I2.PIPE1_DT_42l5r\);
    
    ADO_padl15r : OB33PH
      port map(PAD => ADO(15), A => ADO_cl15r);
    
    \I1.BITCNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BITCNT_317_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BITCNTl0r_net_1\);
    
    \I3.VDBoffb_57\ : OR3
      port map(A => \I3.VDBoffb_57_adt_net_162220_\, B => 
        \I3.VDBoffb_30l5r_adt_net_162179_\, C => 
        \I3.VDBoffb_30l5r_adt_net_162180_\, Y => 
        \I3.VDBoffb_57_net_1\);
    
    \I3.N_1463_i_1_adt_net_855348_\ : BFR
      port map(A => \I3.N_1463_i_1\, Y => 
        \I3.N_1463_i_1_adt_net_855348__net_1\);
    
    \I2.DT_SRAM_0l31r\ : MUX2H
      port map(A => \I2.PIPE5_DTl31r_net_1\, B => 
        \I2.PIPE10_DTl31r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854204__net_1\, Y => 
        \I2.N_899\);
    
    \I1.REG_1_109\ : MUX2H
      port map(A => \REGl208r\, B => \I1.N_1347\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_109_net_1\);
    
    \I2.LSRAM_INl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_396_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl12r_net_1\);
    
    \I2.MIC_REG3L2R_3035\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_319_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3L2R_789\);
    
    \I1.N_238_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_238_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_238_Rd1__net_1\);
    
    \I2.PIPE3_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl8r_net_1\);
    
    \I1.REG_74_0_IVL279R_1940\ : NOR2FT
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l279r_adt_net_122807_\);
    
    \I1.REG_1_287\ : MUX2H
      port map(A => \REGl386r\, B => \I1.REG_74l386r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y => 
        \I1.REG_1_287_net_1\);
    
    \I2.PIPE5_DT_680\ : MUX2L
      port map(A => \I2.PIPE5_DTl4r_net_1\, B => 
        \I2.PIPE5_DT_6l4r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_680_net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2431\ : AO21
      port map(A => \REGl328r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l3r_adt_net_162520_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162552_\);
    
    \I2.EVNT_WORDl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_716_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl3r_net_1\);
    
    \I2.PIPE7_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl21r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl21r_net_1\);
    
    \I3.PIPEA_8_0l21r\ : MUX2L
      port map(A => DPR_cl21r, B => \I3.PIPEA1l21r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855360__net_1\, Y => \I3.N_230\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854192_\ : BFR
      port map(A => \I2.N_4667_1_ADT_NET_1046__35\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854192__net_1\);
    
    \I2.DTO_16_1_IV_0_0L25R_1087\ : AND2
      port map(A => \I2.DTO_1l25r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l25r_adt_net_29614_\);
    
    \I2.PIPE5_DT_698\ : MUX2H
      port map(A => \I2.PIPE4_DTl22r_net_1\, B => 
        \I2.PIPE5_DTl22r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_698_net_1\);
    
    \I2.OFFSETl4r_1569\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_564_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL4R_676\);
    
    REGl184r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_85_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl184r\);
    
    \I3.un146_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.N_641\, B => \I3.N_551\, Y => 
        \I3.un146_reg_ads_0_a2_1_a3_net_1\);
    
    \I2.EVNT_NUM_n5_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl5r_net_1\, B => 
        \I2.EVNT_NUM_c4_net_1\, Y => \I2.EVNT_NUM_n5_tz_i\);
    
    \I1.sstatel4r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl6r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel4r_net_1\);
    
    \I2.SUB8l4r_1601\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_507_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8L4R_708\);
    
    \I2.OFFSET_37_13l1r\ : MUX2L
      port map(A => \I2.N_724\, B => \I2.N_708\, S => 
        \I2.PIPE7_DTL25R_686\, Y => \I2.N_732\);
    
    \I2.DTO_16_1l11r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l11r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l11r_Rd1__net_1\);
    
    \I2.DTE_2_1l15r\ : XOR2
      port map(A => \I2.CRC32l11r_net_1\, B => 
        \I2.CRC32l23r_net_1\, Y => \I2.DTE_2_1l15r_net_1\);
    
    \I2.PIPE4_DTl5r_adt_net_854416_\ : BFR
      port map(A => \I2.PIPE4_DTl5r_net_1\, Y => 
        \I2.PIPE4_DTl5r_adt_net_854416__net_1\);
    
    \I2.RAMADl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l11r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl11r);
    
    \I2.PIPE7_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl26r_net_1\);
    
    \I3.REG_1_149\ : MUX2L
      port map(A => VDB_inl0r, B => REGl48r, S => 
        \I3.N_1935_adt_net_855332__net_1\, Y => \I3.REG_1_149_0\);
    
    \I2.WOFFSET_838\ : MUX2L
      port map(A => \I2.WOFFSETl11r_Rd1__net_1\, B => 
        \I2.N_4254_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835304_Rd1__net_1\, Y
         => \I2.WOFFSETl11r\);
    
    \I2.SUB8l15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_518_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l15r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I137_Y_i\ : OR3FTT
      port map(A => \I2.N_92_0\, B => \I2.N_40_0_adt_net_577293_\, 
        C => \I2.N_40_0_adt_net_577295_\, Y => \I2.N_40_0\);
    
    \I1.N_50_0_ADT_NET_1409__2748\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__200\, B => 
        \I1.N_50_0_ADT_NET_109751__257\, Y => 
        \I1.N_50_0_ADT_NET_1409__21\);
    
    \I2.CHAINB_ERRF1_493\ : MUX2H
      port map(A => CHAINB_ERR_c, B => \I2.CHAINB_ERRF1_net_1\, S
         => \I2.N_3876_adt_net_855252__net_1\, Y => 
        \I2.CHAINB_ERRF1_493_net_1\);
    
    \I2.DTO_1l11r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l11r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l11r_Rd1__net_1\);
    
    \I3.PIPEA_8_0l16r\ : MUX2L
      port map(A => DPR_cl16r, B => \I3.PIPEA1l16r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855348__net_1\, Y => \I3.N_225\);
    
    \I2.REG_1_n15\ : XOR2
      port map(A => \I2.N_3843\, B => \I2.REG_1_n15_0_net_1\, Y
         => \I2.REG_1_n15_net_1\);
    
    \I2.TOKOUTAS\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKOUTAS_3_i_net_1\, 
        Q => \I2.TOKOUTAS_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I148_Y_0\ : XOR2FT
      port map(A => \I2.SUB8l11r_adt_net_855580__net_1\, B => 
        \I2.SUB8l12r_adt_net_855576__net_1\, Y => 
        \I2.ADD_18x18_fast_I148_Y_0\);
    
    \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100_\ : BFR
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855104__net_1\, Y
         => \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100__net_1\);
    
    \I2.STATEel0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATEe_nsl4r_net_1\, CLR
         => \I2.STATEe_i_0l0r_net_1\, Q => \I2.STATEe_ipl0r\);
    
    \I2.ROFFSET_n7\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\, B => 
        \I2.ROFFSET_n7_tz_i\, Y => \I2.ROFFSET_n7_net_1\);
    
    \I2.NWRSRAM_TST\ : DFFS
      port map(CLK => \I2.CLK_sram\, D => \I2.WREi_net_1\, SET
         => \HWRES_3_adt_net_738__net_1\, Q => NWRSRAM_TST_c);
    
    \I3.VDBi_52l1r\ : MUX2H
      port map(A => \I3.VDBil1r_net_1\, B => \FBOUTl1r\, S => 
        \I3.N_57_i_0_0_adt_net_854696__net_1\, Y => 
        \I3.VDBi_52l1r_net_1\);
    
    \I3.VDBi_57_iv_0_0_a2_12l7r\ : AND2
      port map(A => \I3.N_2016\, B => \I3.REGMAPL14R_734\, Y => 
        \I3.N_2045\);
    
    \I3.N_1463_i_1_adt_net_855360_\ : BFR
      port map(A => \I3.N_1463_i_1\, Y => 
        \I3.N_1463_i_1_adt_net_855360__net_1\);
    
    \I2.PIPE4_DTl11r_1148_1736\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL11R_843\);
    
    \I1.REG_18_sqmuxa_adt_net_855476_\ : BFR
      port map(A => \I1.REG_18_sqmuxa\, Y => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\);
    
    \I1.REG_74_0_IVL222R_2005\ : AND2
      port map(A => \FBOUTl1r\, B => \I1.N_12233_i\, Y => 
        \I1.REG_74l222r_adt_net_128480_\);
    
    \I2.PIPE3_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl5r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl5r_net_1\);
    
    \I1.SBYTE_8_i_0l7r\ : OA21
      port map(A => \I1.N_602_i\, B => REGl90r, C => 
        \I1.N_1194_adt_net_106064_\, Y => \I1.N_1194\);
    
    \I5.REG_1_21\ : MUX2H
      port map(A => \I5.TEMPDATAl2r_net_1\, B => REGl438r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_21_net_1\);
    
    \I2.MIC_ERR_REGSl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_353_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl24r_net_1\);
    
    \I3.VDBI_57_0_IVL10R_2214\ : AO21
      port map(A => \I3.PIPEAl10r_net_1\, B => \I3.N_90_i_0_1\, C
         => \I3.VDBi_57l10r_adt_net_141874_\, Y => 
        \I3.VDBi_57l10r_adt_net_141883_\);
    
    \I2.STATE2l5r_1246\ : DFFS
      port map(CLK => CLK_c, D => \I2.N_2796_i_0\, SET => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L5R_508\);
    
    \I2.L2SERV_921\ : MUX2H
      port map(A => \I2.RPAGEl13r\, B => \I2.L2SERV_n1_net_1\, S
         => \I2.L2SERVe\, Y => \I2.L2SERV_921_net_1\);
    
    L1A_pad : IB33
      port map(PAD => L1A, Y => L1A_c);
    
    \I2.RAMDT4L8R_2980\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl8r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L8R_527\);
    
    \I2.L2TYPE_4_IL14R_1616\ : NAND2FT
      port map(A => \I2.N_4455\, B => \I2.N_4456\, Y => 
        \I2.N_4438_adt_net_66932_\);
    
    \I3.REGMAPL28R_2988\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un121_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL28R_535\);
    
    \I2.DTE_21_1_IV_0L13R_1285\ : AND2
      port map(A => \I2.DTE_1l13r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1l13r_adt_net_38171_\);
    
    \I2.DTOSl8r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl8r, Q => 
        \I2.DTOSl8r_net_1\);
    
    \I2.OFFSET_37_2l7r\ : MUX2L
      port map(A => \REGl388r\, B => \REGl324r\, S => 
        \I2.PIPE7_DTL27R_66\, Y => \I2.N_650\);
    
    \I2.END_EVNT5\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT5_net_1\);
    
    \I5.COMMAND_49\ : MUX2H
      port map(A => \I5.COMMANDl12r_net_1\, B => 
        \I5.COMMAND_4l12r_net_1\, S => \I5.sstate1l13r_net_1\, Y
         => \I5.COMMAND_49_net_1\);
    
    \I3.PIPEA_250\ : MUX2L
      port map(A => \I3.PIPEAl19r_net_1\, B => 
        \I3.PIPEA_8l19r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854664__net_1\, Y
         => \I3.PIPEA_250_net_1\);
    
    \I1.REG_1_118\ : MUX2H
      port map(A => \REGl217r\, B => \I1.REG_74l217r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_118_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl13r\ : OR3
      port map(A => \I2.PIPE1_DT_42l13r_adt_net_49201_\, B => 
        \I2.PIPE1_DT_42l13r_adt_net_49210_\, C => 
        \I2.PIPE1_DT_42l13r_adt_net_49211_\, Y => 
        \I2.PIPE1_DT_42l13r\);
    
    \I3.REG_1_279\ : MUX2H
      port map(A => VDB_inl7r, B => \I3.REGl98r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_279_0\);
    
    \I1.REG_16_sqmuxa_0_a2_0_718\ : OR2FT
      port map(A => \I1.PAGECNT_0l9r_adt_net_835132_Rd1__net_1\, 
        B => \I1.REG_74_1_A0_0L228R_100\, Y => \I1.N_253_96\);
    
    \I3.RAMAD_VMEl15r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_39_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl15r);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I91_Y_0\ : AO21TTF
      port map(A => \I2.N_28\, B => \I2.N_2360_tz_tz\, C => 
        \I2.N_17\, Y => \I2.N394\);
    
    \I2.PIPE2_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl20r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl20r_net_1\);
    
    \I5.un1_tick_6_0_a2_0_a2\ : AOI21FTF
      port map(A => \I5.N_155_0_adt_net_983__net_1\, B => 
        \I5.N_81_i_0_i\, C => TICKL0R_556, Y => \I5.N_406\);
    
    \I2.PIPE2_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl6r_net_1\);
    
    SCLB_pad : OB33PH
      port map(PAD => SCLB, A => \I5.N_106\);
    
    \I3.VDBil29r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_369_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil29r_net_1\);
    
    \I2.PIPE1_DT_30l15r\ : MUX2L
      port map(A => \I2.TDCDBSl15r_net_1\, B => 
        \I2.TDCDBSl13r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, Y
         => \I2.PIPE1_DT_30l15r_net_1\);
    
    REGl387r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_288_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl387r\);
    
    \I2.OFFSET_37_27l1r\ : MUX2L
      port map(A => \I2.N_836\, B => \I2.N_820\, S => 
        \I2.PIPE7_DTl25r_net_1\, Y => \I2.N_844\);
    
    \I2.PIPE7_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl22r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl22r_net_1\);
    
    \I2.CRC32_821\ : MUX2L
      port map(A => \I2.CRC32l26r_net_1\, B => \I2.N_3943\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_821_net_1\);
    
    \I1.BYTECNT_i_0_il4r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_310_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.BYTECNT_i_0_il4r_net_1\);
    
    \I2.N_4283_i_0_a2_m1_e_0_666\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__48\, B => 
        \I2.TEMPF_adt_net_855740__net_1\, Y => \I2.N_4283_I_0_44\);
    
    \I2.CRC32_12_i_0_x2l6r\ : XOR2FT
      port map(A => \I2.CRC32l6r_net_1\, B => \I2.N_225_i_i\, Y
         => \I2.N_251_i_i_0\);
    
    DTE_padl16r : IOB33PH
      port map(PAD => DTE(16), A => \I2.DTE_1l16r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl16r);
    
    \I3.VDBi_40_0_i_m2l12r\ : MUX2L
      port map(A => REGl430r, B => REGl446r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_1857\);
    
    \I2.DT_TEMPl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_762_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl1r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0_o2_1\ : OR2
      port map(A => \I2.N_128_0\, B => \I2.N_74_adt_net_55281_\, 
        Y => \I2.N_74\);
    
    \I2.DTE_1_845\ : MUX2L
      port map(A => \I2.DTE_1l5r_net_1\, B => \I2.DTE_21_1l5r\, S
         => \I2.N_2868_1\, Y => \I2.DTE_1_845_net_1\);
    
    \I2.OFFSET_37_8l1r\ : MUX2L
      port map(A => \REGl358r\, B => \REGl294r\, S => 
        \I2.PIPE7_DTL27R_73\, Y => \I2.N_692\);
    
    \I5.REG_1l438r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_21_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl438r);
    
    \I2.MIC_REG3L3R_2967\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_320_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3L3R_484\);
    
    \I3.VDBoffa_31_iv_0l3r\ : AND2
      port map(A => \REGl176r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        Y => \I3.VDBoffa_31l3r_adt_net_164024_\);
    
    \I2.PIPE5_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_684_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl8r_net_1\);
    
    \I2.DT_TEMPl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_787_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl26r_net_1\);
    
    \I1.REG_74_0_IVL355R_1858\ : NOR2FT
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_24_sqmuxa_adt_net_854776__net_1\, Y => 
        \I1.REG_74l355r_adt_net_115687_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I120_Y_0_o2_0_729\ : NAND2
      port map(A => \I2.N_64_0\, B => \I2.N_89_0_110\, Y => 
        \I2.N_72_0_107\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I137_Y_I_1574\ : OAI21
      port map(A => \I2.PIPE4_DTL12R_512\, B => 
        \I2.PIPE4_DTl13r_net_1\, C => \I2.RAMDT4L5R_821\, Y => 
        \I2.N_40_adt_net_57971_\);
    
    \I2.G_EVNT_NUMl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_928_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl6r_net_1\);
    
    \I2.DTE_21_1_IV_0L8R_1314\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.DTE_2_1l8r_net_1\, C
         => \I2.DTE_21_1l8r_adt_net_38735_\, Y => 
        \I2.DTE_21_1l8r_adt_net_38754_\);
    
    \I3.VDBOFFA_31_IV_0L3R_2574\ : AO21
      port map(A => \REGl208r\, B => 
        \I3.REGMAPl23r_adt_net_855012__net_1\, C => 
        \I3.VDBoffa_31l3r_adt_net_164036_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164071_\);
    
    \I3.VDBI_57_0_IVL28R_2145\ : AND2
      port map(A => \I3.PIPEAl28r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l28r_adt_net_138305_\);
    
    \I2.SUB8_506\ : MUX2H
      port map(A => \I2.SUB8l3r_net_1\, B => \I2.SUB8_2l3r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855148__net_1\, Y => 
        \I2.SUB8_506_net_1\);
    
    \I2.PIPE8_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_549_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl21r_net_1\);
    
    \I3.UN2_VSEL_2_I_0_2103\ : AND3FFT
      port map(A => AMB_cl1r, B => \I3.N_2055\, C => AMB_cl0r, Y
         => \I3.N_1510_adt_net_135035_\);
    
    \I2.PIPE1_DT_42_1_iv_2l26r\ : OR2
      port map(A => \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46178_\, 
        B => \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46179_\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il26r\);
    
    \I2.PIPE5_DT_6l3r\ : MUX2L
      port map(A => \I2.PIPE4_DTl3r_adt_net_854544__net_1\, B => 
        \I2.N_1072\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, Y => 
        \I2.PIPE5_DT_6l3r_net_1\);
    
    \I3.REG_1l114r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_295_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl114r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I186_Y\ : XOR2
      port map(A => \I2.N_82_0\, B => 
        \I2.ADD_21x21_fast_I186_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l16r\);
    
    \I3.PIPEA1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_303_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l5r_net_1\);
    
    \I5.AIR_PULSE_0_sqmuxa_1_i_o3\ : AND2
      port map(A => \I5.AIR_START_net_1\, B => 
        \I5.sstate2l3r_net_1\, Y => \I5.N_463\);
    
    \I3.NOEAD_c_i\ : NOR2FT
      port map(A => \I3.MBLTCYC_net_1\, B => \I3.ADACKCYC_net_1\, 
        Y => NOEAD_c_i_0);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I180_un1_Y\ : AND2
      port map(A => \I2.N301_2\, B => 
        \I2.I180_un1_Y_adt_net_215260_\, Y => 
        \I2.I180_un1_Y_adt_net_240062_\);
    
    \I3.NRDMEBi\ : DFFS
      port map(CLK => CLK_c, D => \I3.NRDMEBi_230_net_1\, SET => 
        CLEAR_STAT_i_0, Q => NRDMEB_c);
    
    \I1.REG_74_8_0l380r\ : AND2FT
      port map(A => \I1.N_396\, B => \I1.N_185_9_adt_net_112166_\, 
        Y => \I1.N_185_9\);
    
    \I1.PAGECNTlde_0_o4\ : OAI21TTF
      port map(A => \I1.SSTATEL6R_417\, B => \I1.N_591_1\, C => 
        \I1.N_370_adt_net_106316_\, Y => \I1.N_370\);
    
    \I2.MIC_ERR_REGSl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_357_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl28r_net_1\);
    
    \I2.RAMADl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l2r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl2r);
    
    \I5.SSTATE1SE_4_0_0_907\ : AO21
      port map(A => \I5.sstate1l6r_net_1\, B => \I5.N_67\, C => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.sstate1_ns_el5r_adt_net_9070_\);
    
    \I2.PIPE7_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl27r_net_1\);
    
    \I3.VDBOFFA_49_2546\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal5r_net_1\, Y => 
        \I3.VDBoffa_49_adt_net_163738_\);
    
    \I2.STATE1_NS_0L11R_1035\ : AND3FFT
      port map(A => TDCDRYB_c, B => \I2.N_3889\, C => 
        \I2.N_3887_adt_net_855068__net_1\, Y => 
        \I2.STATE1_nsl11r_adt_net_23387_\);
    
    \I3.N_203_adt_net_854976_\ : BFR
      port map(A => \I3.N_203\, Y => 
        \I3.N_203_adt_net_854976__net_1\);
    
    \I2.PIPE5_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_681_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl5r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L6R_2372\ : AND2
      port map(A => \REGl315r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        Y => \I3.VDBoffb_30l6r_adt_net_161958_\);
    
    \I2.WOFFSETl2r_adt_net_854984_\ : BFR
      port map(A => \I2.WOFFSETl2r\, Y => 
        \I2.WOFFSETl2r_adt_net_854984__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I45_Y\ : AND2
      port map(A => \I2.N235\, B => \I2.N232\, Y => \I2.N310\);
    
    \I2.DTE_21_1_IV_2L0R_1344\ : AND2
      port map(A => GA_cl0r, B => 
        \I2.STATE2l1r_adt_net_855120__net_1\, Y => 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39723_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0_o2_1_948\ : 
        OR3FFT
      port map(A => \I2.N_107_0\, B => \I2.N_13_1\, C => 
        \I2.N_95_0\, Y => \I2.N_74_ADT_NET_55281__326\);
    
    \I5.CHAIN_SELECT_4\ : MUX2L
      port map(A => \I5.AIR_CHAIN_net_1\, B => REGl6r, S => 
        REGl7r, Y => \I5.CHAIN_SELECT_4_net_1\);
    
    \I1.UN1_SBYTE13_I_I_I_1_1773\ : AND2
      port map(A => \I1.N_463_1\, B => 
        \I1.un1_sbyte13_i_i_i_1_adt_net_108180_\, Y => 
        \I1.un1_sbyte13_i_i_i_1_adt_net_108267_\);
    
    \I1.RAMDT_SPI_1l1r\ : DFFC
      port map(CLK => CLK_c, D => \FBOUTl1r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.RAMDT_SPI_1l1r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL22R_1381\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_339\, B => 
        \I2.EVNT_NUMl6r_net_1\, Y => 
        \I2.PIPE1_DT_42l22r_adt_net_46751_\);
    
    \I3.VDBi_343\ : MUX2L
      port map(A => \I3.VDBil3r_net_1\, B => \I3.VDBi_57l3r\, S
         => \I3.un1_STATE1_13_1_adt_net_1351__net_1\, Y => 
        \I3.VDBi_343_net_1\);
    
    \I2.STATE3_NSL8R_1046\ : OR3FTT
      port map(A => \I2.STATE3_il8r\, B => \I2.STATE3l6r_net_1\, 
        C => \I2.N_1170_adt_net_1217__adt_net_855700__net_1\, Y
         => \I2.STATE3_nsl8r_adt_net_24815_\);
    
    \I3.STATE1_NS_1_IV_0L3R_2125\ : NOR3FFT
      port map(A => \I3.SINGCYC_881\, B => \I3.N_638\, C => 
        \I3.N_1905_1_adt_net_855384__net_1\, Y => 
        \I3.STATE1_nsl3r_adt_net_136441_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I138_Y_0_a2\ : NOR3FFT
      port map(A => \I2.N_52_0\, B => \I2.N_100_0_adt_net_58633_\, 
        C => \I2.N_74\, Y => \I2.N_100_0\);
    
    \I2.PIPE9_DT_279\ : MUX2L
      port map(A => \I2.PIPE9_DTl10r_net_1\, B => 
        \I2.PIPE8_DTl10r_net_1\, S => \I2.NWPIPE8_i_0_i_0_0\, Y
         => \I2.PIPE9_DT_279_net_1\);
    
    \I2.OFFSET_37_23l1r\ : MUX2L
      port map(A => \REGl270r\, B => \REGl206r\, S => 
        \I2.PIPE7_DTL27R_91\, Y => \I2.N_812\);
    
    \I3.VDBOFFB_30_IV_0L0R_2491\ : OR3
      port map(A => \I3.VDBoffb_30l0r_adt_net_163127_\, B => 
        \I3.VDBoffb_30l0r_adt_net_163123_\, C => 
        \I3.VDBoffb_30l0r_adt_net_163124_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163130_\);
    
    \I3.PIPEB_105\ : AO21
      port map(A => DPR_cl26r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\, 
        C => \I3.PIPEB_105_adt_net_159621_\, Y => 
        \I3.PIPEB_105_net_1\);
    
    \I5.sstate2l0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate2se_3_i_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.sstate2l0r_net_1\);
    
    \I3.REG1_227\ : OAI21FTF
      port map(A => \I3.REG1l405r_net_1\, B => \I3.N_1563\, C => 
        \I3.REG2_15l405r\, Y => \I3.REG1_227_net_1\);
    
    \I3.UN7_RONLY_0_A2_0_A3_2639\ : AND3
      port map(A => \I3.LWORDS_net_1\, B => \I3.VAS_i_0_il15r\, C
         => \I3.un7_ronly_0_a2_0_a3_adt_net_165586_\, Y => 
        \I3.un7_ronly_0_a2_0_a3_adt_net_165588_\);
    
    \I2.PIPE1_DT_42_1_IVL5R_1491\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        B => \I2.PIPE1_DT_12l5r_net_1\, Y => 
        \I2.PIPE1_DT_42l5r_adt_net_51171_\);
    
    \I3.VDBI_57_IV_0_0L6R_2234\ : NOR2FT
      port map(A => \FBOUTl6r\, B => \I3.N_2047\, Y => 
        \I3.VDBi_57l6r_adt_net_143390_\);
    
    \I2.RAMAD1l13r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_667_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l13r_net_1\);
    
    \I3.REG1_133\ : MUX2L
      port map(A => VDB_inl0r, B => \I3.REG1l0r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG1_133_net_1\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_683\ : AO21
      port map(A => 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855220__net_1\, B
         => \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__870\, 
        C => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_adt_net_19813_\, Y
         => \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_61\);
    
    REGl175r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_76_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl175r\);
    
    \I2.OFFSET_37_19l2r\ : MUX2L
      port map(A => \REGl279r\, B => \REGl215r\, S => 
        \I2.PIPE7_DTL27R_90\, Y => \I2.N_781\);
    
    \I1.REG_1_160\ : MUX2H
      port map(A => \REGl259r\, B => \I1.REG_74l259r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_160_net_1\);
    
    \I2.un2_evnt_word_I_72\ : AND2
      port map(A => \I2.WOFFSETl11r\, B => \I2.N_9_1\, Y => 
        \I2.N_4\);
    
    \I2.DTO_9_IVL22R_1105\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl22r_net_1\, C => 
        \I2.DTO_9l22r_adt_net_30286_\, Y => 
        \I2.DTO_9l22r_adt_net_30294_\);
    
    \I2.G_EVNT_NUM_n7_i_o2\ : AND2
      port map(A => \I2.N_198_551\, B => \I2.G_EVNT_NUMl7r_net_1\, 
        Y => \I2.N_201\);
    
    \I3.VDBI_57_0_IV_0L9R_2216\ : AND2
      port map(A => \I3.VDBil9r_net_1\, B => 
        \I3.N_1764_adt_net_854352__net_1\, Y => 
        \I3.VDBi_57l9r_adt_net_142322_\);
    
    \I1.PAGECNT_0l7r_adt_net_835112_Rd1__adt_net_855516_\ : BFR
      port map(A => \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__363\, Y
         => 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__adt_net_855516__net_1\);
    
    \I1.REG_1_159\ : MUX2H
      port map(A => \REGl258r\, B => \I1.REG_74l258r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_159_net_1\);
    
    \I3.VDBi_29l9r_adt_net_142014_\ : NOR3FFT
      port map(A => REGl41r, B => \I3.REGMAPL7R_460\, C => 
        \I3.N_1907_266\, Y => 
        \I3.VDBi_29l9r_adt_net_142014__net_1\);
    
    \I2.N_2828_adt_net_1062__adt_net_835312_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2828_adt_net_1062__net_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.N_2828_adt_net_1062__adt_net_835312_Rd1__net_1\);
    
    \I1.N_238_RD1__2881\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_238_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_238_RD1__313\);
    
    \I2.DTO_16_1l27r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l27r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l27r_Rd1__net_1\);
    
    \I1.REG_74_0_ivl334r\ : AO21
      port map(A => \REGl334r\, B => \I1.N_209\, C => 
        \I1.REG_74l334r_adt_net_117744_\, Y => \I1.REG_74l334r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0\ : AO21FTF
      port map(A => \I2.N_74_104\, B => 
        \I2.N519_0_adt_net_55614_\, C => \I2.N_70_0\, Y => 
        \I2.N519_0\);
    
    \I2.EVNT_WORD_721\ : MUX2H
      port map(A => \I2.EVNT_WORDl8r_net_1\, B => \I2.I_45\, S
         => \I2.N_2864_0_adt_net_854272__net_1\, Y => 
        \I2.EVNT_WORD_721_net_1\);
    
    VDB_padl7r : IOB33PH
      port map(PAD => VDB(7), A => \I3.N_11\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl7r);
    
    \I3.PIPEA1l26r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_324_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l26r_net_1\);
    
    \I3.REG_1l415r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_222_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl415r);
    
    \I2.DTO_1l13r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l13r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l13r_Rd1__net_1\);
    
    \I2.OFFSET_37_1l4r\ : MUX2L
      port map(A => \REGl353r\, B => \REGl289r\, S => 
        \I2.PIPE7_DTL27R_65\, Y => \I2.N_639\);
    
    \I2.FIDl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_432\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl16r);
    
    CHAINA_ERR_pad : IB33
      port map(PAD => CHAINA_ERR, Y => CHAINA_ERR_c);
    
    \I1.N_223_adt_net_854848_\ : BFR
      port map(A => \I1.N_223\, Y => 
        \I1.N_223_adt_net_854848__net_1\);
    
    \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__2840\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__198\);
    
    FID_padl21r : OB33PH
      port map(PAD => FID(21), A => FID_cl21r);
    
    \I2.PIPE10_DT_635\ : MUX2L
      port map(A => \I2.PIPE10_DTl30r_net_1\, B => 
        \I2.PIPE10_DT_17l30r\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_635_net_1\);
    
    \I2.PIPE6_DT_0_sqmuxa_i\ : NOR2
      port map(A => \I2.N_4551\, B => \I2.N_222_adt_net_63455_\, 
        Y => \I2.N_4526\);
    
    \I2.G_EVNT_NUM_n8_i_o2_1287\ : AND2
      port map(A => \I2.N_201\, B => \I2.G_EVNT_NUMl8r_net_1\, Y
         => \I2.N_207_549\);
    
    \I3.VADm_0_a3l7r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl7r_net_1\, Y => \I3.VADml7r\);
    
    \I2.un78_pipe5_dt_1\ : XOR2
      port map(A => \I2.RAMDT4l9r_net_1\, B => 
        \I2.RAMDT4l8r_net_1\, Y => \I2.un78_pipe5_dt_1_net_1\);
    
    \I2.DTO_16_1_IV_0L21R_1114\ : AO21
      port map(A => \I2.N_197_151\, B => \I2.DT_SRAMl21r_net_1\, 
        C => \I2.DTO_16_1l21r_adt_net_30538_\, Y => 
        \I2.DTO_16_1l21r_adt_net_30548_\);
    
    \I2.DT_SRAM_i_0_m2l9r\ : MUX2L
      port map(A => \I2.N_4045\, B => \I2.PIPE2_DTl9r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.N_4047\);
    
    \I3.VDBOFFB_30_IV_0L1R_2467\ : AO21
      port map(A => \REGl358r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        C => \I3.VDBoffb_30l1r_adt_net_162900_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162932_\);
    
    \I3.N_1910_0_adt_net_854340_\ : BFR
      port map(A => \I3.N_1910_0_adt_net_854348__net_1\, Y => 
        \I3.N_1910_0_adt_net_854340__net_1\);
    
    \I1.REG_74_3_I_A2L172R_1817\ : NOR2
      port map(A => \I1.REG_15_sqmuxa_adt_net_1457__net_1\, B => 
        \I1.N_237_adt_net_854804__net_1\, Y => 
        \I1.N_1370_adt_net_112317_\);
    
    \I1.REG_1_174\ : MUX2H
      port map(A => \REGl273r\, B => \I1.REG_74l273r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y => 
        \I1.REG_1_174_net_1\);
    
    \I0.EV_RESF1\ : DFFC
      port map(CLK => CLK_c, D => EV_RESIN_c, CLR => 
        \I0.un4_hwresi_i\, Q => \I0.EV_RESF1_net_1\);
    
    \I1.PAGECNT_n6_i_i_a4_0\ : OR2FT
      port map(A => \I1.UN1_SBYTE13_1_I_1_207\, B => \I1.N_656\, 
        Y => \I1.N_473\);
    
    ADO_padl6r : OB33PH
      port map(PAD => ADO(6), A => ADO_cl6r);
    
    DPR_padl0r : IB33
      port map(PAD => DPR(0), Y => DPR_cl0r);
    
    \I2.FIDl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_443\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl27r);
    
    \I2.STATE3_NS_O3_0L8R_1038\ : OA21
      port map(A => \I2.un28_sram_empty\, B => 
        \I2.un21_sram_empty_NE_net_1\, C => REGl1r, Y => 
        \I2.N_3012_adt_net_24321_\);
    
    \I2.ROFFSETl4r_1768\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_914_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETL4R_874\);
    
    \I2.RAMADl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l6r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl6r);
    
    \I2.SUB9_1_ADD_18x18_fast_I0_S\ : XOR2
      port map(A => \I2.ca\, B => \I2.G_1_5\, Y => \I2.SUB9_1l3r\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I152_Y_0_1572\ : OA21
      port map(A => \I2.PIPE4_DTl17r_net_1\, B => 
        \I2.PIPE4_DTl18r_net_1\, C => \I2.RAMDT4L12R_799\, Y => 
        \I2.N498_0_adt_net_56940_\);
    
    \I3.REGMAPl12r_1639\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un51_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL12R_746\);
    
    \I2.PIPE9_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_278_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl9r_net_1\);
    
    \I2.un1_STATE1_27_0_0_o3\ : AOI21FTT
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855240__net_1\, 
        B => \I2.N_3891\, C => \I2.STATE1l8r_net_1\, Y => 
        \I2.un1_STATE1_27\);
    
    \I3.DSS\ : DFFS
      port map(CLK => CLK_c, D => \I3.DSSF1_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.DSS_9\);
    
    \I2.PIPE1_DT_12l15r\ : MUX2L
      port map(A => \I2.TDCDASl15r_net_1\, B => 
        \I2.TDCDASl13r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, Y
         => \I2.PIPE1_DT_12l15r_net_1\);
    
    \I2.PIPE10_DT_17_0l29r\ : OR3
      port map(A => \I2.PIPE9_DTl29r_net_1\, B => 
        \I2.PIPE10_DT_17l29r_adt_net_64809_\, C => \I2.N_26\, Y
         => \I2.PIPE10_DT_17l29r\);
    
    \I1.REG_74_0_iv_0_a2l372r\ : AND2
      port map(A => \I1.N_238_Rd1__adt_net_854884__net_1\, B => 
        \I1.N_584\, Y => \I1.N_593\);
    
    \I2.TOKENB_CNT_3_0_a2l0r\ : NOR2
      port map(A => \I2.TOKOUTBS_net_1\, B => \I2.TDCDRYBS_net_1\, 
        Y => \I2.N_177\);
    
    \I2.SUB9_1_ADD_18x18_fast_I4_P0N\ : OR2
      port map(A => \I2.N_3541_i_i\, B => \I2.G_1_1\, Y => 
        \I2.N238\);
    
    \I2.START_GIRO_451\ : MUX2L
      port map(A => \I2.STATE1l18r_net_1\, B => 
        \I2.START_GIRO_net_1\, S => \I2.un1_STATE1_21\, Y => 
        \I2.START_GIRO_451_net_1\);
    
    \I2.GIROT\ : DFFC
      port map(CLK => CLK_c, D => \I2.GIROT_452\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.GIROT_net_1\);
    
    \I1.REG_74_0_IVL376R_1823\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l376r_adt_net_112829_\);
    
    TDCDB_padl9r : IB33
      port map(PAD => TDCDB(9), Y => TDCDB_cl9r);
    
    \I2.PIPE1_DT_12l9r\ : MUX2L
      port map(A => \I2.TDCDASl9r_net_1\, B => 
        \I2.TDCDASl7r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, Y
         => \I2.PIPE1_DT_12l9r_net_1\);
    
    \I2.DTE_21_1_IV_0L9R_1304\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855116__net_1\, B => 
        \I2.EVNT_WORDl5r_net_1\, Y => 
        \I2.DTE_21_1l9r_adt_net_38621_\);
    
    \I3.VDBi_43l9r\ : MUX2L
      port map(A => REGl415r, B => \I3.VDBi_40l9r_net_1\, S => 
        \I3.REGMAPl55r_net_1\, Y => \I3.VDBi_43l9r_net_1\);
    
    \I3.ADACKCYC_112\ : MUX2H
      port map(A => \I3.ADACKCYC_net_1\, B => \I3.VSEL_0\, S => 
        \I3.N_1509\, Y => \I3.ADACKCYC_112_net_1\);
    
    \I2.PIPE5_DT_684\ : MUX2L
      port map(A => \I2.PIPE5_DTl8r_net_1\, B => 
        \I2.PIPE5_DT_6l8r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_684_net_1\);
    
    \I1.REG_74_0_iv_0l179r\ : AO21
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, C => 
        \I1.REG_74l179r_adt_net_132424_\, Y => \I1.REG_74l179r\);
    
    \I3.N_90_i_0_a2\ : AND2
      port map(A => \I3.REGMAPl0r_net_1\, B => 
        \I3.STATE1_IPL9R_11\, Y => \I3.N_90_i_0\);
    
    \I2.PIPE1_DT_42_1_IVL29R_1359\ : AO21FTT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        B => \I2.PIPE1_DT_42l29r_adt_net_45714_\, C => 
        \I2.PIPE1_DT_42l29r_adt_net_45836_\, Y => 
        \I2.PIPE1_DT_42l29r_adt_net_45838_\);
    
    \I1.REG_74_0_iv_i_a2l203r\ : AO21
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_1342_adt_net_130275_\, Y => \I1.N_1342\);
    
    \I2.UN1_PIPE1_DT_1_SQMUXA_2_0_999\ : AND2
      port map(A => \I2.TOKOUTBS_net_1\, B => 
        \I2.STATE1l6r_net_1\, Y => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2_adt_net_20482_\);
    
    \I2.DTO_16_1_IV_0_0L26R_1084\ : AO21
      port map(A => \I2.G_EVNT_NUMl10r_net_1\, B => \I2.N_457\, C
         => \I2.DTO_16_1l26r_adt_net_29426_\, Y => 
        \I2.DTO_16_1l26r_adt_net_29437_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I148_Y\ : XOR2
      port map(A => \I2.N460\, B => \I2.ADD_18x18_fast_I148_Y_0\, 
        Y => \I2.SUB9_1l11r\);
    
    \I2.PIPE1_DT_12l10r\ : MUX2L
      port map(A => \I2.TDCDASl10r_net_1\, B => 
        \I2.TDCDASl8r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, Y
         => \I2.PIPE1_DT_12l10r_net_1\);
    
    \I2.EVNT_NUM_n6_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl6r_net_1\, B => 
        \I2.EVNT_NUM_c5_net_1\, Y => \I2.EVNT_NUM_n6_tz_i\);
    
    \I1.REG_74l324r\ : OR2
      port map(A => \I1.REG_19_sqmuxa\, B => 
        \I1.N_193_adt_net_1425__net_1\, Y => \I1.N_193\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022_\ : NAND2
      port map(A => \I2.WOFFSETl0r_net_1\, B => 
        \I2.STATE2l2r_net_1\, Y => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\);
    
    \I3.REG_1l409r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_216_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl409r);
    
    \I2.DTO_16_1l15r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l15r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l15r_Rd1__net_1\);
    
    \I2.BITCNT_n0_0_a5\ : NOR2
      port map(A => \I2.BITCNT_c0\, B => 
        \I2.ERR_WORDS_RDY_0_sqmuxa\, Y => \I2.BITCNT_n0\);
    
    \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835168_Rd1_\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835168_Rd1__net_1\);
    
    DPR_padl3r : IB33
      port map(PAD => DPR(3), Y => DPR_cl3r);
    
    \I1.REG_24_sqmuxa_adt_net_854780_\ : BFR
      port map(A => \I1.REG_24_sqmuxa\, Y => 
        \I1.REG_24_sqmuxa_adt_net_854780__net_1\);
    
    REGl317r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_218_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl317r\);
    
    \I3.TCNTlde_0\ : OR2FT
      port map(A => \I3.N_1904\, B => \I3.un1_STATE1_10_i_0\, Y
         => \I3.TCNTe\);
    
    \I2.PIPE1_DT_758\ : MUX2L
      port map(A => \I2.PIPE1_DTl31r_net_1\, B => 
        \I2.PIPE1_DT_42l31r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854560__net_1\, 
        Y => \I2.PIPE1_DT_758_net_1\);
    
    TDCDA_padl23r : IB33
      port map(PAD => TDCDA(23), Y => TDCDA_cl23r);
    
    \I5.REG_1_26\ : MUX2H
      port map(A => \I5.TEMPDATAl7r_net_1\, B => REGl443r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_26_net_1\);
    
    \I3.VDBi_40_0_i_m2l6r\ : MUX2L
      port map(A => REGl424r, B => REGl440r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_2269\);
    
    \I2.DTESl31r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl31r, Q => 
        \I2.DTESl31r_net_1\);
    
    \I2.PIPE5_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_692_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl16r_net_1\);
    
    \I2.PHASE_865\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_C_243);
    
    \I1.REG_74_0_IV_0L372R_1829\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.N_593\, Y => 
        \I1.REG_74l372r_adt_net_113310_\);
    
    \I2.OFFSET_37_7l0r\ : MUX2L
      port map(A => \I2.N_675\, B => \I2.N_651\, S => 
        \I2.PIPE7_DTL25R_683\, Y => \I2.N_683\);
    
    \I2.DTE_21_1_IV_0L28R_1235\ : AO21FTT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_290\, B => 
        \I2.DT_SRAMl28r_net_1\, C => 
        \I2.DTE_21_1l28r_adt_net_36757_\, Y => 
        \I2.DTE_21_1l28r_adt_net_36758_\);
    
    \I3.REG_1_278\ : MUX2H
      port map(A => VDB_inl6r, B => \I3.REGl97r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_278_0\);
    
    REGl205r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_106_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl205r\);
    
    REGl208r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_109_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl208r\);
    
    \I2.I_1335_ca\ : NAND2FT
      port map(A => \I2.SUB8L3R_710\, B => \I2.OFFSETL0R_586\, Y
         => \I2.ca\);
    
    \I2.LEAD_FLAG6_642_1601\ : NOR2FT
      port map(A => LEAD_FLAGl5r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_642_adt_net_64068_\);
    
    \I1.REG_1_168\ : MUX2H
      port map(A => \REGl267r\, B => \I1.REG_74l267r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y => 
        \I1.REG_1_168_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I178_Y\ : XOR2
      port map(A => \I2.N_3\, B => \I2.ADD_21x21_fast_I178_Y_0\, 
        Y => \I2.un27_pipe5_dt0l8r\);
    
    \I2.PIPE1_DT_42_1_IVL16R_1411\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040__net_1\, 
        B => \I2.PIPE1_DT_12l16r_net_1\, Y => 
        \I2.PIPE1_DT_42l16r_adt_net_47835_\);
    
    \I2.SUB8l4r_1602\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_507_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8L4R_709\);
    
    \I2.DTO_1_903\ : MUX2L
      port map(A => \I2.DTO_1l29r_net_1\, B => \I2.DTO_16_1l29r\, 
        S => \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => 
        \I2.DTO_1_903_net_1\);
    
    \I3.VDBml13r\ : MUX2L
      port map(A => \I3.VDBil13r_net_1\, B => \I3.N_155\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml13r_net_1\);
    
    \I3.VDBm_0l31r\ : MUX2L
      port map(A => \I3.PIPEAl31r_net_1\, B => 
        \I3.PIPEB_i_0_il31r\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_173\);
    
    \I3.STATE1_420\ : OR2
      port map(A => \I3.STATE1_ipl3r_adt_net_854364__net_1\, B
         => \I3.N_1186_adt_net_1488__net_1\, Y => \I3.N_1186\);
    
    \I2.PIPE5_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_694_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl18r_net_1\);
    
    \I2.N_4646_1_adt_net_19637_Ra1_\ : AOI21
      port map(A => \I2.MIC_REG1_304_net_1\, B => 
        \I2.MIC_REG2_312_net_1\, C => \I2.MIC_REG3_320_net_1\, Y
         => \I2.N_4646_1_adt_net_19637_Ra1__net_1\);
    
    \I2.DTO_1_882\ : MUX2L
      port map(A => \I2.DTO_1l8r_Rd1__net_1\, B => 
        \I2.DTO_16_1l8r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834772_Rd1__net_1\, Y
         => \I2.DTO_1l8r\);
    
    \I3.REGMAP_I_0_IL40R_2933\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un181_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL40R_450\);
    
    TDCDA_padl12r : IB33
      port map(PAD => TDCDA(12), Y => TDCDA_cl12r);
    
    \I0.CLEAR_i\ : NOR2FT
      port map(A => REGl18r, B => \I0.CLEAR_adt_net_15818_\, Y
         => \I0.CLEAR_i_0\);
    
    \I3.PIPEBl29r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEB_108_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl29r_net_1\);
    
    \I3.UN1_NOEDTKI_0_SQMUXA_1_0_2314\ : AND3FFT
      port map(A => \I3.DSS_net_1\, B => \I3.PURGED_net_1\, C => 
        \I3.STATE1_ipl5r\, Y => 
        \I3.un1_NOEDTKi_0_sqmuxa_1_adt_net_159322_\);
    
    \I2.CRC32_12_0_0_m2l5r\ : MUX2H
      port map(A => \I2.DT_SRAMl5r_net_1\, B => 
        \I2.DT_TEMPl5r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854428__net_1\, Y => 
        \I2.N_4267_i_i\);
    
    ADLTC_pad : OB33PH
      port map(PAD => ADLTC, A => \GND\);
    
    \I2.PIPE5_DT_6l10r\ : MUX2L
      port map(A => \I2.PIPE4_DTl10r_net_1\, B => \I2.N_1079\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\, Y
         => \I2.PIPE5_DT_6l10r_net_1\);
    
    NOE64R_pad : OB33PH
      port map(PAD => NOE64R, A => NOEAD_c);
    
    \I2.PIPE9_DT_270\ : MUX2L
      port map(A => \I2.PIPE9_DTl1r_net_1\, B => 
        \I2.PIPE8_DTl1r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_270_net_1\);
    
    \I2.PIPE9_DT_269\ : MUX2L
      port map(A => \I2.PIPE9_DTl0r_net_1\, B => 
        \I2.PIPE8_DTl0r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_269_net_1\);
    
    \I2.TRAIL_MIS7_i\ : DFFS
      port map(CLK => CLK_c, D => \I2.TRAIL_MIS6_i_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.TRAIL_MIS7_i_net_1\);
    
    \I2.N_2828_adt_net_1062__adt_net_835308_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2828_adt_net_1062__net_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.N_2828_adt_net_1062__adt_net_835308_Rd1__net_1\);
    
    \I2.PIPE7_DTl10r_1588\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL10R_695\);
    
    \I2.PIPE5_DTl22r_1559\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_698_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL22R_666\);
    
    \I2.STATE3_ns_o3l10r\ : OR3
      port map(A => \I2.DTOS_i_il31r\, B => \I2.DTOSl29r_net_1\, 
        C => \I2.N_3016_adt_net_24530_\, Y => \I2.N_3016\);
    
    \I3.un156_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_585\, Y => 
        \I3.un156_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.CRC32_12_il1r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_999\, Y => 
        \I2.N_3918\);
    
    \I2.N_2828_adt_net_39957_\ : NAND3FFT
      port map(A => \I2.N_2867_1_338\, B => 
        \I2.N_2828_adt_net_39955__net_1\, C => \I2.N_2870\, Y => 
        \I2.N_2828_adt_net_39957__net_1\);
    
    \I2.REG_1_c3_i\ : AO21
      port map(A => REGl35r, B => \I2.N_3832_adt_net_101495_\, C
         => \I2.N_3832_adt_net_101536_\, Y => \I2.N_3832\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855468_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__21\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\);
    
    \I2.WOFFSET_13_il3r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_13_1\, Y => 
        \I2.N_4246\);
    
    \I2.un1_tdc_res_32_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl409r, Y => 
        \I2.N_4613_i_0\);
    
    \I2.L2ARR_n3\ : XOR2
      port map(A => \I2.L2ARRl3r_net_1\, B => \I2.L2ARR_c2_net_1\, 
        Y => \I2.L2ARR_n3_net_1\);
    
    \I2.RAMAD1l17r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_671_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l17r_net_1\);
    
    \I3.un975_regmap_3_i_0_o2_i_a2\ : AND3FFT
      port map(A => \I3.REGMAPL34R_446\, B => \I3.REGMAPL33R_461\, 
        C => \I3.N_560_adt_net_134484_\, Y => \I3.N_560\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854564_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854564__net_1\);
    
    \I2.G_EVNT_NUM_n10_0\ : MUX2L
      port map(A => \I2.N_285_1\, B => 
        \I2.G_EVNT_NUM_n10_0_a2_0_0_i\, S => \I2.N_218\, Y => 
        \I2.G_EVNT_NUM_n10\);
    
    \I2.OFFSET_37_29l2r\ : MUX2L
      port map(A => \I2.N_853\, B => \I2.N_741\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l2r\);
    
    \I1.SBYTE_8_0_il6r\ : OA21
      port map(A => \I1.N_602_i\, B => REGl89r, C => 
        \I1.N_206_adt_net_105994_\, Y => \I1.N_206\);
    
    \I2.PIPE1_DT_42_1_ivl14r\ : OR3
      port map(A => \I2.PIPE1_DT_42l14r_adt_net_48954_\, B => 
        \I2.PIPE1_DT_42l14r_adt_net_48963_\, C => 
        \I2.PIPE1_DT_42l14r_adt_net_48964_\, Y => 
        \I2.PIPE1_DT_42l14r\);
    
    \I3.VDBOFFB_30_IV_0L6R_2376\ : AO21
      port map(A => \REGl299r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l6r_adt_net_161946_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161981_\);
    
    \I3.PIPEB_81_2342\ : NOR2FT
      port map(A => \I3.PIPEBl2r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_81_adt_net_160629_\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I153_Y_I_O4_1555\ : AO21
      port map(A => \I2.PIPE4_DTl17r_net_1\, B => 
        \I2.PIPE4_DTl16r_net_1\, C => \I2.RAMDT4L5R_820\, Y => 
        \I2.N_33_adt_net_55021_\);
    
    \I2.L2TYPE_4_IL11R_1622\ : AND2FT
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4467\, Y => \I2.N_4441_adt_net_67338_\);
    
    \I2.DTO_16_1_IVL15R_1143\ : AO21
      port map(A => \I2.N_182_adt_net_1007__net_1\, B => 
        \I2.DT_SRAMl15r_net_1\, C => 
        \I2.DTO_16_1l15r_adt_net_31962_\, Y => 
        \I2.DTO_16_1l15r_adt_net_31963_\);
    
    \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855000_\ : 
        BFR
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__net_1\, Y => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855000__net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_2677\ : AND3
      port map(A => \I2.N_107_adt_net_256839_\, B => 
        \I2.N_128_adt_net_54291_\, C => \I2.N525_adt_net_336000_\, 
        Y => \I2.N525_adt_net_335996_\);
    
    \I1.REG_74_0_IVL292R_1927\ : NOR2FT
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l292r_adt_net_121689_\);
    
    \I3.VDBi_16_m_i_2l3r\ : AND2FT
      port map(A => reg_il0r, B => \I3.N_2053\, Y => 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144601_\);
    
    \I2.PIPE5_DT_6_0l13r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l13r\, B => 
        \I2.un27_pipe5_dt0l13r\, S => 
        \I2.dataout_0_adt_net_855804__net_1\, Y => \I2.N_1082\);
    
    \I2.LSRAM_INl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_406_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl22r_net_1\);
    
    \I2.DTOSl9r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl9r, Q => 
        \I2.DTOSl9r_net_1\);
    
    \I2.DTO_9_iv_ml28r_adt_net_28906_\ : NOR2
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl28r_net_1\, Y => 
        \I2.DTO_9_iv_ml28r_adt_net_28906__net_1\);
    
    \I1.REG_74_0_IVL218R_2016\ : AND2
      port map(A => \FBOUTl5r\, B => \I1.REG_7_sqmuxa\, Y => 
        \I1.REG_74l218r_adt_net_128948_\);
    
    \I2.LSRAM_FL_RD7\ : DFFS
      port map(CLK => CLK_c, D => LSRAM_FL_RD, SET => 
        CLEAR_STAT_i_0, Q => \I2.LSRAM_FL_RD7_net_1\);
    
    \I2.MIC_ERR_REGSl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_334_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl5r_net_1\);
    
    \I2.DTE_21_1_0_IV_0_0L29R_1232\ : AO21FTT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_289\, B => 
        \I2.DT_SRAMl29r_net_1\, C => 
        \I2.DTE_21_1l29r_adt_net_36645_\, Y => 
        \I2.DTE_21_1l29r_adt_net_36650_\);
    
    \I3.STATE1_ns_0_iv_0_a3l4r\ : NOR3FFT
      port map(A => \I3.MBLTCYC_423\, B => \I3.N_90_i_0_1\, C => 
        \I3.N_264_0_adt_net_1653_Rd1__net_1\, Y => \I3.N_1516\);
    
    \I5.SENS_ADDR_6l0r\ : AND2
      port map(A => \I5.SENS_ADDR_1_sqmuxa_net_1\, B => 
        \I5.DWACT_ADD_CI_0_partial_suml0r\, Y => 
        \I5.SENS_ADDR_6l0r_net_1\);
    
    \I3.PIPEAl15r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_246_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl15r_net_1\);
    
    \I3.VDBi_57l2r_adt_net_145304_\ : AO21
      port map(A => \I3.N_2046\, B => \I3.REGl135r\, C => 
        \I3.VDBi_57l2r_adt_net_145303__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145304__net_1\);
    
    \I2.DTO_16_1_IV_0L5R_1197\ : AO21
      port map(A => \I2.DTO_1l5r_net_1\, B => \I2.N_196_52\, C
         => \I2.DTO_16_1l5r_adt_net_34199_\, Y => 
        \I2.DTO_16_1l5r_adt_net_34200_\);
    
    \I3.REG_1_172\ : MUX2L
      port map(A => VDB_inl23r, B => REGl71r, S => 
        \I3.N_1935_adt_net_855320__net_1\, Y => \I3.REG_1_172_0\);
    
    \I2.N475_adt_net_87328_\ : AND2FT
      port map(A => \I2.LSRAM_OUTl18r\, B => 
        \I2.PIPE7_DTl18r_net_1\, Y => 
        \I2.N475_adt_net_87328__net_1\);
    
    \I1.REG_74_i_o2l364r\ : OR2
      port map(A => \I1.N_65_12\, B => \I1.N_661_adt_net_114485_\, 
        Y => \I1.N_661\);
    
    \I2.MIC_ERR_REGSl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_344_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl15r_net_1\);
    
    \I3.REG_1_176\ : MUX2L
      port map(A => VDB_inl27r, B => REGl75r, S => 
        \I3.N_1935_adt_net_855316__net_1\, Y => \I3.REG_1_176_0\);
    
    FBOUTl0r : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_58_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \FBOUTl0r\);
    
    \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_STT_M3_996\ : NOR2
      port map(A => \I3.REG2_144_net_1\, B => \I3.REG3_128_net_1\, 
        Y => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_adt_net_19883_Ra1_\);
    
    \I3.PIPEB_102_2321\ : NOR2FT
      port map(A => \I3.PIPEBl23r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_102_adt_net_159747_\);
    
    \I1.REG_13_sqmuxa_0_a2\ : NOR2
      port map(A => 
        \I1.REG_15_sqmuxa_adt_net_1457__adt_net_854380__net_1\, B
         => \I1.N_255\, Y => \I1.REG_13_sqmuxa\);
    
    \I3.N_264_0_adt_net_1653_Ra1_\ : OR2
      port map(A => \I3.SINGCYC_115_net_1\, B => 
        \I3.BLTCYC_113_net_1\, Y => 
        \I3.N_264_0_adt_net_1653_Ra1__net_1\);
    
    \I2.PIPE5_DT_705\ : MUX2L
      port map(A => \I2.PIPE5_DTl29r_net_1\, B => 
        \I2.PIPE4_DTl29r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_705_net_1\);
    
    \I5.SBYTE_69\ : MUX2H
      port map(A => \I5.SBYTEl4r_net_1\, B => \I5.N_22\, S => 
        \I5.N_406\, Y => \I5.SBYTE_69_net_1\);
    
    \I2.REG_1_c6_i_a2_0\ : AND3FFT
      port map(A => REGL37R_566, B => REGL38R_873, C => 
        \I2.N_124\, Y => \I2.N_126\);
    
    \I2.N_4248_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4248\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4248_Rd1__net_1\);
    
    \I2.RAMAD_4l4r\ : MUX2L
      port map(A => \I2.N_531\, B => \I1.BYTECNT_i_0_il4r_net_1\, 
        S => LOAD_RES, Y => \I2.RAMAD_4l4r_net_1\);
    
    \I2.ADO_3l15r\ : MUX2H
      port map(A => \I2.RPAGEl15r\, B => \I2.WPAGEl15r_net_1\, S
         => NOESRAME_c, Y => \I2.ADO_3l15r_net_1\);
    
    REGl395r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_296_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl395r\);
    
    \I3.VDBi_57_0_iv_0_a2_3l8r\ : AND3FTT
      port map(A => \I3.N_1905_1_adt_net_855376__net_1\, B => 
        \I3.REGMAPl16r_net_1\, C => 
        \I3.N_354_0_adt_net_855372__net_1\, Y => \I3.N_2058\);
    
    \I1.BYTECNT_n6_i_0_o2\ : NOR2FT
      port map(A => \I1.BYTECNTl6r_net_1\, B => \I1.N_335\, Y => 
        \I1.N_358\);
    
    \I2.DTO_1_891\ : MUX2L
      port map(A => \I2.DTO_1l17r_Rd1__net_1\, B => 
        \I2.DTO_16_1l17r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834764_Rd1__net_1\, Y
         => \I2.DTO_1l17r\);
    
    \I2.PIPE5_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_690_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl14r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL21R_1387\ : NOR2FT
      port map(A => REGl425r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, Y => 
        \I2.PIPE1_DT_42l21r_adt_net_46867_\);
    
    \I3.TICKil0r_1451\ : DFFC
      port map(CLK => CLK_c, D => \I3.un6_tcnt1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TICKL0R_558);
    
    \I3.TCNT_n2_0_0_o2_0\ : OR2
      port map(A => \I3.N_1911\, B => \I3.TCNTL2R_430\, Y => 
        \I3.N_1912\);
    
    \I3.TCNTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_381_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTl3r_net_1\);
    
    \I5.REG_1_30\ : MUX2H
      port map(A => \I5.REG_12l431r_net_1\, B => REGl447r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_30_net_1\);
    
    \I3.un1_STATE2_13_adt_net_150841_\ : OR3
      port map(A => \I3.STATE2l1r_net_1\, B => \I3.N_1879\, C => 
        \I3.STATE2l3r_net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_150841__net_1\);
    
    \I3.VAS_69\ : MUX2L
      port map(A => VAD_inl7r, B => \I3.VAS_i_0_il7r\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_69_net_1\);
    
    REGl178r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_79_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl178r\);
    
    \I2.CRC32_823\ : MUX2L
      port map(A => \I2.CRC32l28r_net_1\, B => \I2.N_3945\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_823_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I66_Y\ : AO21
      port map(A => \I2.N252_0\, B => 
        \I2.N316_i_i_adt_net_86582_\, C => 
        \I2.N316_i_i_adt_net_86577_\, Y => \I2.N316_i_i\);
    
    \I2.SUB8_1_sqmuxa_0_adt_net_855144_\ : BFR
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855152__net_1\, Y
         => \I2.SUB8_1_sqmuxa_0_adt_net_855144__net_1\);
    
    \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856_\ : BFR
      port map(A => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855860__net_1\, Y => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\);
    
    \I2.N_140_0_ADT_NET_947__2887\ : OR2
      port map(A => \I2.PIPE4_DTl5r_adt_net_854416__net_1\, B => 
        \I2.PIPE4_DTL6R_854\, Y => \I2.N_140_0_ADT_NET_947__328\);
    
    \I1.REG_74_0_ivl335r\ : AO21
      port map(A => \REGl335r\, B => \I1.N_209\, C => 
        \I1.REG_74l335r_adt_net_117658_\, Y => \I1.REG_74l335r\);
    
    \I3.REGMAPl56r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un227_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPl56r_net_1\);
    
    \I3.VDBI_16_M_I_2L3R_2255\ : OAI21FTF
      port map(A => GA_cl3r, B => \I3.N_2042\, C => 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144610_\, Y => 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144611_\);
    
    \I2.PIPE10_DT_17_i_a3_2l13r\ : OR3
      port map(A => \I2.N_3822_adt_net_64766_\, B => 
        \I2.N_3822_adt_net_64764_\, C => 
        \I2.N_3822_adt_net_64765_\, Y => \I2.N_3822\);
    
    \I2.FID_7_0_ivl25r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl25r_net_1\, 
        C => \I2.FID_7l25r_adt_net_19029_\, Y => \I2.FID_7l25r\);
    
    \I2.EVNT_NUMl0r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_963_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl0r_net_1\);
    
    ADO_padl11r : OB33PH
      port map(PAD => ADO(11), A => ADO_cl11r);
    
    \I3.REGMAP_i_0_il19r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un76_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il19r_net_1\);
    
    \I2.PIPE6_DT_472\ : MUX2H
      port map(A => \I2.PIPE5_DTl18r_net_1\, B => 
        \I2.PIPE6_DTl18r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_472_net_1\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2511\ : AND2
      port map(A => \REGl243r\, B => \I3.REGMAPl27r_net_1\, Y => 
        \I3.N_2070_adt_net_163458_\);
    
    \I5.sstate1se_4_0_0\ : MUX2H
      port map(A => \I5.sstate1l8r_net_1\, B => 
        \I5.sstate1_ns_el5r_adt_net_9070_\, S => TICKl0r, Y => 
        \I5.sstate1_ns_el5r\);
    
    \I2.MIC_REG2_i_0_il4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_313_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2_i_0_il4r_net_1\);
    
    \I1.REG_74_0_ivl178r\ : AO21
      port map(A => \REGl178r\, B => \I1.N_49\, C => 
        \I1.REG_74l178r_adt_net_132510_\, Y => \I1.REG_74l178r\);
    
    \I3.REGMAPl9r_adt_net_854328_\ : BFR
      port map(A => \I3.REGMAPl9r_adt_net_854332__net_1\, Y => 
        \I3.REGMAPl9r_adt_net_854328__net_1\);
    
    \I2.PIPE2_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl15r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl15r_net_1\);
    
    \I2.PIPE1_DT_42_1_iv_0l24r\ : OAI21TTF
      port map(A => REGl444r, B => 
        \I2.N_3234_adt_net_855648__net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_0_il24r_adt_net_46513_\, Y => 
        \I2.PIPE1_DT_42_1_iv_0_il24r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I122_Y_0\ : OAI21
      port map(A => \I2.N_107_adt_net_276024_\, B => \I2.N394\, C
         => \I2.N_64\, Y => \I2.N537_i\);
    
    \I2.PIPE9_DT_293\ : MUX2L
      port map(A => \I2.PIPE9_DTl24r_net_1\, B => 
        \I2.PIPE8_DTl24r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_293_net_1\);
    
    \I2.OFFSET_37_11l4r\ : MUX2L
      port map(A => \REGl377r\, B => \REGl313r\, S => 
        \I2.PIPE7_DTL27R_80\, Y => \I2.N_719\);
    
    \I2.MIC_ERR_REGSl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_335_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl6r_net_1\);
    
    \I1.PAGECNT_320\ : MUX2H
      port map(A => \I1.PAGECNTl7r_net_1\, B => \I1.N_1378\, S
         => \I1.PAGECNTe_adt_net_854892__net_1\, Y => 
        \I1.PAGECNT_320_net_1\);
    
    \I2.L2TYPEl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_600_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl11r_net_1\);
    
    \I1.REG_74_0_ivl266r\ : AO21
      port map(A => \REGl266r\, B => 
        \I1.N_137_adt_net_854760__net_1\, C => 
        \I1.REG_74l266r_adt_net_124199_\, Y => \I1.REG_74l266r\);
    
    \I5.TEMP_ACK_73\ : MUX2L
      port map(A => \I5.TEMP_ACK_net_1\, B => REGl118r, S => 
        \I5.N_443\, Y => \I5.TEMP_ACK_73_net_1\);
    
    \I3.REG_44_IL89R_2302\ : AOI21FTT
      port map(A => REGl89r, B => \I3.N_98_0\, C => \I3.N_1673\, 
        Y => \I3.N_1635_adt_net_150153_\);
    
    \I2.RAMADl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l3r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl3r);
    
    \I2.MIC_ERR_REGS_337\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl9r_net_1\, B => 
        \I2.MIC_ERR_REGSl8r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_337_net_1\);
    
    \I2.FID_7_0_ivl27r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl27r_net_1\, 
        C => \I2.FID_7l27r_adt_net_18841_\, Y => \I2.FID_7l27r\);
    
    \I2.CRC32l8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_803_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l8r_net_1\);
    
    \I2.EVNT_NUM_963\ : MUX2L
      port map(A => \I2.EVNT_NUMl0r_net_1\, B => 
        \I2.EVNT_NUM_n0_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_963_net_1\);
    
    \I2.DTESl13r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl13r, Q => 
        \I2.DTESl13r_net_1\);
    
    \I3.REG_1l88r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_269_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl88r);
    
    \I2.RESYN_0_I2_TRGCNT_C2_I_941\ : AOI21
      port map(A => \I2.TRGCNTl2r_net_1\, B => \I2.N_3765\, C => 
        \I2.un9_tdctrgi_i_0\, Y => \I2.N_3763_adt_net_16097_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_1005\ : OR2FT
      port map(A => \I2.N_45_0\, B => \I2.N525_adt_net_57834_\, Y
         => \I2.N525_383\);
    
    \I5.AIR_WDATA_56\ : MUX2H
      port map(A => \I5.sstate2l3r_net_1\, B => 
        \I5.AIR_WDATAl1r_net_1\, S => \I5.N_461\, Y => 
        \I5.AIR_WDATA_56_net_1\);
    
    REGl236r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_137_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl236r\);
    
    \I5.COMMANDl1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_13_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl1r_net_1\);
    
    \I2.PIPE5_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_693_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl17r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I109_Y_0\ : AO21
      port map(A => \I2.N288\, B => \I2.N291\, C => \I2.N287\, Y
         => \I2.ADD_18x18_fast_I109_Y_0\);
    
    \I2.G_EVNT_NUM_934\ : MUX2L
      port map(A => \I2.G_EVNT_NUM_i_0_il0r_net_1\, B => 
        \I2.G_EVNT_NUM_n0\, S => \I2.N_3769\, Y => 
        \I2.G_EVNT_NUM_934_net_1\);
    
    \I1.LUT_0_sqmuxa_i_0_o2_i_0\ : NOR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__186\, B
         => \I1.N_325\, Y => \I1.N_328_i_0\);
    
    \I1.BYTECNTlde_i_a2_i_845\ : AO21
      port map(A => \I1.N_628\, B => 
        \I1.sstate_ns_i_0_a4_0_1l0r_adt_net_107171_\, C => 
        \I1.N_223_226\, Y => \I1.N_1383_223\);
    
    \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112_\ : BFR
      port map(A => \I2.un3_tdcgda1_1_adt_net_821__net_1\, Y => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\);
    
    \I2.WOFFSETl4r_adt_net_854980_\ : BFR
      port map(A => \I2.WOFFSETl4r\, Y => 
        \I2.WOFFSETl4r_adt_net_854980__net_1\);
    
    \I1.PAGECNT_0l8r_adt_net_834720__adt_net_835724_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_319_adt_net_854860__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0l8r_adt_net_834720__adt_net_835724_Rd1__net_1\);
    
    \I1.REG_74_0_ivl397r\ : AO21
      port map(A => \REGl397r\, B => \I1.N_273\, C => 
        \I1.REG_74l397r_adt_net_110358_\, Y => \I1.REG_74l397r\);
    
    \I2.OFFSET_37_4l0r\ : MUX2L
      port map(A => \REGl365r\, B => \REGl301r\, S => 
        \I2.PIPE7_DTL27R_74\, Y => \I2.N_659\);
    
    \I3.PIPEA_8_0l13r\ : MUX2L
      port map(A => DPR_cl13r, B => \I3.PIPEA1l13r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855348__net_1\, Y => \I3.N_222\);
    
    \I1.N_50_0_ADT_NET_109751__2862\ : NOR3FFT
      port map(A => \I1.N_232_1_296\, B => 
        \I1.N_50_0_adt_net_109760__net_1\, C => \I1.N_435_1_284\, 
        Y => \I1.N_50_0_ADT_NET_109751__257\);
    
    \I2.PIPE1_DT_42_i_0l15r\ : OR2FT
      port map(A => \I2.N_3283_adt_net_855064__net_1\, B => 
        \I2.N_3238_adt_net_48555_\, Y => \I2.N_3238\);
    
    \I1.REG_74_0_ivl318r\ : AO21
      port map(A => \REGl318r\, B => \I1.N_193\, C => 
        \I1.REG_74l318r_adt_net_119217_\, Y => \I1.REG_74l318r\);
    
    \I3.UN1_STATE2_11_0_0_2309\ : AO21
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, B => 
        \I3.un1_STATE2_11_adt_net_1401__net_1\, C => 
        \I3.STATE2l4r_net_1\, Y => 
        \I3.un1_STATE2_11_adt_net_153728_\);
    
    \I2.PIPE3_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl19r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl19r_net_1\);
    
    \I2.N_140_0_adt_net_947_\ : OR2
      port map(A => \I2.PIPE4_DTl5r_adt_net_854420__net_1\, B => 
        \I2.PIPE4_DTL6R_479\, Y => 
        \I2.N_140_0_adt_net_947__net_1\);
    
    \I1.REG_74_0_ivl240r\ : AO21
      port map(A => \REGl240r\, B => \I1.N_113\, C => 
        \I1.REG_74l240r_adt_net_126727_\, Y => \I1.REG_74l240r\);
    
    \I2.DTOSl1r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl1r, Q => 
        \I2.DTOSl1r_net_1\);
    
    \I2.DTO_16_1_iv_0l31r\ : OR2
      port map(A => \I2.DTO_16_1l31r_adt_net_28255_\, B => 
        \I2.DTO_16_1l31r_adt_net_28256_\, Y => \I2.DTO_16_1l31r\);
    
    \I2.DTO_16_1_iv_0l27r\ : OR2
      port map(A => \I2.DTO_16_1l27r_adt_net_29251_\, B => 
        \I2.DTO_16_1l27r_adt_net_29252_\, Y => \I2.DTO_16_1l27r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_o2_727\ : AND3FFT
      port map(A => \I2.N_3_0_adt_net_1070__net_1\, B => 
        \I2.N_95_0\, C => \I2.N_45_1_adt_net_271427_\, Y => 
        \I2.N_45_1_105\);
    
    \I2.DT_TEMP_7l14r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854244__net_1\, B => 
        \I2.DT_SRAMl14r_net_1\, Y => \I2.DT_TEMP_7l14r_net_1\);
    
    \I1.un1_sbyte13_2_i_i_a2_i_849\ : OR2FT
      port map(A => \I1.N_436_i_i\, B => 
        \I1.N_223_adt_net_108707_\, Y => \I1.N_223_227\);
    
    \I1.REG_74_1_380_M8_I_0_RD1__2893\ : DFFC
      port map(CLK => CLK_c, D => \I1.REG_74_1_380_m8_i_0_Ra1_\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.REG_74_1_380_M8_I_0_RD1__336\);
    
    \I2.G_EVNT_NUM_n11_0_a2\ : NAND3FFT
      port map(A => EV_RES_C_568, B => \I2.N_287_adt_net_26828_\, 
        C => \I2.G_EVNT_NUMl11r_net_1\, Y => \I2.N_287\);
    
    \I2.CRC32l6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_801_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l6r_net_1\);
    
    \I2.un78_pipe5_dt\ : XOR2
      port map(A => \I2.RAMDT4l12r_net_1\, B => 
        \I2.un78_pipe5_dt_4_net_1\, Y => \I2.dataout_1\);
    
    RAMDT_padl5r : IOB33PH
      port map(PAD => RAMDT(5), A => \I1.RAMDT_SPI_1l5r_net_1\, 
        EN => \I1.RAMDT_SPI_e_net_1\, Y => RAMDT_inl5r);
    
    \I2.DT_TEMP_7l13r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854244__net_1\, B => 
        \I2.N_4048\, Y => \I2.DT_TEMP_7l13r_net_1\);
    
    REGl293r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_194_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl293r\);
    
    \I2.N_70_adt_net_255801_\ : OR2FT
      port map(A => \I2.N_95\, B => 
        \I2.N_70_adt_net_54406__net_1\, Y => 
        \I2.N_70_adt_net_255801__net_1\);
    
    \I3.REG_1l164r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_212_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl164r\);
    
    \I2.RAMDT4L12R_3072\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_826\);
    
    \I2.PIPE1_DT_42_1_IVL30R_1354\ : AO21FTT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        B => \I2.PIPE1_DT_12l30r_net_1\, C => 
        \I2.PIPE1_DT_42l30r_adt_net_45594_\, Y => 
        \I2.PIPE1_DT_42l30r_adt_net_45595_\);
    
    \I3.VDBi_16_m_i_o3l3r_888\ : OR2
      port map(A => \I3.REGMAPL8R_740\, B => \I3.REGMAPL9R_786\, 
        Y => \I3.N_1907_266\);
    
    \I2.DTESl28r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl28r, Q => 
        \I2.DTESl28r_net_1\);
    
    \I2.CRC32_12_il24r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_128_i_0_i_0\, Y => 
        \I2.N_3941\);
    
    \I3.PIPEBl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_82_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl3r_net_1\);
    
    \I1.REG_74_0_IVL384R_1809\ : AND2
      port map(A => \FBOUTl3r\, B => \I1.REG_28_sqmuxa\, Y => 
        \I1.REG_74l384r_adt_net_111663_\);
    
    \I3.VDBml0r\ : MUX2L
      port map(A => \I3.VDBil0r_net_1\, B => \I3.N_142\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml0r_net_1\);
    
    \I3.REGMAPl8r_1632\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un37_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL8R_739\);
    
    \I2.PIPE5_DT_6l0r\ : MUX2L
      port map(A => \I2.PIPE4_DTl0r_net_1\, B => \I2.N_1069\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, Y
         => \I2.PIPE5_DT_6l0r_net_1\);
    
    \I2.DTO_16_1_iv_0_o2_0l12r\ : AO21FTT
      port map(A => \I2.N_4283_i_0_adt_net_854968__net_1\, B => 
        \I2.DT_TEMPl12r_net_1\, C => \I2.N_3966_adt_net_32562_\, 
        Y => \I2.N_3966\);
    
    \I3.VDBi_29l3r\ : NOR3
      port map(A => \I3.REGMAPL14R_734\, B => 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144601_\, C => 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144611_\, Y => 
        \I3.VDBi_29l3r_adt_net_510711_\);
    
    \I3.VDBoffl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_120_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl4r_net_1\);
    
    \I3.CYCSF1\ : DFFC
      port map(CLK => CLK_c, D => \I3.CYCSF1_60_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.CYCSF1_net_1\);
    
    \I2.PIPE8_DT_552\ : MUX2L
      port map(A => \I2.PIPE8_DTl24r_net_1\, B => 
        \I2.PIPE8_DT_21l24r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_552_net_1\);
    
    \I1.REG_74_0_ivl270r\ : AO21
      port map(A => \REGl270r\, B => 
        \I1.N_145_adt_net_854768__net_1\, C => 
        \I1.REG_74l270r_adt_net_123818_\, Y => \I1.REG_74l270r\);
    
    \I5.BITCNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.BITCNT_85_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.BITCNTl1r_net_1\);
    
    \I2.DTESl24r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl24r, Q => 
        \I2.DTESl24r_net_1\);
    
    \I5.DATA_12l10r\ : MUX2L
      port map(A => REGl127r, B => \I5.SBYTEl2r_net_1\, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l10r_net_1\);
    
    \I2.DT_TEMPl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_775_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl14r_net_1\);
    
    \I1.REG_0_sqmuxa_i_0_o2_0\ : AND3FFT
      port map(A => \I1.BYTECNT_307_net_1\, B => 
        \I1.BYTECNT_308_net_1\, C => 
        \I1.N_304_adt_net_105325_Ra1_\, Y => \I1.N_304_Ra1_\);
    
    REGl276r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_177_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl276r\);
    
    \I3.PIPEAl7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_238_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl7r_net_1\);
    
    \I3.un10_tcnt2\ : OR3FTT
      port map(A => \I3.un6_tcnt1_net_1\, B => 
        \I3.un10_tcnt2_adt_net_135290_\, C => 
        \I3.un10_tcnt2_adt_net_135291_\, Y => 
        \I3.un10_tcnt2_net_1\);
    
    \I1.REG_74_0_IVL380R_1819\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l380r_adt_net_112485_\);
    
    REGl285r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_186_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl285r\);
    
    REGl288r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_189_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl288r\);
    
    \I1.REG_74_0_IVL298R_1920\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l298r_adt_net_121040_\);
    
    \I3.VDBi_16_m_i_m2l12r\ : MUX2H
      port map(A => REGl28r, B => REGl44r, S => 
        \I3.REGMAPl7r_net_1\, Y => \I3.N_280\);
    
    \I2.UN1_DTO_CL_0_SQMUXA_0_0_O2_1_1021\ : AO21TTF
      port map(A => \I2.STATE2l5r_net_1\, B => \I2.N_237\, C => 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, Y => 
        \I2.un1_DTO_cl_0_sqmuxa_adt_net_22686_\);
    
    \I2.OFFSET_37_15l5r\ : MUX2L
      port map(A => \REGl234r\, B => \REGl170r\, S => 
        \I2.PIPE7_DTL27R_69\, Y => \I2.N_752\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I10_G0N_0_o2\ : NAND2
      port map(A => \I2.RAMDT4L5R_818\, B => 
        \I2.PIPE4_DTL10R_792\, Y => \I2.N_66\);
    
    \I2.EVNT_WORD_715\ : MUX2H
      port map(A => \I2.EVNT_WORDl2r_net_1\, B => \I2.I_9_0\, S
         => \I2.N_2864_0_adt_net_854276__net_1\, Y => 
        \I2.EVNT_WORD_715_net_1\);
    
    \I2.PIPE6_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_471_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl17r_net_1\);
    
    \I2.TOKENA_CNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TOKENA_CNT_4l0r_net_1\, CLR
         => \I2.un6_clear_stat_i\, Q => \I2.TOKENA_CNTl0r_net_1\);
    
    RAMAD_padl3r : OB33PH
      port map(PAD => RAMAD(3), A => RAMAD_cl3r);
    
    \I3.TCNT_n4_0_0\ : OAI21
      port map(A => \I3.un1_STATE1_10_i_0\, B => \I3.N_263_i\, C
         => \I3.N_1966_1\, Y => \I3.TCNT_n4\);
    
    \I5.un1_sdaa_0_a2\ : NOR2
      port map(A => \I5.CHAIN_SELECT_net_1\, B => 
        \I5.SDAnoe_net_1\, Y => un1_sdaa_0_a2);
    
    \I2.ROFFSET_911\ : MUX2H
      port map(A => \I2.ROFFSETl7r_net_1\, B => 
        \I2.ROFFSET_n7_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_911_net_1\);
    
    \I1.PAGECNTlde_0\ : OR2
      port map(A => \I1.N_292\, B => 
        \I1.PAGECNTe_adt_net_106660_\, Y => \I1.PAGECNTe\);
    
    \I2.END_EVNT1_710\ : OA21TTF
      port map(A => \I2.N_3798\, B => \I2.END_EVNT1_net_1\, C => 
        \I2.STATE1l17r_net_1\, Y => \I2.END_EVNT1_710_net_1\);
    
    \I2.DTE_21_1_ivl23r\ : AO21
      port map(A => \I2.DTE_1l23r_Rd1__net_1\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835168_Rd1__net_1\, 
        C => \I2.DTE_21_1l23r_adt_net_37285_Rd1__net_1\, Y => 
        \I2.DTE_21_1l23r_Rd1_\);
    
    \I2.DT_TEMP_763\ : MUX2H
      port map(A => \I2.DT_TEMPl2r_net_1\, B => 
        \I2.DT_TEMP_7l2r_net_1\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.DT_TEMP_763_net_1\);
    
    \I2.WPAGE_n1\ : XOR2
      port map(A => \I2.WPAGEl13r_net_1\, B => 
        \I2.WPAGEl12r_net_1\, Y => \I2.WPAGE_n1_net_1\);
    
    \I3.VDBOFFB_30_IV_0L6R_2377\ : AO21
      port map(A => \REGl347r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        C => \I3.VDBoffb_30l6r_adt_net_161950_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161982_\);
    
    \I2.RAMDT4L12R_2818\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_146\);
    
    \I2.MIC_REG3_320\ : MUX2H
      port map(A => \I2.MIC_REG3l3r_net_1\, B => 
        \I2.MIC_REG3l4r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_net_1\, Y => 
        \I2.MIC_REG3_320_net_1\);
    
    \I2.ADEl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl3r);
    
    \I2.FIDl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_417_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl1r);
    
    \I2.PIPE8_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_530_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl2r_net_1\);
    
    \I2.L2ARR_c2\ : NOR2FT
      port map(A => \I2.L2ARRl2r_net_1\, B => \I2.N_4454\, Y => 
        \I2.L2ARR_c2_net_1\);
    
    \I2.DTE_21_1_iv_0l13r\ : OR3
      port map(A => \I2.DTE_21_1l13r_adt_net_38171_\, B => 
        \I2.DTE_21_1l13r_adt_net_38179_\, C => 
        \I2.DTE_21_1l13r_adt_net_38180_\, Y => \I2.DTE_21_1l13r\);
    
    \I3.VDBi_31l3r\ : MUX2L
      port map(A => \I3.REGl136r\, B => \I3.VDBi_29l3r_net_1\, S
         => \I3.REGMAPl17r_adt_net_854292__net_1\, Y => 
        \I3.VDBi_31l3r_net_1\);
    
    \I3.VDBI_57_IV_0L5R_2245\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854360__net_1\, B
         => \I3.VDBoffl5r_net_1\, Y => 
        \I3.VDBi_57l5r_adt_net_143850_\);
    
    \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072_\ : BFR
      port map(A => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855076__net_1\, Y
         => \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\);
    
    \I2.PIPE1_DT_42_1_IVL10R_1465\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\, B => 
        \I2.PIPE1_DT_30l10r_net_1\, C => 
        \I2.PIPE1_DT_42l10r_adt_net_49936_\, Y => 
        \I2.PIPE1_DT_42l10r_adt_net_49952_\);
    
    \I3.REG_1_187\ : MUX2L
      port map(A => VDB_inl6r, B => \I3.REGl139r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, Y => 
        \I3.REG_1_187_0\);
    
    \I3.PIPEAl9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_240_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl9r_net_1\);
    
    \I1.REG_74_0_ivl294r\ : AO21
      port map(A => \REGl294r\, B => \I1.N_169\, C => 
        \I1.REG_74l294r_adt_net_121384_\, Y => \I1.REG_74l294r\);
    
    \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096_\ : BFR
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855104__net_1\, Y
         => \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096__net_1\);
    
    \I1.REG_74l220r\ : OR3
      port map(A => \I1.N_89_adt_net_128732_\, B => 
        \I1.N_97_6_adt_net_854712__net_1\, C => 
        \I1.N_89_adt_net_128736_\, Y => \I1.N_89\);
    
    DTE_padl7r : IOB33PH
      port map(PAD => DTE(7), A => \I2.DTE_1l7r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl7r);
    
    REGl199r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_100_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl199r\);
    
    \I3.PULSE_338\ : MUX2L
      port map(A => PULSEl8r, B => \I3.PULSE_46l8r\, S => 
        \I3.N_1409_adt_net_854740__net_1\, Y => 
        \I3.PULSE_338_net_1\);
    
    \I2.DTE_21_1_IVL23R_1251\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l23r\, C
         => \I2.DTE_21_1l23r_adt_net_37284_\, Y => 
        \I2.DTE_21_1l23r_adt_net_37285_\);
    
    \I1.REG_1_124\ : MUX2H
      port map(A => \REGl223r\, B => \I1.REG_74l223r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\, Y => 
        \I1.REG_1_124_net_1\);
    
    \I1.BYTECNT_n8_i_0_x2\ : XOR2
      port map(A => \I1.BYTECNTl8r_net_1\, B => \I1.N_363\, Y => 
        \I1.N_413_i_0\);
    
    \I3.N_1186_adt_net_1488_\ : OR2
      port map(A => \I3.STATE1_IPL2R_886\, B => \I3.N_1180\, Y
         => \I3.N_1186_adt_net_1488__net_1\);
    
    \I2.OFFSET_37_21l4r\ : MUX2L
      port map(A => \I2.N_791\, B => \I2.N_767\, S => 
        \I2.PIPE7_DTL25R_685\, Y => \I2.N_799\);
    
    \I3.VDBil17r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_357_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil17r_net_1\);
    
    \I5.REG_1l422r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_35_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl422r);
    
    \PULSEl0r_adt_net_854532__adt_net_855544_\ : BFR
      port map(A => \PULSEl0r_adt_net_854532__net_1\, Y => 
        \PULSEl0r_adt_net_854532__adt_net_855544__net_1\);
    
    \I3.VDBi_57_iv_0_0_a2_10l7r_939\ : OR2FT
      port map(A => \I3.N_2016_319\, B => \I3.REGMAPL14R_733\, Y
         => \I3.N_2017_317\);
    
    \I2.OFFSET_37_3l5r\ : MUX2L
      port map(A => \I2.N_648\, B => \I2.N_640\, S => 
        \I2.PIPE7_DTL26R_349\, Y => \I2.N_656\);
    
    \I3.PIPEB_100\ : AO21
      port map(A => DPR_cl21r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\, 
        C => \I3.PIPEB_100_adt_net_159831_\, Y => 
        \I3.PIPEB_100_net_1\);
    
    \I2.OFFSETl7r_1563\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_567_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL7R_670\);
    
    \I2.L2SERVl3r_1255\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_517\);
    
    \I1.ISI_7_i_0\ : AND2
      port map(A => \I1.N_1193_adt_net_1562__net_1\, B => 
        \I1.N_1193_adt_net_134015_\, Y => \I1.N_1193\);
    
    \I2.DTE_21_1_IV_0L20R_1258\ : AND2FT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855200__net_1\, 
        B => \I2.DT_TEMPl20r_net_1\, Y => 
        \I2.DTE_21_1l20r_adt_net_37603_\);
    
    \I3.TCNT3_377\ : MUX2H
      port map(A => \I3.TCNT3_i_0_il2r_net_1\, B => 
        \I3.TCNT3_n2_net_1\, S => \TICKl1r\, Y => 
        \I3.TCNT3_377_net_1\);
    
    \I2.PIPE8_DT_528\ : MUX2L
      port map(A => \I2.PIPE8_DTl0r_net_1\, B => 
        \I2.PIPE8_DT_21l0r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_528_net_1\);
    
    \I2.DTE_0_sqmuxa_i_o2tt_N_8_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.DTE_0_sqmuxa_i_o2tt_N_8_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.DTE_0_sqmuxa_i_o2tt_N_8_Rd1__net_1\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854480_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854492__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854480__net_1\);
    
    \I2.DT_TEMP_765\ : MUX2H
      port map(A => \I2.DT_TEMPl4r_net_1\, B => 
        \I2.DT_TEMP_7l4r_net_1\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.DT_TEMP_765_net_1\);
    
    \I2.L2TYPEl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_604_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl15r_net_1\);
    
    N_1_I3_TCNT2_c3 : AND2
      port map(A => \I3.TCNT2l3r_net_1\, B => \I3.TCNT2_c2\, Y
         => \I3.TCNT2_c3\);
    
    \I3.VDBOFFA_31_IV_0L5R_2545\ : OR3
      port map(A => \I3.VDBoffa_31l5r_adt_net_163697_\, B => 
        \I3.VDBoffa_31l5r_adt_net_163693_\, C => 
        \I3.VDBoffa_31l5r_adt_net_163694_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163700_\);
    
    \I1.REG_74_0_ivl333r\ : AO21
      port map(A => \REGl333r\, B => \I1.N_209\, C => 
        \I1.REG_74l333r_adt_net_117830_\, Y => \I1.REG_74l333r\);
    
    \I5.REG_1_35\ : MUX2L
      port map(A => \I5.TEMPDATAl2r_net_1\, B => REGl422r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_35_net_1\);
    
    \I3.PIPEA1_316\ : MUX2L
      port map(A => \I3.PIPEA1l18r_net_1\, B => 
        \I3.PIPEA1_12l18r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__252\, Y => 
        \I3.PIPEA1_316_net_1\);
    
    \I2.OFFSETl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_561_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl1r_net_1\);
    
    \I1.BYTECNT_n8_i_0\ : NOR2
      port map(A => \I1.N_223_adt_net_854844__net_1\, B => 
        \I1.N_413_i_0\, Y => \I1.N_1162\);
    
    F_SCK_c : DFFC
      port map(CLK => CLK_c, D => \I1.ISCK_53_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \F_SCK_c\);
    
    \I2.MIC_REG2l3r_adt_net_834020_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.MIC_REG2_312_adt_net_855644__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2l3r_adt_net_834020_Rd1__net_1\);
    
    \I2.PIPE8_DT_16_0l6r\ : MUX2H
      port map(A => \I2.PIPE8_DTl6r_net_1\, B => 
        \I2.PIPE7_DTl6r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_572\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__2763\ : NAND3FFT
      port map(A => \I2.ENDF_837\, B => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__236\, C => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_net_1\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__46\);
    
    TDCDB_padl6r : IB33
      port map(PAD => TDCDB(6), Y => TDCDB_cl6r);
    
    \I2.WOFFSET_835\ : MUX2L
      port map(A => \I2.WOFFSETl8r_Rd1__net_1\, B => 
        \I2.N_4251_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835308_Rd1__net_1\, Y
         => \I2.WOFFSETl8r\);
    
    \I3.TCNT1_c4\ : NAND2
      port map(A => \I3.TCNT1l4r_net_1\, B => \I3.TCNT1_c3_net_1\, 
        Y => \I3.TCNT1_c4_net_1\);
    
    \I2.DTO_16_1_IV_0_0L12R_1160\ : AO21
      port map(A => \I2.N_457\, B => \I2.N_93_i_0\, C => 
        \I2.DTO_16_1l12r_adt_net_32624_\, Y => 
        \I2.DTO_16_1l12r_adt_net_32633_\);
    
    \I1.REG_74_0_ivl311r\ : AO21
      port map(A => \REGl311r\, B => \I1.N_185\, C => 
        \I1.REG_74l311r_adt_net_119819_\, Y => \I1.REG_74l311r\);
    
    \I3.VDBOFFB_30_IV_0L2R_2448\ : AO21
      port map(A => \REGl295r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l2r_adt_net_162706_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162741_\);
    
    \I2.DT_SRAMl8r\ : MUX2L
      port map(A => \I2.N_876\, B => \I2.PIPE2_DTl8r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672__net_1\, 
        Y => \I2.DT_SRAMl8r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I144_Y\ : AND2
      port map(A => \I2.N319_0\, B => \I2.N323_0\, Y => 
        \I2.N510_adt_net_220872_\);
    
    \I3.VDBOFFA_31_IV_0L7R_2494\ : AND2
      port map(A => \REGl204r\, B => \I3.REGMAPl22r_net_1\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163272_\);
    
    \I3.VDBOFFA_31_IV_0L3R_2577\ : AO21
      port map(A => \REGl168r\, B => \I3.REGMAPl18r_net_1\, C => 
        \I3.VDBoffa_31l3r_adt_net_164048_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164074_\);
    
    \I2.PIPE2_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl18r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl18r_net_1\);
    
    \I3.un126_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.N_641\, B => \I3.N_553\, Y => 
        \I3.un126_reg_ads_0_a2_1_a3_net_1\);
    
    \I3.N_57_i_0_0_adt_net_854688_\ : BFR
      port map(A => \I3.N_57_i_0_0\, Y => 
        \I3.N_57_i_0_0_adt_net_854688__net_1\);
    
    \I2.PIPE8_DT_16l15r\ : AND2
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\, B => 
        \I2.N_581\, Y => \I2.PIPE8_DT_16l15r_net_1\);
    
    \I2.PIPE10_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_610_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl5r_net_1\);
    
    \I1.BYTECNTlde_i_a2_i_o2_1\ : NAND3FTT
      port map(A => \I1.BYTECNT_311_net_1\, B => 
        \I1.BYTECNT_312_net_1\, C => \I1.BYTECNT_313_net_1\, Y
         => \I1.N_333_Ra1_\);
    
    \I3.STATE1_NS_0_IV_0L1R_2078\ : NOR3FFT
      port map(A => \I3.N_268\, B => \I3.STATE1l10r_net_1\, C => 
        \I3.DSS_net_1\, Y => \I3.STATE1_nsl1r_adt_net_134332_\);
    
    \I2.PIPE5_DT_6l12r\ : MUX2L
      port map(A => \I2.PIPE4_DTl12r_net_1\, B => \I2.N_1081\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\, Y
         => \I2.PIPE5_DT_6l12r_net_1\);
    
    \I2.MIC_ERR_REGSl41r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_370_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl41r_net_1\);
    
    \I4.RESYN_0_I4_UN1_BCNT_2_928\ : OR2
      port map(A => \I4.bcnt_i_0_il2r_net_1\, B => 
        \I4.bcntl1r_net_1\, Y => \I4.N_48_3_adt_net_14719_\);
    
    \I3.STATE1l8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl2r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL8R_10\);
    
    \I2.MIC_REG2l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_309_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2l0r_net_1\);
    
    \I1.REG_74_0_IVL177R_2057\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, Y => 
        \I1.REG_74l177r_adt_net_132596_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I4_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L4R_764\, B => \I2.PIPE4_DTL4R_852\, 
        Y => \I2.N_64\);
    
    \I2.DTE_21_1_IV_0L20R_1260\ : OAI21FTF
      port map(A => \I2.STATE2l1r_adt_net_855128__net_1\, B => 
        \I2.N_3283\, C => \I2.DTE_21_1l20r_adt_net_37603_\, Y => 
        \I2.DTE_21_1l20r_adt_net_37612_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I173_Y\ : XOR2
      port map(A => \I2.N_2358_tz_tz_adt_net_854952__net_1\, B
         => \I2.ADD_21x21_fast_I173_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l3r\);
    
    \I2.MIC_ERR_REGSl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_351_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl22r_net_1\);
    
    \I2.G_EVNT_NUMl2r_955\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_932_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUML2R_333\);
    
    \I3.VDBOFFA_31_IV_0L3R_2579\ : OR2
      port map(A => \I3.VDBoffa_31l3r_adt_net_164071_\, B => 
        \I3.VDBoffa_31l3r_adt_net_164072_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164077_\);
    
    \I2.N_4283_i_0_a2_m1_e_0_856\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__46\, B => 
        \I2.TEMPF_adt_net_855744__net_1\, Y => 
        \I2.N_4283_I_0_234\);
    
    \I2.PIPE10_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_612_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl7r_net_1\);
    
    \I2.OFFSET_37_19l5r\ : MUX2L
      port map(A => \REGl282r\, B => \REGl218r\, S => 
        \I2.PIPE7_DTL27R_88\, Y => \I2.N_784\);
    
    \I1.REG_74_0_IVL288R_1931\ : NOR2FT
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l288r_adt_net_122033_\);
    
    \I1.REG_74_0_ivl292r\ : AO21
      port map(A => \REGl292r\, B => \I1.N_161\, C => 
        \I1.REG_74l292r_adt_net_121689_\, Y => 
        \I1.REG_74l292r_net_1\);
    
    \I2.STATE3_ns_il7r\ : AND2
      port map(A => \I2.STATE3L7R_391\, B => PULSEl3r, Y => 
        \I2.STATE3_ns_il7r_net_1\);
    
    \I3.PIPEA1_321\ : MUX2L
      port map(A => \I3.PIPEA1l23r_net_1\, B => 
        \I3.PIPEA1_12l23r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__251\, Y => 
        \I3.PIPEA1_321_net_1\);
    
    \I2.DTE_2_1_0l4r\ : XOR2
      port map(A => \I2.CRC32l12r_net_1\, B => 
        \I2.CRC32l0r_net_1\, Y => \I2.DTE_2_1_0l4r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I36_Y\ : AND2FT
      port map(A => \I2.SUB8l11r_adt_net_855580__net_1\, B => 
        \I2.N301_1_adt_net_70232_\, Y => \I2.N301_1\);
    
    \I2.EVNT_WORD_719\ : MUX2H
      port map(A => \I2.EVNT_WORDl6r_net_1\, B => \I2.I_31\, S
         => \I2.N_2864_0_adt_net_854272__net_1\, Y => 
        \I2.EVNT_WORD_719_net_1\);
    
    \I3.REG_1_216\ : MUX2L
      port map(A => VDB_inl3r, B => REGl409r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_216_0\);
    
    \I3.VDBi_29l1r\ : MUX2L
      port map(A => \I3.REGl92r\, B => 
        \I3.VDBi_23l1r_adt_net_145581_\, S => \I3.REGMAPL14R_734\, 
        Y => \I3.VDBi_29l1r_adt_net_411517_\);
    
    \I3.REG_44_il89r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_1635_adt_net_150153_\, Y => \I3.N_1635\);
    
    \I2.DT_TEMP_7l17r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854240__net_1\, B => 
        \I2.N_188\, Y => \I2.DT_TEMP_7l17r_net_1\);
    
    \I2.PIPE5_DT_681\ : MUX2L
      port map(A => \I2.PIPE5_DTl5r_net_1\, B => 
        \I2.PIPE5_DT_6l5r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_681_net_1\);
    
    \I2.RAMDT4L4R_3010\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl4r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L4R_764\);
    
    \I1.REG_1_172\ : MUX2H
      port map(A => \REGl271r\, B => \I1.REG_74l271r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y => 
        \I1.REG_1_172_net_1\);
    
    \I5.DATAl11r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l11r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl128r);
    
    \I2.PIPE7_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl24r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl24r_net_1\);
    
    \I2.ROFFSET_n2\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855700__net_1\, B => 
        \I2.ROFFSET_n2_tz_i\, Y => \I2.ROFFSET_n2_net_1\);
    
    \I2.CRC32l18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_813_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l18r_net_1\);
    
    \I2.PIPE5_DT_6_dl20r\ : MUX2L
      port map(A => \I2.PIPE4_DTl20r_net_1\, B => 
        \I2.un27_pipe5_dt1l20r\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855616__net_1\, Y => 
        \I2.PIPE5_DT_6_dl20r_net_1\);
    
    \I1.REG_1_240\ : MUX2H
      port map(A => \REGl339r\, B => \I1.REG_74l339r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\, Y => 
        \I1.REG_1_240_net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__2994\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__541\);
    
    \I3.STATE1_ipl3r_adt_net_854368_\ : BFR
      port map(A => \I3.STATE1_ipl3r_net_1\, Y => 
        \I3.STATE1_ipl3r_adt_net_854368__net_1\);
    
    \I2.LSRAM_IN_389\ : MUX2L
      port map(A => \I2.PIPE5_DTl5r_net_1\, B => 
        \I2.LSRAM_INl5r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_389_net_1\);
    
    \I4.resyn_0_I4_LSRAM_FL_RADDR_11\ : MUX2L
      port map(A => \I4.bcnt_i_0_il2r_net_1\, B => 
        \LSRAM_FL_RADDRl2r\, S => \I4.LSRAM_FL_RADDR_0_sqmuxa_1\, 
        Y => \I4.LSRAM_FL_RADDR_11\);
    
    \I2.CRC32_796\ : MUX2L
      port map(A => \I2.CRC32l1r_net_1\, B => \I2.N_3918\, S => 
        \I2.N_2826_1_adt_net_794__net_1\, Y => 
        \I2.CRC32_796_net_1\);
    
    \I1.SBYTE_8_0_a2_i_m2l0r\ : MUX2L
      port map(A => F_SO_c, B => REGl83r, S => 
        \I1.sstatel2r_net_1\, Y => \I1.N_405\);
    
    \I3.PIPEB_93\ : AO21
      port map(A => DPR_cl14r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_93_adt_net_160125_\, Y => 
        \I3.PIPEB_93_net_1\);
    
    \I1.REG_74_0_IVL392R_1798\ : NOR2FT
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, Y => 
        \I1.REG_74l392r_adt_net_110870_\);
    
    \I3.PIPEA1l4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_302_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l4r_net_1\);
    
    \I2.PLL_LOCK\ : AND2
      port map(A => \I2.PLL_LOCK_sram\, B => \I2.PLL_LOCK_tdc\, Y
         => PLL_LOCK);
    
    \I2.FID_7_0_IVL23R_989\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl23r_net_1\, 
        Y => \I2.FID_7l23r_adt_net_19209_\);
    
    \I2.MIC_ERR_REGS_338\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl10r_net_1\, B => 
        \I2.MIC_ERR_REGSl9r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_338_net_1\);
    
    FBOUTl3r : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_61_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \FBOUTl3r\);
    
    \I2.REG_1_c2_i\ : NAND2
      port map(A => \I2.N_122\, B => \I2.N_3832_adt_net_101495_\, 
        Y => \I2.N_3831\);
    
    \I3.REG_1l93r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_274_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl93r\);
    
    \I2.STATEe_illegalpipe1\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_3457_ip\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATEe_illegalpipe1_net_1\);
    
    \I3.VDBOFFB_30_IV_0L2R_2455\ : OR3
      port map(A => \I3.VDBoffb_30l2r_adt_net_162747_\, B => 
        \I3.VDBoffb_30l2r_adt_net_162743_\, C => 
        \I3.VDBoffb_30l2r_adt_net_162744_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162750_\);
    
    \I2.FIDl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_441\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl25r);
    
    REGl196r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_97_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl196r\);
    
    \I2.PIPE1_DT_42_1_IVL29R_1360\ : OAI21FTF
      port map(A => \I2.FIRST_TDC_1_sqmuxa_net_1\, B => 
        \I2.TDCDBSl28r_net_1\, C => 
        \I2.PIPE1_DT_42l29r_adt_net_45837_\, Y => 
        \I2.PIPE1_DT_42l29r_adt_net_45839_\);
    
    \I2.N_152_i_0_adt_net_55693_\ : OA21
      port map(A => \I2.PIPE4_DTL17R_635\, B => 
        \I2.PIPE4_DTL15R_637\, C => \I2.RAMDT4L12R_824\, Y => 
        \I2.N_152_i_0_adt_net_55693__net_1\);
    
    \I2.DTE_21_1_IV_0_A2_4_27_M2_E_1000\ : NOR2
      port map(A => \I2.NWPIPE5_305\, B => 
        \I2.REG_0L3R_ADT_NET_848__49\, Y => 
        \I2.N_4030_adt_net_20660_\);
    
    \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834756_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_0_sqmuxa_i_0_N_3_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834756_Rd1__net_1\);
    
    \I3.VDBI_57_IV_0L5R_2246\ : AND2FT
      port map(A => \I3.N_1905_1_adt_net_855384__net_1\, B => 
        \I3.VDBi_43l5r_net_1\, Y => 
        \I3.VDBi_57l5r_adt_net_143854_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I23_G0N\ : AND2FT
      port map(A => \I2.LSRAM_OUTl2r\, B => \I2.PIPE7_DTL2R_702\, 
        Y => \I2.N236\);
    
    \I2.EVNT_NUMl11r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_952_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl11r_net_1\);
    
    \I3.EVREADi_1455\ : DFFC
      port map(CLK => CLK_c, D => \I3.EVREADi_225_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => EVREAD_562);
    
    \I2.PIPE1_DT_42_1_IVL14R_1440\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855224__net_1\, B => 
        \I2.MIC_ERR_REGSl14r_net_1\, C => 
        \I2.PIPE1_DT_42l14r_adt_net_48962_\, Y => 
        \I2.PIPE1_DT_42l14r_adt_net_48963_\);
    
    \I1.REG_74_3_4L380R_1944\ : NAND2FT
      port map(A => \I1.REG_74_5_404_m1_e_0_net_1\, B => 
        \I1.REG_74_12_220_m9_i_a6_0\, Y => 
        \I1.REG_74_3_4_il380r_adt_net_123086_\);
    
    \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855756_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_1_1_net_1\, Y => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855756__net_1\);
    
    \I2.PIPE3_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl4r_net_1\);
    
    \I3.un1_STATE1_11_i\ : AO21FTT
      port map(A => \I3.STATE1_ipl9r\, B => \I3.STATE1_ipl8r\, C
         => \I3.N_1902_adt_net_160759_\, Y => \I3.N_1902\);
    
    \I2.CHB_DATA8_2_i_o2\ : AND2FT
      port map(A => \I2.N_4401\, B => \I2.PIPE7_DTl29r_net_1\, Y
         => \I2.N_4402\);
    
    \I5.SBYTE_9_0l7r\ : MUX2L
      port map(A => \I5.COMMANDl15r_net_1\, B => 
        \I5.SBYTEl6r_net_1\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.SBYTE_9l7r\);
    
    \I3.VDBOFFB_30_IV_0L2R_2446\ : AO21
      port map(A => \REGl335r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l2r_adt_net_162698_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162739_\);
    
    \I3.STATE1_ipl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl8r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl2r_net_1\);
    
    \I2.STATE5_ns_a2_0_a5l1r\ : AND2
      port map(A => \I2.N_4338_1\, B => \I2.STATE5l3r_net_1\, Y
         => \I2.STATE5_ns_il1r\);
    
    \I2.CRC32_12_i_x2l20r\ : XOR2FT
      port map(A => \I2.CRC32l20r_net_1\, B => \I2.N_3962_i_i\, Y
         => \I2.N_111_i_i_0\);
    
    \I2.N_4283_i_0_a2_m1_e_0_662\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__46\, B => 
        \I2.TEMPF_net_1\, Y => \I2.N_4283_I_0_40\);
    
    \I2.OFFSET_37_25l5r\ : MUX2L
      port map(A => \REGl258r\, B => \REGl194r\, S => 
        \I2.PIPE7_DTL27R_89\, Y => \I2.N_832\);
    
    \I3.VDBI_57_0_IV_0L18R_2177\ : AO21
      port map(A => REGl66r, B => \I3.N_1839\, C => 
        \I3.VDBi_57l18r_adt_net_139489_\, Y => 
        \I3.VDBi_57l18r_adt_net_139494_\);
    
    \I1.BYTECNTlde_i_a2_i_847\ : AO21
      port map(A => \I1.N_628\, B => 
        \I1.sstate_ns_i_0_a4_0_1l0r_adt_net_107171_\, C => 
        \I1.N_223_227\, Y => \I1.N_1383_225\);
    
    \I1.BYTECNT_n3_0_a4_0\ : NAND3FFT
      port map(A => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854912__net_1\, B
         => \I1.N_321\, C => \I1.sstatel7r_net_1\, Y => 
        \I1.N_485\);
    
    \I2.RAMDT4l8r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl8r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l8r_net_1\);
    
    \I2.DTE_2_1_0_x2l14r\ : XOR2
      port map(A => \I2.CRC32l10r_net_1\, B => 
        \I2.CRC32l22r_net_1\, Y => \I2.N_126_i_0\);
    
    \I2.PIPE4_DT_I_IL1R_2956\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DT_I_IL1R_473\);
    
    \I3.VDBI_29L4R_2722\ : AO21FTT
      port map(A => \I3.REGMAPL14R_735\, B => 
        \I3.VDBi_20l4r_adt_net_514155_\, C => 
        \I3.VDBi_29l4r_adt_net_621921_\, Y => 
        \I3.VDBi_29l4r_adt_net_144161_\);
    
    \I3.PIPEA_262\ : MUX2L
      port map(A => \I3.PIPEAl31r_net_1\, B => 
        \I3.PIPEA_8l31r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854652__net_1\, Y
         => \I3.PIPEA_262_net_1\);
    
    \I2.N_1170_adt_net_1217__adt_net_855696_\ : BFR
      port map(A => \I2.N_1170_adt_net_1217__net_1\, Y => 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\);
    
    \I2.DT_SRAM_0_i_m2l24r\ : MUX2L
      port map(A => \I2.PIPE10_DTl24r_net_1\, B => 
        \I2.PIPE5_DTl24r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, Y => 
        \I2.N_4192\);
    
    \I2.OFFSET_564\ : MUX2L
      port map(A => \I2.OFFSETl4r_net_1\, B => \I2.OFFSET_37l4r\, 
        S => \I2.UN1_NWPIPE7_2_297\, Y => \I2.OFFSET_564_net_1\);
    
    \I3.REG_1l411r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_218_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl411r);
    
    \I3.STATE1l10r_1621\ : DFFS
      port map(CLK => CLK_c, D => \I3.STATE1_nsl0r\, SET => 
        \I3.N_1311_0\, Q => \I3.STATE1L10R_728\);
    
    \I1.N_41_9_ADT_NET_3739__2799\ : NAND2
      port map(A => \I1.REG_15_SQMUXA_275\, B => 
        \I1.REG_16_SQMUXA_95\, Y => \I1.N_41_9_ADT_NET_3739__93\);
    
    \I5.BITCNT_n1_i\ : OA21FTT
      port map(A => \I5.N_65\, B => \I5.N_94\, C => 
        \I5.N_52_adt_net_9528_\, Y => \I5.N_52\);
    
    \I2.DTE_21_1_IV_0L8R_1310\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855128__net_1\, B => 
        \I2.EVNT_WORDl4r_net_1\, Y => 
        \I2.DTE_21_1l8r_adt_net_38737_\);
    
    \I3.un181_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_558\, B => \I3.N_582\, Y => 
        \I3.un181_reg_ads_0_a2_0_a3_net_1\);
    
    \I1.REG_74_0_IVL240R_1986\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_10_sqmuxa_adt_net_854720__net_1\, Y => 
        \I1.REG_74l240r_adt_net_126727_\);
    
    REGl297r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_198_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl297r\);
    
    INTR1_pad : OB33PH
      port map(PAD => INTR1, A => \GND\);
    
    \I1.REG_1_243\ : MUX2H
      port map(A => \REGl342r\, B => \I1.REG_74l342r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\, Y => 
        \I1.REG_1_243_net_1\);
    
    \I1.REG_30_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_267\, B => 
        \I1.REG_15_sqmuxa_adt_net_1457__net_1\, Y => 
        \I1.REG_30_sqmuxa\);
    
    \I1.REG_1_69\ : MUX2H
      port map(A => \REGl168r\, B => \I1.REG_74l168r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, Y => 
        \I1.REG_1_69_net_1\);
    
    \I2.RAMAD1l9r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_663_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l9r_net_1\);
    
    \I3.PIPEB_106_2317\ : NOR2FT
      port map(A => \I3.PIPEBl27r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_106_adt_net_159579_\);
    
    \I3.VDBoffa_45\ : OR3
      port map(A => \I3.VDBoffa_45_adt_net_164498_\, B => 
        \I3.VDBoffa_31l1r_adt_net_164459_\, C => 
        \I3.VDBoffa_31l1r_adt_net_164460_\, Y => 
        \I3.VDBoffa_45_net_1\);
    
    \I1.REG_1_100\ : MUX2H
      port map(A => \REGl199r\, B => \I1.N_1338\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\, Y => 
        \I1.REG_1_100_net_1\);
    
    REGl215r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_116_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl215r\);
    
    \I3.STATE1_NS_0L0R_2117\ : OA21FTT
      port map(A => \I3.N_268\, B => \I3.DSS_9\, C => 
        \I3.STATE1l10r_net_1\, Y => 
        \I3.STATE1_nsl0r_adt_net_135920_\);
    
    REGl218r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_119_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl218r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I32_Y\ : OA21TTF
      port map(A => \I2.SUB8l11r_adt_net_855580__net_1\, B => 
        \I2.SUB8l12r_adt_net_855576__net_1\, C => 
        \I2.SUB8l13r_adt_net_855564__net_1\, Y => \I2.N297\);
    
    \I3.PIPEA_8l10r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854476__net_1\, B => 
        \I3.N_219\, Y => \I3.PIPEA_8l10r_net_1\);
    
    \I2.SUB8l5r_1600\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_508_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8L5R_707\);
    
    \I2.G_EVNT_NUM_N11_0_1057\ : NOR3FTT
      port map(A => \I2.N_285_1\, B => \I2.N_218\, C => 
        \I2.G_EVNT_NUMl11r_net_1\, Y => 
        \I2.G_EVNT_NUM_n11_adt_net_26872_\);
    
    \I1.ISCK_0_sqmuxa_0_0\ : OR2FT
      port map(A => \I1.N_656\, B => 
        \I1.ISCK_0_sqmuxa_adt_net_134155_\, Y => 
        \I1.ISCK_0_sqmuxa\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I136_Y_0_O2_M4_1570\ : 
        OR3FFT
      port map(A => \I2.N_2358_tz_tz_adt_net_854952__net_1\, B
         => \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_2_adt_net_56515_\, 
        C => \I2.N_74_103\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_adt_net_56806_\);
    
    DTO_padl31r : IOB33PH
      port map(PAD => DTO(31), A => \I2.DTO_1l31r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl31r);
    
    \I3.STATE2_ns_i_i_a5_0_a3l1r\ : AND2FT
      port map(A => \I3.N_1622_1\, B => 
        \I3.STATE2_ns_i_i_a5_0_a3l1r_adt_net_135757_\, Y => 
        \I3.STATE2_ns_i_i_a5_0_a3l1r_net_1\);
    
    \I2.MIC_REG1L2R_2947\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_303_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1L2R_464\);
    
    \I2.DTO_1l8r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l8r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l8r_Rd1__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I48_Y\ : AO21
      port map(A => \I2.N279\, B => \I2.N300_0_adt_net_87046_\, C
         => \I2.N296_0_adt_net_86403_\, Y => \I2.N298_0\);
    
    \I3.STATE1_NS_1_IV_0L5R_2123\ : AND3FTT
      port map(A => \I3.SINGCYC_881\, B => \I3.BLTCYC_net_1\, C
         => \I3.N_90_i_0_1\, Y => 
        \I3.STATE1_nsl5r_adt_net_136320_\);
    
    \I3.REG_1l141r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_189_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl141r\);
    
    \I1.REG_74_0_IVL277R_1942\ : NOR2FT
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l277r_adt_net_122979_\);
    
    \I2.OFFSET_37_18l0r\ : MUX2L
      port map(A => \REGl245r\, B => \REGl181r\, S => 
        \I2.PIPE7_DTL27R_86\, Y => \I2.N_771\);
    
    \I2.DTE_21_1_IV_0L12R_1289\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855124__net_1\, B => 
        \I2.EVNT_WORDl8r_net_1\, Y => 
        \I2.DTE_21_1l12r_adt_net_38281_\);
    
    \I2.BNCID_VECTROR_8_TZ_0_1417\ : AND2
      port map(A => \I2.BNCID_VECTra12_1_net_1\, B => 
        \I2.BNCID_VECTro_8\, Y => 
        \I2.BNCID_VECTror_8_tz_0_i_adt_net_48007_\);
    
    \I5.REG_1l443r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_26_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl443r);
    
    \I3.LWORDS\ : DFFC
      port map(CLK => CLK_c, D => \I3.LWORDS_61_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.LWORDS_net_1\);
    
    \I2.PIPE1_DT_42_1_IV_1L1R_997\ : OA21
      port map(A => \I2.N_148\, B => \I2.N_3870\, C => 
        \I2.CHAINA_EN244_i_adt_net_855260__net_1\, Y => 
        \I2.N_12169_i_adt_net_20407_\);
    
    \I2.WOFFSETl8r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl8r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl8r_Rd1__net_1\);
    
    \I2.DTO_16_1l18r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l18r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l18r_Rd1__net_1\);
    
    \I3.STATE2_ns_i_i_a5_0_a3_1l1r\ : NAND2
      port map(A => \I3.N_203\, B => \I3.STATE2l4r_net_1\, Y => 
        \I3.N_1622_1\);
    
    \I3.LED_R_i_a3\ : OR2FT
      port map(A => TRM_BUSY_c, B => EVRDY_c, Y => LED_R_i_a3);
    
    \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855220_\ : BFR
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__806\, Y => 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855220__net_1\);
    
    \I2.INT_ERRBF1_495\ : OAI21TTF
      port map(A => \I2.N_3876_adt_net_855252__net_1\, B => 
        INT_ERRB_c, C => \I2.INT_ERRBF1_495_adt_net_90378_\, Y
         => \I2.INT_ERRBF1_495_net_1\);
    
    L2R_pad : IB33
      port map(PAD => L2R, Y => L2R_c);
    
    FID_padl30r : OB33PH
      port map(PAD => FID(30), A => FID_cl30r);
    
    \I2.SUB9l6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_574_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l6r_net_1\);
    
    \I2.REG_1_c2_i_a2_0\ : OR2FT
      port map(A => \I2.N_3824_adt_net_90291_\, B => \I2.N_121\, 
        Y => \I2.N_122\);
    
    DPR_padl1r : IB33
      port map(PAD => DPR(1), Y => DPR_cl1r);
    
    \I3.VDBOFFA_31_IV_0L3R_2565\ : AND2
      port map(A => \REGl240r\, B => \I3.REGMAPl27r_net_1\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164028_\);
    
    \I2.OFFSET_37_19l7r\ : MUX2L
      port map(A => \REGl284r\, B => \REGl220r\, S => 
        \I2.PIPE7_DTL27R_86\, Y => \I2.N_786\);
    
    \I2.RAMDT4l7r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl7r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l7r_net_1\);
    
    \I3.PULSE_46_0_iv_i_il3r\ : AO21
      port map(A => PULSEl3r, B => 
        \I3.N_311_adt_net_854752__net_1\, C => \I3.N_1935\, Y => 
        \I3.N_49\);
    
    \I3.PIPEB_92_2331\ : NOR2FT
      port map(A => \I3.PIPEBl13r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_92_adt_net_160167_\);
    
    \I3.RAMAD_VMEl0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_24_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl0r);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__3092\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__862\);
    
    \I2.SUB9l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_573_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l5r_net_1\);
    
    \I2.RAMAD_4_0l4r\ : MUX2H
      port map(A => \I2.RAMAD1l4r_net_1\, B => RAMAD_VMEl4r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_531\);
    
    \I2.CRC32_12_i_0_m2l30r\ : MUX2L
      port map(A => \I2.DT_TEMPl30r_net_1\, B => 
        \I2.DT_SRAMl30r_adt_net_854200__net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854188__net_1\, Y => 
        \I2.N_231_i_i\);
    
    \I3.un136_reg_ads_0_a2_2_a2_0\ : NAND2FT
      port map(A => \I3.VASl2r_net_1\, B => \I3.N_548_366\, Y => 
        \I3.N_549\);
    
    \I2.BNCID_VECTrff_0_265_0\ : AO21
      port map(A => \I2.BNCID_VECTwa12_1_net_1\, B => 
        \I2.BNCID_VECTrff_3_262_0_a2_0\, C => \I2.BNCID_VECTro_0\, 
        Y => \I2.BNCID_VECTrff_0_265_0_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL16R_1414\ : OAI21FTF
      port map(A => REGl436r, B => 
        \I2.N_3234_adt_net_855652__net_1\, C => 
        \I2.PIPE1_DT_42l16r_adt_net_47850_\, Y => 
        \I2.PIPE1_DT_42l16r_adt_net_47851_\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I112_Y_1667\ : AOI21FTT
      port map(A => \I2.N344\, B => 
        \I2.I112_un1_Y_adt_net_71518_\, C => \I2.N328\, Y => 
        \I2.N448_i_adt_net_71546_\);
    
    \I2.PIPE1_DT_42_1_IVL23R_1378\ : OAI21FTF
      port map(A => REGl443r, B => 
        \I2.N_3234_adt_net_855648__net_1\, C => 
        \I2.PIPE1_DT_42l23r_adt_net_46647_\, Y => 
        \I2.PIPE1_DT_42l23r_adt_net_46653_\);
    
    \I3.PIPEB_105_2318\ : NOR2FT
      port map(A => \I3.PIPEBl26r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_105_adt_net_159621_\);
    
    \I3.TCNTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_380_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTl4r_net_1\);
    
    \I2.PIPE5_DT_6l4r\ : MUX2L
      port map(A => \I2.PIPE4_DTl4r_net_1\, B => \I2.N_1073\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, Y
         => \I2.PIPE5_DT_6l4r_net_1\);
    
    \I2.DTE_1_858\ : MUX2L
      port map(A => \I2.DTE_1l20r_Rd1__net_1\, B => 
        \I2.DTE_21_1l20r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\, Y => 
        \I2.DTE_1l20r\);
    
    \I2.LEAD_FLAG6_638_1605\ : NOR2FT
      port map(A => LEAD_FLAGl1r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_638_adt_net_64516_\);
    
    \I2.DTO_cl_63l31r\ : DFFS
      port map(CLK => CLK_c, D => \I2.DTO_cl_63_871_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.DTO_cl_32l31r\);
    
    \I2.FIDl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_428\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl12r);
    
    \I2.DTE_cl_0_sqmuxa_2_0_a2_0_a2_0_910\ : OR2FT
      port map(A => \I2.N_4241_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, Y => 
        \I2.DTE_CL_0_SQMUXA_2_0_288\);
    
    TDCDA_padl28r : IB33
      port map(PAD => TDCDA(28), Y => TDCDA_cl28r);
    
    \I2.DT_TEMP_773\ : MUX2H
      port map(A => \I2.DT_TEMPl12r_net_1\, B => 
        \I2.DT_TEMP_7l12r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_773_net_1\);
    
    \I2.DTE_2_1l9r\ : XOR2
      port map(A => \I2.CRC32l29r_net_1\, B => 
        \I2.DTE_2_1_0l9r_net_1\, Y => \I2.DTE_2_1l9r_net_1\);
    
    \I3.PIPEA_8_0l26r\ : MUX2L
      port map(A => DPR_cl26r, B => \I3.PIPEA1l26r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855356__net_1\, Y => \I3.N_235\);
    
    \I2.DTO_1l24r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l24r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l24r_Rd1__net_1\);
    
    \I2.un2_evnt_word_I_9\ : XOR2
      port map(A => \I2.N_50\, B => 
        \I2.WOFFSETl2r_adt_net_854984__net_1\, Y => \I2.I_9_0\);
    
    \I2.CRC32_12_0_0_m2l21r\ : MUX2L
      port map(A => \I2.DT_TEMPl21r_net_1\, B => 
        \I2.DT_SRAMl21r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854192__net_1\, Y => 
        \I2.N_4039_i_i\);
    
    \I3.VDBi_40_0_i_m2l7r\ : MUX2L
      port map(A => REGl425r, B => REGl441r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_2270\);
    
    \I2.L2TYPE_4_IL5R_1632\ : NAND2FT
      port map(A => \I2.N_4457\, B => \I2.N_4460\, Y => 
        \I2.N_4447_adt_net_68073_\);
    
    \I2.N411_adt_net_4092_\ : AO21
      port map(A => \I2.N411_adt_net_194931__net_1\, B => 
        \I2.N411_adt_net_194981__net_1\, C => \I2.N233\, Y => 
        \I2.N411_adt_net_4092__net_1\);
    
    \I3.REG_1l48r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_149_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl48r);
    
    \I2.ROFFSETl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_913_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl5r_net_1\);
    
    \I2.LSRAM_IN_413\ : MUX2L
      port map(A => \I2.PIPE5_DTl29r_net_1\, B => 
        \I2.LSRAM_INl29r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_413_net_1\);
    
    \I3.REGMAP_i_0_il42r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un191_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il42r_net_1\);
    
    \I1.REG_74_0_iv_i_a2l198r\ : AO21
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_1337_adt_net_130705_\, Y => \I1.N_1337\);
    
    \I2.N_163_adt_net_1241_\ : OA21
      port map(A => \I2.PIPE4_DTL13R_642\, B => 
        \I2.PIPE4_DTL14R_640\, C => \I2.RAMDT4L5R_816\, Y => 
        \I2.N_163_adt_net_1241__net_1\);
    
    \I2.MIC_REG1_0_sqmuxa_0\ : AND2
      port map(A => COM_SERS_561, B => \I2.STATE5l2r_net_1\, Y
         => \I2.MIC_REG1_0_sqmuxa_0_net_1\);
    
    \I1.N_137_adt_net_854760_\ : BFR
      port map(A => \I1.N_137\, Y => 
        \I1.N_137_adt_net_854760__net_1\);
    
    \I2.PIPE8_DT_21l10r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl10r\, B => \I2.N_576\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l10r_net_1\);
    
    DTE_padl5r : IOB33PH
      port map(PAD => DTE(5), A => \I2.DTE_1l5r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl5r);
    
    \I2.DTO_16_1_ivl28r\ : AND2FT
      port map(A => \I2.DTO_16_1_iv_0l28r_net_1\, B => 
        \I2.DTO_16_1_ivl28r_adt_net_28982_\, Y => 
        \I2.DTO_16_1_ivl28r_net_1\);
    
    \I2.OFFSET_37_29l5r\ : MUX2L
      port map(A => \I2.N_856\, B => \I2.N_744\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l5r\);
    
    \I2.DT_TEMPl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_790_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl29r_net_1\);
    
    \I5.sstate2l2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate2_ns_el2r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate2l2r_net_1\);
    
    \I2.N258_0_adt_net_854936_\ : BFR
      port map(A => \I2.N258_0\, Y => 
        \I2.N258_0_adt_net_854936__net_1\);
    
    \I1.REG_74_0_ivl192r\ : AO21
      port map(A => \REGl192r\, B => \I1.N_65\, C => 
        \I1.REG_74l192r_adt_net_131269_\, Y => \I1.REG_74l192r\);
    
    \I1.REG_74L220R_2007\ : AND2FT
      port map(A => \I1.N_1169_adt_net_854820__net_1\, B => 
        \I1.N_89_adt_net_128728_\, Y => \I1.N_89_adt_net_128717_\);
    
    \I3.REGMAP_I_0_IL24R_3023\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un101_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL24R_777\);
    
    \I1.PAGECNT_0l9r_adt_net_835132_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854852__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0l9r_adt_net_835132_Rd1__net_1\);
    
    \I2.ROFFSET_916\ : MUX2H
      port map(A => \I2.ROFFSETl2r_net_1\, B => 
        \I2.ROFFSET_n2_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_916_net_1\);
    
    \I2.PIPE4_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl18r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl18r_net_1\);
    
    \I2.STATE1l12r_adt_net_855176_\ : BFR
      port map(A => \I2.STATE1L12R_646\, Y => 
        \I2.STATE1l12r_adt_net_855176__net_1\);
    
    \I3.UN1_EVREAD_DS_1_SQMUXA_1_2311\ : AND3FTT
      port map(A => \I3.N_281\, B => \I3.un15_anycyc_net_1\, C
         => \I3.N_1860_2\, Y => 
        \I3.un1_EVREAD_DS_1_sqmuxa_1_adt_net_158292_\);
    
    \I2.PIPE5_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_680_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl4r_net_1\);
    
    CHAINB_EN244_pad : OB33PH
      port map(PAD => CHAINB_EN244, A => 
        \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\);
    
    \I2.PIPE4_DTl14r_1532\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL14R_639\);
    
    \I1.PAGECNTL7R_2978\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_320_adt_net_854876__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL7R_525\);
    
    \I2.SUB9_1_ADD_18x18_fast_I152_Y_0\ : XOR2FT
      port map(A => \I2.N_3558_i_adt_net_855584__net_1\, B => 
        \I2.SUB8l15r_adt_net_855572__net_1\, Y => 
        \I2.ADD_18x18_fast_I152_Y_0\);
    
    \I5.REG_1_20\ : MUX2H
      port map(A => \I5.TEMPDATAl1r_net_1\, B => REGl437r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\, Y
         => \I5.REG_1_20_net_1\);
    
    \I2.RAMDT4L12R_3070\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_824\);
    
    \I2.I_1337_G_1\ : XOR2FT
      port map(A => \I2.SUB8L5R_707\, B => \I2.OFFSETL2R_678\, Y
         => \I2.G_1_4\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I154_Y_0_2693\ : NAND2FT
      port map(A => \I2.N502_i_0_adt_net_490392_\, B => 
        \I2.N498_0_adt_net_598321_\, Y => \I2.N502_i_0\);
    
    \I1.BYTECNT_314\ : MUX2H
      port map(A => \I1.BYTECNTl0r_net_1\, B => \I1.BYTECNT_n0\, 
        S => \I1.N_1383\, Y => \I1.BYTECNT_314_net_1\);
    
    \I1.REG_74_0_IVL304R_1914\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l304r_adt_net_120524_\);
    
    \I3.VDBI_57_0_IVL31R_2140\ : AO21
      port map(A => \I3.VDBil31r_net_1\, B => 
        \I3.N_1910_0_adt_net_854340__net_1\, C => 
        \I3.VDBi_57l31r_adt_net_137838_\, Y => 
        \I3.VDBi_57l31r_adt_net_137844_\);
    
    \I2.DT_TEMP_775\ : MUX2H
      port map(A => \I2.DT_TEMPl14r_net_1\, B => 
        \I2.DT_TEMP_7l14r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_775_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I121_Y_i_a3_0\ : AO21TTF
      port map(A => \I2.RAMDT4L12R_146\, B => 
        \I2.PIPE4_DTl5r_adt_net_854412__net_1\, C => \I2.N_67\, Y
         => \I2.ADD_21x21_fast_I121_Y_i_a3_0_i_0\);
    
    \I1.REG_74_0_IVL396R_1794\ : NOR2FT
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, Y => 
        \I1.REG_74l396r_adt_net_110526_\);
    
    \I4.bcntl0r\ : DFFC
      port map(CLK => CLK_c, D => \I4.bcnt_5_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I4.bcntl0r_net_1\);
    
    \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344_\ : BFR
      port map(A => \I3.STATE1_ipl3r_adt_net_854364__net_1\, Y
         => 
        \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344__net_1\);
    
    \I2.DTOSl14r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl14r, Q => 
        \I2.DTOSl14r_net_1\);
    
    \I2.DTO_16_1_IV_0_0L29R_1073\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.N_4159\, C => \I2.DTO_16_1l29r_adt_net_28732_\, Y => 
        \I2.DTO_16_1l29r_adt_net_28739_\);
    
    \I1.REG_1_215\ : MUX2H
      port map(A => \REGl314r\, B => \I1.REG_74l314r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_215_net_1\);
    
    \I1.REG_1_108\ : MUX2H
      port map(A => \REGl207r\, B => \I1.N_1346\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_108_net_1\);
    
    \I2.un3_tdcgda1_1_adt_net_821__adt_net_855104_\ : BFR
      port map(A => \I2.un3_tdcgda1_1_adt_net_821__net_1\, Y => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855104__net_1\);
    
    \I2.DTE_21_1_iv_0l20r\ : AO21
      port map(A => \I2.DTE_1l20r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.DTE_21_1l20r_adt_net_37615_\, Y => \I2.DTE_21_1l20r\);
    
    \I2.PIPE8_DT_16_0l3r\ : MUX2H
      port map(A => \I2.PIPE8_DTl3r_net_1\, B => 
        \I2.PIPE7_DTl3r_net_1\, S => 
        \I2.N_565_0_adt_net_855728__net_1\, Y => \I2.N_569\);
    
    \I3.VDBi_40_0_i_m2l13r\ : MUX2L
      port map(A => REGl431r, B => REGl447r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_2276\);
    
    \I2.OFFSET_37_1l6r\ : MUX2L
      port map(A => \REGl355r\, B => \REGl291r\, S => 
        \I2.PIPE7_DTL27R_65\, Y => \I2.N_641\);
    
    \I1.un1_sbyte13_1_i_0_s\ : AO21
      port map(A => \I1.N_370\, B => 
        \I1.un1_sbyte13_1_i_1_adt_net_106369_\, C => 
        \PULSE_0L0R_ADT_NET_834380_RD1__199\, Y => 
        \I1.un1_sbyte13_1_i_1\);
    
    \I3.REG_1_ml71r\ : AND2
      port map(A => REGl71r, B => 
        \I3.REGMAPl9r_adt_net_854312__net_1\, Y => 
        \I3.VDBi_20l23r\);
    
    \I1.REG_74_0_IV_0_0L254R_1971\ : AND2
      port map(A => \FBOUTl1r\, B => \I1.N_596\, Y => 
        \I1.REG_74l254r_adt_net_125314_\);
    
    \I2.PIPE4_DTl0r_1149\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL0R_411\);
    
    \I2.CRC32l17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_812_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l17r_net_1\);
    
    \I1.SBYTE_8_0_i_a2_0l3r\ : OR2FT
      port map(A => \I1.sstatel2r_net_1\, B => 
        \I1.sstatel9r_net_1\, Y => \I1.N_603_i\);
    
    \I3.REG_1l78r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_179_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl78r);
    
    \I2.BNCID_VECTrff_6_259_0\ : AO21
      port map(A => \I2.BNCID_VECTwa14_1_net_1\, B => 
        \I2.BNCID_VECTrff_7_258_0_a2_0\, C => \I2.BNCID_VECTro_6\, 
        Y => \I2.BNCID_VECTrff_6_259_0_net_1\);
    
    \I2.SUB9l10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_578_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l10r_net_1\);
    
    \I2.FCNTe_i\ : AOI21FTT
      port map(A => \I2.N_3267_adt_net_25763_\, B => \I2.N_3277\, 
        C => \I2.STATE1l13r_net_1\, Y => \I2.N_3267\);
    
    \I2.UN5_TDCGDA1_1012\ : NOR2
      port map(A => \I2.un7_tdcgda1_1_i_i\, B => 
        \I2.un7_tdcgda1_0_i_i\, Y => 
        \I2.un5_tdcgda1_adt_net_21626_\);
    
    \I3.un2_vsel_1_i_0_a2\ : NAND3FFT
      port map(A => \I3.N_1918\, B => \I3.N_2055_adt_net_134992_\, 
        C => \I3.SELBASE32_net_1\, Y => \I3.N_2055\);
    
    \I2.un1_NWPIPE7_2_919\ : OR2FT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855160__net_1\, B
         => \I2.UN1_NWPIPE7_2_ADT_NET_73606__324\, Y => 
        \I2.UN1_NWPIPE7_2_297\);
    
    \I3.VSEL_0_a3_0_a3_0\ : NOR2
      port map(A => \I3.ASBS_net_1\, B => \I3.N_1918\, Y => 
        \I3.VSEL_0\);
    
    \I2.DTE_2_1_0l6r\ : XOR2
      port map(A => \I2.CRC32l14r_net_1\, B => 
        \I2.CRC32l2r_net_1\, Y => \I2.DTE_2_1_0l6r_net_1\);
    
    \I2.CRC32_12_il22r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_130_i_0_i_0\, Y => 
        \I2.N_3939\);
    
    \I2.MTDCRESB\ : DFFC
      port map(CLK => CLK_c, D => \I2.MTDCRESB_379_net_1\, CLR
         => \I2.un15_clear_stat_i\, Q => MTDCRESB_c);
    
    \I1.REG_1_98\ : MUX2H
      port map(A => \REGl197r\, B => \I1.N_129\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\, Y => 
        \I1.REG_1_98_net_1\);
    
    \I3.PULSE_46_0_IV_0_0L8R_2289\ : AND3
      port map(A => VDB_inl0r, B => \I3.REGMAPl56r_net_1\, C => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        Y => \I3.PULSE_46l8r_adt_net_146836_\);
    
    \I2.un7_bnc_id_1_I_8\ : AND2
      port map(A => \I2.BNC_IDL1R_394\, B => \I2.BNC_IDL0R_395\, 
        Y => \I2.N_45\);
    
    \I1.un1_sbyte13_1_i_0_s_829\ : AO21
      port map(A => \I1.N_370_adt_net_854904__net_1\, B => 
        \I1.un1_sbyte13_1_i_1_adt_net_106369__adt_net_854528__net_1\, 
        C => \PULSE_0L0R_ADT_NET_834380_RD1__199\, Y => 
        \I1.UN1_SBYTE13_1_I_1_207\);
    
    \I2.FCNT_n2_tz\ : XOR2FT
      port map(A => \I2.FCNT_c1\, B => \I2.FCNTl2r_net_1\, Y => 
        \I2.FCNT_n2_tz_i\);
    
    \I2.END_EVNT5_1144_1732\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT5_839\);
    
    \I3.REG3l6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_131_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l6r_net_1\);
    
    \I2.N_40_adt_net_589963_\ : NOR3FFT
      port map(A => \I2.N_45_0\, B => 
        \I2.N_40_adt_net_589803__net_1\, C => 
        \I2.N525_adt_net_57834_\, Y => 
        \I2.N_40_adt_net_589963__net_1\);
    
    \I2.DTE_21_1_IV_0L12R_1288\ : AND2
      port map(A => \I2.STATE2L3R_440\, B => \I2.N_3966\, Y => 
        \I2.DTE_21_1l12r_adt_net_38279_\);
    
    \I2.L2RF2\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2RF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L2RF2_net_1\);
    
    \I2.FID_7_0_ivl9r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl9r_net_1\, 
        C => \I2.FID_7l9r_adt_net_92653_\, Y => \I2.FID_7l9r\);
    
    \I1.BYTECNTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_308_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTl6r_net_1\);
    
    \I3.VDBI_57_0_IV_0L27R_2149\ : AO21
      port map(A => REGl75r, B => \I3.N_1839\, C => 
        \I3.VDBi_57l27r_adt_net_138433_\, Y => 
        \I3.VDBi_57l27r_adt_net_138440_\);
    
    \I2.PIPE4_DTl12r_1248\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL12R_510\);
    
    \I2.PIPE8_DT_21l20r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl20r\, B => 
        \I2.PIPE8_DT_16l20r_net_1\, S => \I2.NWPIPE7_net_1\, Y
         => \I2.PIPE8_DT_21l20r_net_1\);
    
    \I2.N_40_adt_net_1100_\ : NAND3FFT
      port map(A => \I2.N_70_adt_net_54406__net_1\, B => 
        \I2.N_40_adt_net_589963__net_1\, C => 
        \I2.N_114_adt_net_275711_\, Y => 
        \I2.N_40_adt_net_1100__net_1\);
    
    ADO_padl10r : OB33PH
      port map(PAD => ADO(10), A => ADO_cl10r);
    
    \I4.STATE1l1r\ : DFFC
      port map(CLK => CLK_c, D => \I4.STATE1_nsl1r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I4.STATE1l1r_net_1\);
    
    \I2.PIPE1_DTl2r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_729_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl2r_net_1\);
    
    \I2.DTO_9_IVL1R_1208\ : NOR2
      port map(A => \I2.N_4283_I_0_235\, B => 
        \I2.DT_TEMPl1r_net_1\, Y => 
        \I2.DTO_9_ivl1r_adt_net_35072_\);
    
    \I3.STATE1_ILLEGAL_2130\ : AO21
      port map(A => \I3.STATE1_ipl4r\, B => \I3.N_1174\, C => 
        \I3.N_1193_ip_adt_net_136552_\, Y => 
        \I3.N_1193_ip_adt_net_136553_\);
    
    REGl170r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_71_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl170r\);
    
    \I1.REG_74_0_ivl195r\ : AO21
      port map(A => \REGl195r\, B => \I1.N_65_92\, C => 
        \I1.REG_74l195r_adt_net_131011_\, Y => \I1.REG_74l195r\);
    
    \I2.DTO_16_1_IV_0_O7L29R_1070\ : AND2FT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl29r_net_1\, Y => \I2.N_4159_adt_net_28676_\);
    
    \I3.TICKil0r_1448\ : DFFC
      port map(CLK => CLK_c, D => \I3.un6_tcnt1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TICKL0R_555);
    
    \I1.BYTECNTL2R_2844\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_312_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTL2R_213\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2517\ : AO21
      port map(A => \REGl203r\, B => \I3.REGMAPl22r_net_1\, C => 
        \I3.N_2070_adt_net_163454_\, Y => 
        \I3.N_2070_adt_net_163498_\);
    
    \I3.VDBI_57_0_IV_0_0L8R_2224\ : AND2FT
      port map(A => \I3.REGMAPl55r_net_1\, B => 
        \I3.VDBi_57l8r_adt_net_142678_\, Y => 
        \I3.VDBi_57l8r_adt_net_142786_\);
    
    \I2.MIC_ERR_REGS_333\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl5r_net_1\, B => 
        \I2.MIC_ERR_REGSl4r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_333_net_1\);
    
    \I1.sstate_ns_0_iv_0_0l1r\ : OAI21TTF
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.N_346\, C => \I1.sstate_nsl1r_adt_net_107663_\, Y => 
        \I1.sstate_nsl1r\);
    
    \I2.SUB9_569\ : MUX2H
      port map(A => \I2.SUB9l1r_net_1\, B => \I2.SUB8l2r_net_1\, 
        S => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_569_net_1\);
    
    \I3.REG_1_266\ : MUX2H
      port map(A => REGl85r, B => \I3.N_1631\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_266_0\);
    
    \I2.PIPE1_DT_42_1_iv_2l25r\ : OA21FTF
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, B => 
        \I2.TDCDBSl25r_net_1\, C => \I2.PIPE1_DT_42_1_iv_1_il25r\, 
        Y => \I2.PIPE1_DT_42_1_iv_2l25r_net_1\);
    
    \I2.SUB9_571\ : MUX2H
      port map(A => \I2.SUB9l3r_net_1\, B => \I2.SUB9_1l3r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_571_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl30r\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, B => 
        \I2.PIPE1_DT_30l30r_net_1\, C => 
        \I2.PIPE1_DT_42l30r_adt_net_45595_\, Y => 
        \I2.PIPE1_DT_42l30r\);
    
    \I2.OFFSET_37_28l0r\ : MUX2L
      port map(A => \I2.N_843\, B => \I2.N_795\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_851\);
    
    \I2.L2ARR_n1\ : XOR2
      port map(A => \I2.L2ARRl1r_net_1\, B => \I2.L2ARRl0r_net_1\, 
        Y => \I2.L2ARR_n1_net_1\);
    
    \I2.DT_TEMPl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_789_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl28r_net_1\);
    
    \I3.REG_1l103r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_284_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl103r);
    
    \I2.SUB8_523_2739\ : AND3
      port map(A => \I2.N288_0\, B => 
        \I2.N475_adt_net_4127__net_1\, C => 
        \I2.SUB8_523_adt_net_566364_\, Y => 
        \I2.SUB8_523_adt_net_670055_\);
    
    \I2.G_EVNT_NUM_927\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl7r_net_1\, B => \I2.N_4639\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_927_net_1\);
    
    \I2.un1_STATE1_40_0_o2_2\ : NOR3FTT
      port map(A => \I2.CHAINA_EN244_i_adt_net_855264__net_1\, B
         => \I2.END_CHAINA1_net_1\, C => \I2.N_3272_345\, Y => 
        \I2.N_3898_i\);
    
    \I3.PIPEA_8l5r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854480__net_1\, B => 
        \I3.N_214\, Y => \I3.PIPEA_8l5r_net_1\);
    
    \I3.REG_1l92r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_273_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl92r\);
    
    \I2.PIPE1_DT_42_1_IVL8R_1476\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855228__net_1\, B => 
        \I2.MIC_ERR_REGSl8r_net_1\, C => 
        \I2.PIPE1_DT_42l8r_adt_net_50444_\, Y => 
        \I2.PIPE1_DT_42l8r_adt_net_50445_\);
    
    \I2.DTE_1l11r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l11r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l11r_Rd1__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I163_Y_1692\ : OA21FTF
      port map(A => \I2.N350\, B => \I2.N357_1\, C => \I2.N349\, 
        Y => \I2.N492_i_adt_net_89450_\);
    
    \I2.DTE_21_1_iv_0_a2_4_27_m2_e\ : OAI21FTF
      port map(A => \I2.REG_0L3R_ADT_NET_848__49\, B => 
        \I2.NWPIPE10_net_1\, C => \I2.N_4030_adt_net_20660_\, Y
         => \I2.N_4030\);
    
    \I2.PIPE7_DTl25r_1577\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL25R_684\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_782\ : AO21
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__26\, B => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_a5_2_i_adt_net_2404__net_1\, C
         => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__162\, 
        Y => \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_160\);
    
    \I2.OFFSET_37_29l7r\ : MUX2L
      port map(A => \I2.N_858\, B => \I2.N_746\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l7r\);
    
    
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536_\ : 
        BFR
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__net_1\, 
        Y => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536__net_1\);
    
    \I3.PIPEB_89\ : AO21
      port map(A => DPR_cl10r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_89_adt_net_160293_\, Y => 
        \I3.PIPEB_89_net_1\);
    
    \I3.un224_reg_ads_0_a2_3_a2_996\ : NAND2
      port map(A => \I3.LWORDS_788\, B => \I3.N_545\, Y => 
        \I3.N_546_374\);
    
    \I3.REGMAPL57R_3054\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un231_reg_ads_0_a2_4_a3_net_1\, Q => 
        \I3.REGMAPL57R_808\);
    
    \I2.G_EVNT_NUM_m_1_i_0_o2l8r_676\ : OR2FT
      port map(A => \I2.N_176_i\, B => \I2.N_4641_56\, Y => 
        \I2.N_223_54\);
    
    \I5.COMMAND_4l12r\ : MUX2L
      port map(A => \I5.AIR_WDATAl8r_net_1\, B => REGl113r, S => 
        REGl7r, Y => \I5.COMMAND_4l12r_net_1\);
    
    \I2.RAMDT4L0R_3016\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl0r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L0R_770\);
    
    \I2.PIPE1_DT_42_1_IVL16R_1410\ : AND2
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl48r_net_1\, Y => 
        \I2.PIPE1_DT_42l16r_adt_net_47833_\);
    
    \I2.N475_adt_net_4127_\ : AO21
      port map(A => \I2.I180_un1_Y_adt_net_240115_\, B => 
        \I2.N475_adt_net_378647__net_1\, C => 
        \I2.N475_adt_net_460353__net_1\, Y => 
        \I2.N475_adt_net_4127__net_1\);
    
    \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__2828\ : OAI21TTF
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100__net_1\, B
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        C => \I2.FIRST_TDC_1_sqmuxa_net_1\, Y => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__172\);
    
    \I2.REG_1_n4\ : XOR2FT
      port map(A => \I2.N_3832\, B => \I2.REG_1_n4_0_net_1\, Y
         => \I2.REG_1_n4_net_1\);
    
    \I1.REG_1_150\ : MUX2H
      port map(A => \REGl249r\, B => \I1.REG_74l249r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_150_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I178_Y_2728\ : AND2
      port map(A => \I2.N297_0\, B => \I2.N301_2\, Y => 
        \I2.N479_adt_net_642172_\);
    
    \PULSEl0r_adt_net_854532_\ : BFR
      port map(A => \PULSEl0r_adt_net_854536__net_1\, Y => 
        \PULSEl0r_adt_net_854532__net_1\);
    
    \I2.N475_adt_net_378647_\ : AND3
      port map(A => \I2.N285\, B => \I2.N479_adt_net_642172_\, C
         => \I2.I180_un1_Y_adt_net_215260_\, Y => 
        \I2.N475_adt_net_378647__net_1\);
    
    \I2.FCNTl0r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_947_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.FCNT_c0\);
    
    \I1.REG_74_0_ivl213r\ : AO21
      port map(A => \REGl213r\, B => \I1.N_89_165\, C => 
        \I1.REG_74l213r_adt_net_129378_\, Y => \I1.REG_74l213r\);
    
    \I2.DTE_1l22r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l22r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l22r_Rd1__net_1\);
    
    \I1.PAGECNT_n7_i_i_o2\ : NOR2
      port map(A => \I1.N_310_Rd1__net_1\, B => 
        \I1.N_299_adt_net_833868_Rd1__net_1\, Y => \I1.N_345\);
    
    \I2.G_EVNT_NUM_n3_i_0_o2\ : AND2FT
      port map(A => \I2.N_187\, B => \I2.G_EVNT_NUML3R_399\, Y
         => \I2.N_189\);
    
    DTO_padl3r : IOB33PH
      port map(PAD => DTO(3), A => \I2.DTO_1l3r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl3r);
    
    \I1.REG_74_0_IVL193R_2041\ : AND2
      port map(A => \FBOUTl4r\, B => \I1.REG_4_sqmuxa\, Y => 
        \I1.REG_74l193r_adt_net_131183_\);
    
    \I1.REG_74_0_IVL290R_1929\ : NOR2FT
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l290r_adt_net_121861_\);
    
    \I1.REG_74_0_iv_i_a2l207r\ : AO21
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, C => 
        \I1.N_1346_adt_net_129931_\, Y => \I1.N_1346\);
    
    \I2.DTO_16_1_IVL23R_1100\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.G_EVNT_NUMl7r_net_1\, Y
         => \I2.DTO_16_1l23r_adt_net_30106_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I184_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTL14R_640\, Y => \I2.ADD_21x21_fast_I184_Y_0\);
    
    \I2.REG_0l3r_adt_net_848__adt_net_854224_\ : BFR
      port map(A => 
        \I2.REG_0l3r_adt_net_848__adt_net_854228__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__adt_net_854224__net_1\);
    
    \I2.PIPE5_DTl22r_1558\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_698_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL22R_665\);
    
    \I2.DT_SRAM_0l20r\ : MUX2L
      port map(A => \I2.PIPE10_DTl20r_net_1\, B => 
        \I2.PIPE5_DTl20r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, Y => 
        \I2.N_888\);
    
    \I3.un68_reg_ads_0_a2_3_a3\ : AND2
      port map(A => \I3.N_545\, B => 
        \I3.un68_reg_ads_0_a2_3_a3_adt_net_166224_\, Y => 
        \I3.un68_reg_ads_0_a2_3_a3_net_1\);
    
    PULSEl0r : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854736__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \PULSEl0r\);
    
    \I3.VADm_0_a3l12r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl12r_net_1\, Y => \I3.VADml12r\);
    
    \I2.FIDl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_430\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl14r);
    
    \I1.BYTECNT_n5_i_0\ : AND2FT
      port map(A => \I1.N_223_227\, B => 
        \I1.N_75_adt_net_109200_\, Y => \I1.N_75\);
    
    \I2.DT_TEMPl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_765_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl4r_net_1\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_m9_i_a5\ : AND3FTT
      port map(A => \I2.REG_0L3R_ADT_NET_848__49\, B => 
        \I2.END_EVNT5_839\, C => 
        \I2.N_4646_1_ADT_NET_1645_RD1__890\, Y => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_N_20_i\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__2849\ : NOR3FFT
      port map(A => \I2.END_EVNT5_840\, B => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\, C => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_M3_238\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__236\);
    
    \I2.TOKOUT_FL_674_adt_net_1115_\ : AO21
      port map(A => \I2.TOKOUTAS_net_1\, B => 
        \I2.STATE1l10r_net_1\, C => 
        \I2.TOKOUT_FL_674_adt_net_61290__net_1\, Y => 
        \I2.TOKOUT_FL_674_adt_net_1115__net_1\);
    
    \I2.DTO_16_1l20r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l20r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l20r_Rd1__net_1\);
    
    \I2.CRC32_805\ : MUX2L
      port map(A => \I2.CRC32l10r_net_1\, B => \I2.N_3927\, S => 
        \I2.N_2826_1_ADT_NET_794__332\, Y => \I2.CRC32_805_net_1\);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854660_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854660__net_1\);
    
    \I2.LSRAM_RADDRl0r\ : MUX2L
      port map(A => \LSRAM_FL_RADDRl0r\, B => 
        \I2.LSRAM_RADDRil0r_net_1\, S => FLUSH, Y => 
        \I2.LSRAM_RADDRl0r_net_1\);
    
    \I2.PIPE9_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_279_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl10r_net_1\);
    
    \I1.REG_19_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_127_i\, B => \I1.N_242\, Y => 
        \I1.REG_19_sqmuxa\);
    
    \I3.UN15_TCNT4_2644\ : NOR2
      port map(A => \I3.TCNT4_i_0_il0r_net_1\, B => 
        \I3.TCNT4l3r_net_1\, Y => \I3.un15_tcnt4_adt_net_165650_\);
    
    \I5.AIR_WDATA_60\ : MUX2L
      port map(A => \I5.AIR_WDATAl10r_net_1\, B => 
        \I5.AIR_WDATA_9l10r_net_1\, S => \I5.N_461\, Y => 
        \I5.AIR_WDATA_60_net_1\);
    
    \I3.N_178_ADT_NET_1360__2807\ : OR2FT
      port map(A => \I3.N_2083\, B => 
        \I3.N_178_adt_net_134608__net_1\, Y => 
        \I3.N_178_ADT_NET_1360__127\);
    
    \I1.RAMDT_SPI_1l4r\ : DFFC
      port map(CLK => CLK_c, D => \FBOUTl4r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.RAMDT_SPI_1l4r_net_1\);
    
    \I3.TCNT1_c1\ : AND2
      port map(A => \I3.TCNT1l0r_net_1\, B => 
        \I3.TCNT1_i_0_il1r_net_1\, Y => \I3.TCNT1_c1_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I198_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl2r\, B => 
        \I2.PIPE7_DTl2r_net_1\, Y => \I2.SUB_21x21_fast_I198_Y_0\);
    
    \I2.DTO_16_1_IV_0L8R_1180\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.N_3967\, C => \I2.DTO_16_1l8r_adt_net_33478_\, Y => 
        \I2.DTO_16_1l8r_adt_net_33488_\);
    
    \I2.PIPE5_DT_689\ : MUX2L
      port map(A => \I2.PIPE5_DTl13r_net_1\, B => 
        \I2.PIPE5_DT_6l13r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_689_net_1\);
    
    \I2.OFFSET_37_15l4r\ : MUX2L
      port map(A => \REGl233r\, B => \REGl169r\, S => 
        \I2.PIPE7_DTL27R_70\, Y => \I2.N_751\);
    
    \I2.REG_1_c4_i_o2\ : NAND3
      port map(A => REGL35R_564, B => REGL36R_565, C => 
        \I2.N_3845\, Y => \I2.N_3847\);
    
    \I1.REG_74_0_iv_0l359r\ : AO21
      port map(A => \REGl359r\, B => \I1.N_661\, C => 
        \I1.REG_74l359r_adt_net_114955_\, Y => \I1.REG_74l359r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I203_Y\ : XOR2FT
      port map(A => \I2.N510\, B => \I2.SUB_21x21_fast_I203_Y_0\, 
        Y => \I2.SUB8_2l7r\);
    
    \I1.PAGECNTL9R_3079\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854856__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL9R_835\);
    
    \I3.PIPEA_8l20r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854464__net_1\, B => 
        \I3.N_229\, Y => \I3.PIPEA_8l20r_net_1\);
    
    \I1.sstatel6r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl4r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel6r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I23_Y\ : AND2
      port map(A => \I2.N268\, B => \I2.N288_adt_net_68878_\, Y
         => \I2.N288\);
    
    \I2.ENDF_1140\ : DFFC
      port map(CLK => CLK_c, D => \I2.ENDF_712_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ENDF_402\);
    
    \I2.L2SERVl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_920_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEl14r\);
    
    \I1.LUT_55\ : AO21FTT
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.N_606_Rd1__net_1\, C => \I1.LUT_55_adt_net_133935_\, 
        Y => \I1.LUT_55_net_1\);
    
    DPR_padl23r : IB33
      port map(PAD => DPR(23), Y => DPR_cl23r);
    
    \I2.G_EVNT_NUM_n7_i_a2\ : NOR2
      port map(A => \I2.N_198\, B => \I2.G_EVNT_NUMl7r_net_1\, Y
         => \I2.N_281\);
    
    \I3.PULSE_46_0_IV_0_0L6R_2290\ : NOR2FT
      port map(A => PULSEl6r, B => \I3.N_291\, Y => 
        \I3.PULSE_46l6r_adt_net_147009_\);
    
    \I1.REG_74_0_IVL348R_1865\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l348r_adt_net_116326_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I91_Y_0\ : OR2FT
      port map(A => \I2.N_17_0\, B => \I2.N_93_0\, Y => 
        \I2.N394_0\);
    
    \I3.TCNT1l4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT1_n4_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT1l4r_net_1\);
    
    TICKl3r : DFFC
      port map(CLK => CLK_c, D => \I3.un15_tcnt4_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \TICKl3r\);
    
    \I1.REG_0_sqmuxa_i_0_a2\ : AND3
      port map(A => \I1.sstatel0r_net_1\, B => \I1.N_324_24\, C
         => \I1.BITCNTl2r_net_1\, Y => \I1.N_598\);
    
    \I2.EVNT_NUMl6r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_957_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl6r_net_1\);
    
    \I1.BYTECNT_N4_I_1779\ : XOR2
      port map(A => \I1.BYTECNT_i_0_il4r_net_1\, B => \I1.N_327\, 
        Y => \I1.N_1381_adt_net_109130_\);
    
    \I3.VDBoffb_55\ : OR3
      port map(A => \I3.VDBoffb_55_adt_net_162600_\, B => 
        \I3.VDBoffb_30l3r_adt_net_162559_\, C => 
        \I3.VDBoffb_30l3r_adt_net_162560_\, Y => 
        \I3.VDBoffb_55_net_1\);
    
    \I1.REG_74_9_0_o2l372r\ : NAND2
      port map(A => \I1.N_273_5_i\, B => 
        \I1.REG_74_4_i_a2_404_N_4_i\, Y => \I1.N_374\);
    
    \I3.PULSEl9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_339_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl9r);
    
    \I1.REG_1_302\ : MUX2H
      port map(A => \REGl401r\, B => \I1.REG_74l401r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\, Y => 
        \I1.REG_1_302_net_1\);
    
    \I3.VDBi_31l22r\ : MUX2L
      port map(A => \I3.REGl155r\, B => \I3.VDBi_20l22r\, S => 
        \I3.REGMAPl17r_adt_net_854280__net_1\, Y => 
        \I3.VDBi_31l22r_net_1\);
    
    \I3.REG_1l413r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_220_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl413r);
    
    \I2.un7_bnc_id_1_I_65\ : AND2
      port map(A => \I2.BNC_IDl10r_net_1\, B => \I2.N_11_1\, Y
         => \I2.N_4_0\);
    
    \I2.BNC_IDl11r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_66_0\, CLR => 
        \I2.N_4618_i_0\, SET => \I2.N_4606_i_0\, Q => 
        \I2.BNC_IDl11r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I151_Y_i_a4_0\ : OR3
      port map(A => \I2.N_41_adt_net_54984_\, B => 
        \I2.N_163_adt_net_1241__net_1\, C => 
        \I2.N_41_adt_net_54991_\, Y => \I2.N_41\);
    
    \I2.PIPE8_DT_16_0l2r\ : MUX2H
      port map(A => \I2.PIPE8_DTl2r_net_1\, B => 
        \I2.PIPE7_DTl2r_net_1\, S => 
        \I2.N_565_0_adt_net_855728__net_1\, Y => \I2.N_568\);
    
    \I2.PIPE4_DTL9R_3081\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL9R_845\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__3104\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__890\);
    
    \I3.VDBi_57_0_ivl14r\ : OR2
      port map(A => \I3.VDBi_57l14r_adt_net_140192_\, B => 
        \I3.VDBi_57l14r_adt_net_140197_\, Y => \I3.VDBi_57l14r\);
    
    \I1.REG_1_122\ : MUX2H
      port map(A => \REGl221r\, B => \I1.REG_74l221r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_122_net_1\);
    
    \I2.SUB8_1_sqmuxa_0_adt_net_855156_\ : BFR
      port map(A => \I2.SUB8_1_sqmuxa_0\, Y => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855156__net_1\);
    
    TDCDA_padl30r : IB33
      port map(PAD => TDCDA(30), Y => TDCDA_cl30r);
    
    \I3.VDBi_16_m_i_o3l3r\ : OR2
      port map(A => \I3.REGMAPL8R_741\, B => \I3.REGMAPl9r_net_1\, 
        Y => \I3.N_1907\);
    
    NOEMIC_pad : OB33PH
      port map(PAD => NOEMIC, A => NOEMIC_c);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I53_Y_1281\ : NAND2
      port map(A => \I2.N273_547\, B => \I2.N270_0_545\, Y => 
        \I2.N303_0_543\);
    
    \I2.FID_7_0_IVL30R_975\ : AND2
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTES_i_0_il30r\, 
        Y => \I2.FID_7l30r_adt_net_18551_\);
    
    \I2.SRAM_EVNT_n4\ : XOR2
      port map(A => \I2.N_3828\, B => \I2.SRAM_EVNT_n4_0_net_1\, 
        Y => \I2.SRAM_EVNT_n4_net_1\);
    
    \I5.REG_1_25\ : MUX2H
      port map(A => \I5.TEMPDATAl6r_net_1\, B => REGl442r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_25_net_1\);
    
    \I1.PAGECNTlde_0_o2\ : OAI21FTF
      port map(A => \I1.SSTATEL10R_882\, B => \I1.N_328_I_0_498\, 
        C => \PULSE_0L0R_ADT_NET_834380_RD1__201\, Y => 
        \I1.N_292\);
    
    \I3.VDBoffb_30_iv_0l4r\ : AND2
      port map(A => \REGl369r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162314_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I182_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl12r_net_1\, Y => 
        \I2.ADD_21x21_fast_I182_Y_0\);
    
    \I2.FID_7_ivl3r\ : OR2
      port map(A => \I2.FID_7l3r_adt_net_93258_\, B => 
        \I2.FID_7l3r_adt_net_93259_\, Y => \I2.FID_7l3r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I59_Y\ : AND2
      port map(A => \I2.N261_0\, B => \I2.N264_0\, Y => 
        \I2.N309_0\);
    
    \I2.OFFSET_37_7l5r\ : MUX2L
      port map(A => \I2.N_680\, B => \I2.N_656\, S => 
        \I2.PIPE7_DTL25R_682\, Y => \I2.N_688\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I179_Y\ : XOR2
      port map(A => \I2.N525_0\, B => 
        \I2.ADD_21x21_fast_I179_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l9r\);
    
    \I1.REG_1_158\ : MUX2H
      port map(A => \REGl257r\, B => \I1.REG_74l257r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_158_net_1\);
    
    \I1.REG_1_277\ : MUX2H
      port map(A => \REGl376r\, B => \I1.REG_74l376r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_277_net_1\);
    
    \I2.STATEe_ns_i_0l1r\ : OA21TTF
      port map(A => \I2.STATEe_ipl3r\, B => \I2.INT_ERRS_net_1\, 
        C => \I2.STATEe_ipl1r\, Y => \I2.STATEe_ns_i_0_il1r\);
    
    \I2.FID_7_0_IVL0R_1733\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl0r_net_1\, 
        Y => \I2.FID_7l0r_adt_net_93569_\);
    
    \I2.LSRAM_IN_404\ : MUX2L
      port map(A => \I2.PIPE5_DTl20r_net_1\, B => 
        \I2.LSRAM_INl20r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_404_net_1\);
    
    \I3.VDBI_57_IVL3R_2256\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854360__net_1\, B
         => \I3.VDBoffl3r_net_1\, Y => 
        \I3.VDBi_57l3r_adt_net_145062_\);
    
    \I1.REG_74_0_IVL352R_1861\ : NOR2FT
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_24_sqmuxa_adt_net_854780__net_1\, Y => 
        \I1.REG_74l352r_adt_net_115945_\);
    
    \I3.VDBi_57_0_ivl29r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l29r_net_1\, C
         => \I3.VDBi_57l29r_adt_net_138175_\, Y => 
        \I3.VDBi_57l29r\);
    
    \I2.ADE_4l15r\ : MUX2L
      port map(A => \I2.RPAGEl15r\, B => \I2.WPAGEl15r_net_1\, S
         => NOESRAME_c, Y => \I2.ADE_4l15r_net_1\);
    
    \I2.DTE_21_1_IV_0_0_18_M7_1215\ : AND2
      port map(A => \I2.DTE_1l18r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35891_\);
    
    \I2.DTO_16_1_iv_0l9r\ : OR2
      port map(A => \I2.DTO_16_1l9r_adt_net_33251_\, B => 
        \I2.DTO_16_1l9r_adt_net_33252_\, Y => \I2.DTO_16_1l9r\);
    
    \I2.un7_tdcgda1_0\ : XOR2
      port map(A => \I2.TDCDASl24r_net_1\, B => \I2.TDCl0r_net_1\, 
        Y => \I2.un7_tdcgda1_0_i_i\);
    
    \I2.G_EVNT_NUMl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_926_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl8r_net_1\);
    
    \I2.STATEE_NSL0R_1026\ : NOR3FFT
      port map(A => BNC_RES_E, B => \I2.STATEe_ipl0r\, C => 
        \I2.INT_ERRS_net_1\, Y => 
        \I2.STATEe_nsl0r_adt_net_23014_\);
    
    \I1.PAGECNT_n8_i_i_x2\ : XOR2
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        B => \I1.N_369\, Y => \I1.N_409_i_i_0_i\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I209_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl13r_adt_net_854940__net_1\, B
         => \I2.PIPE7_DTl13r_net_1\, Y => 
        \I2.SUB_21x21_fast_I209_Y_0\);
    
    \I2.DTO_9_IV_0_O2L0R_1211\ : NOR2
      port map(A => \I2.CRC32_1_SQMUXA_0_38\, B => 
        \I2.DT_SRAML0R_376\, Y => \I2.DTO_9_ivl0r_adt_net_35332_\);
    
    \I2.DTE_21_1_ivl1r\ : AOI21FTT
      port map(A => \I2.DTE_1l1r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, C => 
        \I2.DTE_21_1_iv_2_il1r\, Y => \I2.DTE_21_1_iv_i_0l1r\);
    
    \I3.REG_1l135r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_183_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl135r\);
    
    \I2.L2ARRl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_943_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRl1r_net_1\);
    
    \I2.END_EVNT3\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT3_net_1\);
    
    \I2.PIPE8_DT_21l18r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl18r\, B => 
        \I2.PIPE8_DT_16l18r_net_1\, S => \I2.NWPIPE7_net_1\, Y
         => \I2.PIPE8_DT_21l18r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L0R_2621\ : AND2
      port map(A => \REGl213r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.VDBoffa_31l0r_adt_net_164606_\);
    
    \I2.DTE_1l6r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l6r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l6r_Rd1__net_1\);
    
    NOEAD_pad : OB33PH
      port map(PAD => NOEAD, A => NOEAD_C_I_0_13);
    
    \I2.CRC32_12_I_0_M2L27R_1348\ : AND2
      port map(A => \I2.DT_TEMPl27r_net_1\, B => 
        \I2.N_4667_1_ADT_NET_1046__35\, Y => 
        \I2.N_230_i_i_adt_net_41076_\);
    
    \I2.REG_1l35r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n3_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl35r);
    
    REGl338r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_239_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl338r\);
    
    \I3.PIPEA1l19r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_317_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l19r_net_1\);
    
    \I3.VDBi_57l6r_adt_net_143325_\ : AO21
      port map(A => \I3.N_2037\, B => \I3.N_2269\, C => 
        \I3.VDBi_57l6r_adt_net_143308__net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143325__net_1\);
    
    \I1.REG_1_265\ : MUX2H
      port map(A => \REGl364r\, B => \I1.REG_74l364r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_265_net_1\);
    
    \I5.sstate2se_4_o2\ : NAND2
      port map(A => TICKL0R_557, B => REGl7r, Y => \I5.N_464\);
    
    \I2.SUB9_583\ : MUX2H
      port map(A => \I2.SUB9_i_0_il15r\, B => \I2.SUB9_1l15r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_583_net_1\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2278\ : AND3
      port map(A => REGl48r, B => \I3.N_590\, C => 
        \I3.N_2044_316\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146432_\);
    
    N_1_I3_TCNT3_n7 : XOR2FT
      port map(A => \I3.TCNT3l7r_net_1\, B => \N_1.I3.TCNT3_c6\, 
        Y => \N_1.I3.TCNT3_n7\);
    
    \I2.G_EVNT_NUMl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_929_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl5r_net_1\);
    
    \I3.VDBi_43l10r\ : MUX2L
      port map(A => REGl416r, B => \I3.VDBi_40l10r_net_1\, S => 
        \I3.REGMAPl55r_net_1\, Y => \I3.VDBi_43l10r_net_1\);
    
    \I1.SSTATEL0R_2875\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_ns_il10r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL0R_307\);
    
    \I2.EVNT_WORD_713_1533\ : AND2FT
      port map(A => 
        \I2.WOFFSETl0r_adt_net_854636__adt_net_855712__net_1\, B
         => \I2.N_2864_0_adt_net_854264__net_1\, Y => 
        \I2.EVNT_WORD_713_adt_net_53148_\);
    
    \I2.MIC_ERR_REGS_332\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl4r_net_1\, B => 
        \I2.MIC_ERR_REGSl3r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_332_net_1\);
    
    \I2.FCNT_n1\ : XOR2FT
      port map(A => \I2.N_1236\, B => \I2.N_1237\, Y => 
        \I2.FCNT_n1_net_1\);
    
    \I3.LED_G_0_a3\ : AND2
      port map(A => REGl27r, B => TRM_BUSY_c, Y => LED_G_c);
    
    \I3.VDBi_40_0_i_m2l10r\ : MUX2L
      port map(A => REGl428r, B => REGl444r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_1855\);
    
    \I2.DTE_1l13r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l13r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l13r_Rd1__net_1\);
    
    \I2.PIPE8_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_529_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl1r_net_1\);
    
    \I1.REG_1_242\ : MUX2H
      port map(A => \REGl341r\, B => \I1.REG_74l341r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\, Y => 
        \I1.REG_1_242_net_1\);
    
    \I3.PIPEB_98_2325\ : NOR2FT
      port map(A => \I3.PIPEBl19r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_98_adt_net_159915_\);
    
    \I2.MIC_REG1l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_308_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1l7r_net_1\);
    
    \I2.FID_7_0_IVL28R_979\ : AND2
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl28r_net_1\, 
        Y => \I2.FID_7l28r_adt_net_18739_\);
    
    \I2.UN1_STATE3_0_SQMUXA_1_1061\ : AND3
      port map(A => \I2.un28_sram_empty\, B => 
        \I2.STATE3l5r_net_1\, C => 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26951_\, Y => 
        \I2.L2SERVe_adt_net_26991_\);
    
    \I2.DT_SRAM_0l21r\ : MUX2L
      port map(A => \I2.PIPE10_DTl21r_net_1\, B => 
        \I2.PIPE5_DTL21R_626\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854220__net_1\, Y => 
        \I2.N_889\);
    
    \I2.PIPE6_DT_0_sqmuxa_i_m2\ : MUX2L
      port map(A => LEAD_FLAGl2r, B => LEAD_FLAGl0r, S => 
        \I2.PIPE5_DTL22R_665\, Y => \I2.N_4542\);
    
    \I1.REG_74l308r\ : NAND2FT
      port map(A => \I1.REG_17_sqmuxa\, B => \I1.REG_74_1l308r\, 
        Y => \I1.N_177\);
    
    \I2.OFFSET_37_2l6r\ : MUX2L
      port map(A => \REGl387r\, B => \REGl323r\, S => 
        \I2.PIPE7_DTL27R_67\, Y => \I2.N_649\);
    
    \I2.STATE3_nsl10r\ : AO21
      port map(A => \I2.STATE3l2r_net_1\, B => \I2.N_3016\, C => 
        \I2.N_4676\, Y => \I2.STATE3_nsl10r_net_1\);
    
    \I3.N_57_i_0_0_adt_net_854692_\ : BFR
      port map(A => \I3.N_57_i_0_0_adt_net_854700__net_1\, Y => 
        \I3.N_57_i_0_0_adt_net_854692__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I212_Y\ : XOR2FT
      port map(A => \I2.I180_un1_Y\, B => 
        \I2.SUB_21x21_fast_I212_Y_0\, Y => \I2.SUB8_2_i_i_0l16r\);
    
    \I3.VADm_0_a3l20r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl20r_net_1\, Y => \I3.VADml20r\);
    
    \I2.PIPE6_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_462_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl8r_net_1\);
    
    \I3.VDBi_57_0_ivl11r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855380__net_1\, B => 
        \I3.VDBi_43l11r_net_1\, C => 
        \I3.VDBi_57l11r_adt_net_141441_\, Y => \I3.VDBi_57l11r\);
    
    \I2.DTO_1l14r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l14r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l14r_Rd1__net_1\);
    
    \I1.REG_1_244\ : MUX2H
      port map(A => \REGl343r\, B => \I1.REG_74l343r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_244_net_1\);
    
    \I2.EVNT_WORD_717\ : MUX2H
      port map(A => \I2.EVNT_WORDl4r_net_1\, B => \I2.I_20\, S
         => \I2.N_2864_0_adt_net_854276__net_1\, Y => 
        \I2.EVNT_WORD_717_net_1\);
    
    TDC_RESA_pad : OB33PH
      port map(PAD => TDC_RESA, A => TDC_RES_c_c);
    
    \I2.CRC32_815\ : MUX2L
      port map(A => \I2.CRC32l20r_net_1\, B => \I2.N_3937\, S => 
        \I2.N_2826_1_ADT_NET_794__330\, Y => \I2.CRC32_815_net_1\);
    
    \I2.SUB8_511\ : MUX2H
      port map(A => \I2.SUB8l8r_net_1\, B => \I2.SUB8_2_i_i_0l8r\, 
        S => \I2.SUB8_1_sqmuxa_0_adt_net_855144__net_1\, Y => 
        \I2.SUB8_511_net_1\);
    
    DTO_padl10r : IOB33PH
      port map(PAD => DTO(10), A => \I2.DTO_1l10r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl10r);
    
    \I3.REG_1_ml65r\ : AND2
      port map(A => REGl65r, B => 
        \I3.REGMAPl9r_adt_net_854312__net_1\, Y => 
        \I3.VDBi_20l17r\);
    
    \I3.VDBI_57_0_IVL26R_2152\ : AO21
      port map(A => \I3.VDBil26r_net_1\, B => 
        \I3.N_1910_0_adt_net_854344__net_1\, C => 
        \I3.VDBi_57l26r_adt_net_138571_\, Y => 
        \I3.VDBi_57l26r_adt_net_138577_\);
    
    \I2.WOFFSETl1r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.WOFFSETl1r_adt_net_854992__net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl1r_Rd1__net_1\);
    
    \I2.N_201_adt_net_855048_\ : BFR
      port map(A => \I2.N_201\, Y => 
        \I2.N_201_adt_net_855048__net_1\);
    
    \I3.PIPEA1_305\ : MUX2L
      port map(A => \I3.PIPEA1l7r_net_1\, B => 
        \I3.PIPEA1_12l7r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__254\, Y => 
        \I3.PIPEA1_305_net_1\);
    
    \I3.VDBOFFB_30_IV_0L6R_2381\ : OR2
      port map(A => \I3.VDBoffb_30l6r_adt_net_161981_\, B => 
        \I3.VDBoffb_30l6r_adt_net_161982_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161987_\);
    
    \I2.DT_TEMPl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_778_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl17r_net_1\);
    
    \I3.STATE2l0r_1000\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE2_nsl4r\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.STATE2L0R_378\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I206_Y\ : XOR2
      port map(A => \I2.N501_i\, B => 
        \I2.SUB_21x21_fast_I206_Y_0\, Y => \I2.SUB8_2l10r\);
    
    \I3.VDBi_57_0_iv_0_0_a2l8r_940\ : NOR2
      port map(A => \I3.N_2015_120\, B => \I3.REGMAPL55R_782\, Y
         => \I3.N_2016_318\);
    
    \I3.PIPEA1_12l6r\ : AND2
      port map(A => DPR_cl6r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854508__net_1\, Y => 
        \I3.PIPEA1_12l6r_net_1\);
    
    \I2.PIPE7_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl8r_net_1\);
    
    \I1.SSTATEL9R_2916\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl1r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL9R_433\);
    
    \I3.REG_1L6R_925\ : OA21
      port map(A => \I3.REG1l6r_net_1\, B => \I3.REG2l6r_net_1\, 
        C => \I3.REG3l6r_net_1\, Y => \REGl6r_adt_net_14043_\);
    
    \I2.OFFSET_37_25l4r\ : MUX2L
      port map(A => \REGl257r\, B => \REGl193r\, S => 
        \I2.PIPE7_DTL27R_89\, Y => \I2.N_831\);
    
    \I2.G_EVNT_NUM_n1_i_a2\ : NOR2
      port map(A => \I2.G_EVNT_NUM_i_0_il0r_net_1\, B => 
        \I2.G_EVNT_NUMl1r_net_1\, Y => \I2.N_279\);
    
    \I3.VDBOFFB_30_IV_0L4R_2418\ : OR3
      port map(A => \I3.VDBoffb_30l4r_adt_net_162365_\, B => 
        \I3.VDBoffb_30l4r_adt_net_162359_\, C => 
        \I3.VDBoffb_30l4r_adt_net_162360_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162369_\);
    
    \I2.EVRDYi_496\ : OAI21FTT
      port map(A => EVRDY_c, B => \I2.N_3824_adt_net_90281_\, C
         => \I2.un8_evread_1_adt_net_855796__net_1\, Y => 
        \I2.EVRDYi_496_net_1\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855452_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__292\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\);
    
    \I3.VDBI_57_0_IVL14R_2192\ : AO21
      port map(A => \I3.VDBil14r_net_1\, B => 
        \I3.N_1910_0_adt_net_854348__net_1\, C => 
        \I3.VDBi_57l14r_adt_net_140190_\, Y => 
        \I3.VDBi_57l14r_adt_net_140197_\);
    
    \I3.STATE1l10r\ : DFFS
      port map(CLK => CLK_c, D => \I3.STATE1_nsl0r\, SET => 
        \I3.N_1311_0\, Q => \I3.STATE1l10r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2540\ : AO21
      port map(A => \REGl170r\, B => \I3.REGMAPl18r_net_1\, C => 
        \I3.VDBoffa_31l5r_adt_net_163664_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163693_\);
    
    \I3.REG2_146\ : MUX2L
      port map(A => VDB_inl5r, B => \I3.REG2l5r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG2_146_net_1\);
    
    \I1.REG_74_0_IV_0L173R_2061\ : AND2
      port map(A => \REGl173r\, B => \I1.N_49_267\, Y => 
        \I1.REG_74l173r_adt_net_132940_\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I152_Y_0_1567\ : OAI21
      port map(A => \I2.PIPE4_DTl17r_net_1\, B => 
        \I2.PIPE4_DTl16r_net_1\, C => \I2.RAMDT4l5r_net_1\, Y => 
        \I2.N498_adt_net_56484_\);
    
    \I2.un12_tokoutas_i_0_o2\ : NOR2
      port map(A => \I2.TOKOUTAS_509\, B => \I2.TOKOUT_FL_644\, Y
         => \I2.N_3881\);
    
    \I2.N_4671_adt_net_854596_\ : BFR
      port map(A => \I2.N_4671\, Y => 
        \I2.N_4671_adt_net_854596__net_1\);
    
    REGl378r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_279_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl378r\);
    
    \I1.REG_74_i_o2_0_0_364_m9_i_1\ : AND2
      port map(A => \I1.REG_74_8_308_m9_i_1\, B => 
        \I1.REG_74_i_o2_0_0_364_m9_i_1_adt_net_114039_\, Y => 
        \I1.REG_74_i_o2_0_0_364_m9_i_1_net_1\);
    
    \I2.UN1_STATE1_39_6_1528\ : AO21FTT
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855244__net_1\, 
        B => \I2.STATE1l9r_net_1\, C => \I2.N_3358\, Y => 
        \I2.un1_STATE1_39_6_i_adt_net_52471_\);
    
    \I2.FID_7_0_IVL28R_980\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl76r, C => 
        \I2.FID_7l28r_adt_net_18739_\, Y => 
        \I2.FID_7l28r_adt_net_18747_\);
    
    \I2.PIPE6_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_459_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl5r_net_1\);
    
    TDCDA_padl29r : IB33
      port map(PAD => TDCDA(29), Y => TDCDA_cl29r);
    
    \I3.VDBOFFA_31_IV_0L2R_2596\ : AO21
      port map(A => \REGl183r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.VDBoffa_31l2r_adt_net_164258_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164265_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I5_P0N_i_a4_731\ : OR2
      port map(A => \I2.RAMDT4L12R_143\, B => 
        \I2.PIPE4_DTl5r_adt_net_854416__net_1\, Y => 
        \I2.N_89_0_109\);
    
    \I2.FID_7_0_IVL24R_987\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl24r_net_1\, 
        Y => \I2.FID_7l24r_adt_net_19115_\);
    
    \I2.DTE_21_1_iv_0l16r\ : OR3
      port map(A => \I2.DTE_21_1l16r_adt_net_37823_\, B => 
        \I2.DTE_21_1l16r_adt_net_37833_\, C => 
        \I2.DTE_21_1l16r_adt_net_37834_\, Y => \I2.DTE_21_1l16r\);
    
    \I1.REG_74_0_IVL338R_1878\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l338r_adt_net_117400_\);
    
    \I2.L2TYPE_4_IL12R_1620\ : NAND2FT
      port map(A => \I2.N_4455\, B => \I2.N_4458\, Y => 
        \I2.N_4440_adt_net_67210_\);
    
    \I2.OFFSET_37_12l6r\ : MUX2L
      port map(A => \REGl347r\, B => \I2.N_721\, S => 
        \I2.PIPE7_DTL26R_356\, Y => \I2.N_729\);
    
    \I2.PIPE1_DT_42_1_IVL0R_1521\ : AND2FT
      port map(A => \I2.N_3279_0_adt_net_855232__net_1\, B => 
        \I2.MIC_ERR_REGSl0r_net_1\, Y => 
        \I2.PIPE1_DT_42l0r_adt_net_52239_\);
    
    \I4.END_FLUSH\ : DFFC
      port map(CLK => CLK_c, D => \I4.END_FLUSH_2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => END_FLUSH);
    
    \I2.PIPE6_DT_487\ : MUX2L
      port map(A => \I2.PIPE6_DTl33r_net_1\, B => \I2.N_4526\, S
         => \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_487_net_1\);
    
    \I2.RAMAD1l12r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_666_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l12r_net_1\);
    
    \I2.PIPE5_DT_6l1r\ : MUX2L
      port map(A => \I2.PIPE4_DT_i_il1r_net_1\, B => \I2.N_1070\, 
        S => \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, Y
         => \I2.PIPE5_DT_6l1r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I145_Y_0\ : XOR2
      port map(A => \I2.N_3543_i_i\, B => \I2.G_1_0\, Y => 
        \I2.ADD_18x18_fast_I145_Y_0\);
    
    \I3.VDBI_57_0_IVL29R_2143\ : AND2
      port map(A => \I3.PIPEAl29r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l29r_adt_net_138169_\);
    
    \I3.REG_1_281_e\ : NAND3
      port map(A => \I3.REGMAPl14r_net_1\, B => 
        \I3.STATE1_IPL8R_10\, C => \I3.N_127\, Y => \I3.N_2297_i\);
    
    \I2.PIPE1_DT_42_1_IVL18R_1404\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\, B => 
        \I2.PIPE1_DT_30l18r_net_1\, C => 
        \I2.PIPE1_DT_42l18r_adt_net_47441_\, Y => 
        \I2.PIPE1_DT_42l18r_adt_net_47456_\);
    
    DTE_padl29r : IOB33PH
      port map(PAD => DTE(29), A => \I2.DTE_1l29r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl29r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_a2_3\ : AND2
      port map(A => \I2.RAMDT4L12R_822\, B => 
        \I2.N_139_0_adt_net_55124_\, Y => \I2.N_139_0\);
    
    \I2.PIPE1_DT_42_1_IVL12R_1450\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl8r\, Y => 
        \I2.PIPE1_DT_42l12r_adt_net_49448_\);
    
    REGl173r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_74_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl173r\);
    
    \I3.PIPEA1_318\ : MUX2L
      port map(A => \I3.PIPEA1l20r_net_1\, B => 
        \I3.PIPEA1_12l20r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__251\, Y => 
        \I3.PIPEA1_318_net_1\);
    
    \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672_\ : BFR
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__489\, Y => 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672__net_1\);
    
    \I3.VDBi_340\ : MUX2L
      port map(A => \I3.VDBil0r_net_1\, B => \I3.VDBi_57l0r\, S
         => \I3.un1_STATE1_13_1_adt_net_1351__net_1\, Y => 
        \I3.VDBi_340_net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2597\ : OR2
      port map(A => \I3.VDBoffa_31l2r_adt_net_164261_\, B => 
        \I3.VDBoffa_31l2r_adt_net_164262_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164267_\);
    
    \I2.PIPE6_DT_il33r\ : INV
      port map(A => \I2.PIPE6_DTl33r_net_1\, Y => 
        \I2.PIPE6_DT_il33r_net_1\);
    
    \I2.PIPE10_DT_607\ : MUX2L
      port map(A => \I2.PIPE10_DTl2r_net_1\, B => 
        \I2.PIPE9_DTl2r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_607_net_1\);
    
    \I2.PIPE7_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl5r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl5r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I39_Y\ : AND2
      port map(A => \I2.N241\, B => \I2.N244\, Y => \I2.N304\);
    
    \I2.un1_DTO_cl_0_sqmuxa_0_a2_0_a2_0_a2_0\ : OR3FFT
      port map(A => \I2.STATE2l5r_net_1\, B => 
        \I2.WR_SRAM_2_ADT_NET_748__39\, C => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__181\, Y => 
        \I2.N_2870\);
    
    \I2.TRGCNT_n0_0\ : XOR2
      port map(A => \I2.N_3794\, B => \I2.TRGCNTl0r_net_1\, Y => 
        \I2.TRGCNT_n0_0_net_1\);
    
    \I2.DTOSl29r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl29r, Q => 
        \I2.DTOSl29r_net_1\);
    
    \I3.un211_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_558\, B => \I3.N_586\, Y => 
        \I3.un211_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.ROFFSETl3r_1510\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_915_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETL3R_617\);
    
    \I3.un60_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_632\, B => \I3.un60_reg_ads_3\, Y => 
        \I3.un60_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.CRC32l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_800_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l5r_net_1\);
    
    \I3.VDBil11r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_351_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil11r_net_1\);
    
    \I2.PIPE4_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl26r_net_1\);
    
    REGl291r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_192_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl291r\);
    
    \I1.REG_74_8_0_o4_a0_0l324r_721\ : OR2
      port map(A => \I1.PAGECNTL5R_309\, B => \I1.PAGECNTL6R_248\, 
        Y => \I1.REG_74_1_A0_0L228R_99\);
    
    \I2.STATEe_nsl4r\ : AO21
      port map(A => \I2.STATEe_ipl2r\, B => \I2.N_3510\, C => 
        \I2.STATEe_nsl4r_adt_net_22922_\, Y => 
        \I2.STATEe_nsl4r_net_1\);
    
    \I3.RAMDTSl11r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl11r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl11r_net_1\);
    
    \I2.FID_7_0_iv_0l1r\ : OAI21FTF
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl1r_net_1\, 
        C => \I2.FID_7_0_iv_0l1r_adt_net_93441_\, Y => 
        \I2.FID_7_0_iv_0l1r_net_1\);
    
    \I3.PIPEB_4l28r\ : NAND2FT
      port map(A => DPR_cl28r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855280__net_1\, 
        Y => \I3.PIPEB_4l28r_net_1\);
    
    \I3.un106_reg_ads_0_a2_0_a2_0\ : NOR2FT
      port map(A => \I3.VASl12r_net_1\, B => \I3.N_547_369\, Y
         => \I3.N_548\);
    
    \I3.VDBi_57_0_iv_0_0_a2l13r_744\ : NAND2FT
      port map(A => \I3.REGMAPL16R_444\, B => \I3.N_354_0_130\, Y
         => \I3.N_2014_122\);
    
    \I3.PIPEA_8_0l23r\ : MUX2L
      port map(A => DPR_cl23r, B => \I3.PIPEA1l23r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855360__net_1\, Y => \I3.N_232\);
    
    \I2.un7_bnc_id_1_I_24\ : XOR2
      port map(A => \I2.BNC_IDl5r_net_1\, B => \I2.N_34_0\, Y => 
        \I2.I_24_0\);
    
    \I2.SRAM_EVNT_n2\ : XOR2
      port map(A => \I2.N_3826\, B => \I2.SRAM_EVNT_n2_0_net_1\, 
        Y => \I2.SRAM_EVNT_n2_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2392\ : AO21
      port map(A => \REGl322r\, B => \I3.REGMAPl37r_net_1\, C => 
        \I3.VDBoffb_30l5r_adt_net_162128_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162169_\);
    
    \I1.sstatel8r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl2r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel8r_net_1\);
    
    \I4.un4_bcnt_I_5\ : XOR2
      port map(A => \I4.bcntl1r_net_1\, B => \I4.bcntl0r_net_1\, 
        Y => \I4.I_5\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854456_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854472__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854456__net_1\);
    
    \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m3_860\ : MUX2H
      port map(A => \I2.MIC_REG2L3R_ADT_NET_834020_RD1__215\, B
         => \I2.MIC_REG3L3R_804\, S => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Rd1__net_1\, Y => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_M3_238\);
    
    \I2.PIPE5_DT_677\ : MUX2L
      port map(A => \I2.PIPE5_DTl1r_net_1\, B => 
        \I2.PIPE5_DT_6l1r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_677_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I0_S_0_x2\ : XOR2
      port map(A => \I2.RAMDT4l0r_net_1\, B => 
        \I2.PIPE4_DTl0r_net_1\, Y => \I2.un27_pipe5_dt0l0r\);
    
    \I2.un2_evnt_word_I_48\ : AND2
      port map(A => \I2.WOFFSETl7r\, B => \I2.N_29\, Y => 
        \I2.DWACT_FINC_E_0l4r\);
    
    \I3.PIPEA_8_0l3r\ : MUX2L
      port map(A => DPR_cl3r, B => \I3.PIPEA1l3r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855364__net_1\, Y => \I3.N_212\);
    
    \I2.N_4539_i_0_o2\ : NOR2FT
      port map(A => \I2.PIPE5_DTL23R_624\, B => 
        \I2.PIPE5_DTL21R_894\, Y => \I2.N_215\);
    
    \I2.PIPE6_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_474_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl20r_net_1\);
    
    \I2.STATE1_ns_il5r\ : NOR2
      port map(A => \I2.CHAINA_EN244_i_adt_net_855264__net_1\, B
         => \I2.N_3287_i_0\, Y => \I2.STATE1_ns_il5r_net_1\);
    
    \I1.ISI_0_sqmuxa_1_0_i_o2\ : NAND2
      port map(A => \I1.sstatel9r_net_1\, B => \I1.N_321\, Y => 
        \I1.N_346\);
    
    \I3.VDBI_57_0_IV_0_0L15R_2183\ : AND2
      port map(A => \I3.PIPEAl15r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l15r_adt_net_139959_\);
    
    \I2.PIPE9_DT_289\ : MUX2L
      port map(A => \I2.PIPE9_DTl20r_net_1\, B => 
        \I2.PIPE8_DTl20r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_289_net_1\);
    
    \I2.STATE3_ns_o3_0l12r\ : NAND2FT
      port map(A => \I2.FIFO_FULL_592\, B => NOESRAME_C_833, Y
         => \I2.N_3015\);
    
    \I2.STATE2_ns_0l4r\ : NAND2FT
      port map(A => \I2.N_2864_0_adt_net_835284_Rd1__net_1\, B
         => \I2.N_4293_Rd1__net_1\, Y => \I2.STATE2l1r\);
    
    \I3.VDBOFFB_30_IV_0L1R_2461\ : AND2
      port map(A => \REGl310r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        Y => \I3.VDBoffb_30l1r_adt_net_162904_\);
    
    \I2.N479_adt_net_296182_\ : NOR2FT
      port map(A => \I2.N363\, B => \I2.N356\, Y => 
        \I2.N479_adt_net_296182__net_1\);
    
    \I2.OFFSETl7r_1564\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_567_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL7R_671\);
    
    \I3.STATE1l9r_1165\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL9R_427\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854588_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854588__net_1\);
    
    \I2.N_4646_1_ADT_NET_19637_RD1__2976\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_19637_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_19637_RD1__523\);
    
    \I3.VDBOFFA_31_IV_0L7R_2503\ : AO21
      port map(A => \REGl260r\, B => \I3.REGMAPl29r_net_1\, C => 
        \I3.VDBoffa_31l7r_adt_net_163280_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163312_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I44_Y\ : AND2
      port map(A => \I2.G_1_2\, B => \I2.N309_adt_net_70030_\, Y
         => \I2.N309\);
    
    DPR_padl20r : IB33
      port map(PAD => DPR(20), Y => DPR_cl20r);
    
    \I2.END_CHAINA1_708_1539\ : AO21
      port map(A => \I2.END_CHAINA1_net_1\, B => \I2.N_3288\, C
         => \I2.END_CHAINA1_708_adt_net_53509_\, Y => 
        \I2.END_CHAINA1_708_adt_net_53513_\);
    
    \I2.PIPE10_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_608_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl3r_net_1\);
    
    \I3.VDBI_57_IVL4R_2250\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854360__net_1\, B
         => \I3.VDBoffl4r_net_1\, Y => 
        \I3.VDBi_57l4r_adt_net_144429_\);
    
    \I3.REGMAPl6r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un29_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl6r_net_1\);
    
    TRM_DRDY_pad : OB33PH
      port map(PAD => TRM_DRDY, A => EVRDY_c);
    
    \I2.CRC32l11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_806_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l11r_net_1\);
    
    \I2.DT_TEMP_7l29r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854232__net_1\, B => 
        \I2.DT_SRAMl29r_net_1\, Y => \I2.DT_TEMP_7l29r_net_1\);
    
    \I1.REG_74_0_ivl238r\ : AO21
      port map(A => \REGl238r\, B => \I1.N_113\, C => 
        \I1.REG_74l238r_adt_net_126899_\, Y => \I1.REG_74l238r\);
    
    \I5.SBYTEl7r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_72_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl7r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I174_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l11r_net_1\, B => 
        \I2.PIPE4_DTl4r_net_1\, Y => 
        \I2.ADD_21x21_fast_I174_Y_0_0\);
    
    \I2.REG_1_c7_i\ : AO21
      port map(A => REGl39r, B => 
        \I2.N_3836_i_0_adt_net_2390__net_1\, C => 
        \I2.N_3836_i_0_adt_net_101388_\, Y => \I2.N_3836_i_0\);
    
    \I2.REG_0l3r_adt_net_848__adt_net_854216_\ : BFR
      port map(A => 
        \I2.REG_0l3r_adt_net_848__adt_net_854228__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__adt_net_854216__net_1\);
    
    \I2.SUB8_513\ : MUX2H
      port map(A => \I2.SUB8l10r_net_1\, B => \I2.SUB8_2l10r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855144__net_1\, Y => 
        \I2.SUB8_513_net_1\);
    
    \I5.un1_sdab_0_a2\ : NOR2FT
      port map(A => \I5.CHAIN_SELECT_net_1\, B => 
        \I5.SDAnoe_net_1\, Y => un1_sdab_0_a2);
    
    \I2.CRC32_12_i_m2l8r\ : MUX2H
      port map(A => \I2.DT_SRAMl8r_net_1\, B => 
        \I2.DT_TEMPl8r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854436__net_1\, Y => 
        \I2.N_3956_i_i\);
    
    \I2.un78_pipe5_dt_0\ : XOR2
      port map(A => \I2.RAMDT4l7r_net_1\, B => 
        \I2.RAMDT4l13r_net_1\, Y => \I2.un78_pipe5_dt_0_net_1\);
    
    \I2.EVNT_REJ_2_sqmuxa\ : AND2
      port map(A => \I2.un28_sram_empty\, B => 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26951_\, Y => 
        \I2.EVNT_REJ_2_sqmuxa_net_1\);
    
    \I2.BNCID_VECTrff_14_251_0\ : AO21
      port map(A => \I2.BNCID_VECTwa14_1_net_1\, B => 
        \I2.BNCID_VECTrff_12_253_0_a2_0\, C => 
        \I2.BNCID_VECTro_14\, Y => 
        \I2.BNCID_VECTrff_14_251_0_net_1\);
    
    \I2.PIPE4_DTL10R_3087\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL10R_851\);
    
    \I3.PIPEA1_312\ : MUX2L
      port map(A => \I3.PIPEA1l14r_net_1\, B => 
        \I3.PIPEA1_12l14r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__253\, Y => 
        \I3.PIPEA1_312_net_1\);
    
    \I2.PIPE4_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl21r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl21r_net_1\);
    
    \I1.NOELUTi\ : DFFS
      port map(CLK => CLK_c, D => \I1.NOELUTi_51_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => NOELUT_c);
    
    \I3.TCNT1_c3\ : AND2
      port map(A => \I3.TCNT1_i_0_il3r_net_1\, B => 
        \I3.TCNT1_c2_net_1\, Y => \I3.TCNT1_c3_net_1\);
    
    \I2.un1_STATE2_15_i_0_o2\ : NOR2
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__181\, B => 
        \I2.N_4184\, Y => \I2.N_4282\);
    
    \I3.VDBOFFA_31_IV_0L4R_2552\ : AND2
      port map(A => \REGl169r\, B => \I3.REGMAPl18r_net_1\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163858_\);
    
    \I1.REG_74_0_ivl386r\ : AO21
      port map(A => \REGl386r\, B => \I1.N_257\, C => 
        \I1.REG_74l386r_adt_net_111491_\, Y => \I1.REG_74l386r\);
    
    \I1.REG_74_0_ivl348r\ : AO21
      port map(A => \REGl348r\, B => \I1.N_217\, C => 
        \I1.REG_74l348r_adt_net_116326_\, Y => 
        \I1.REG_74l348r_net_1\);
    
    \I2.TEMPF_adt_net_855740__adt_net_855896_\ : BFR
      port map(A => \I2.TEMPF_adt_net_855740__net_1\, Y => 
        \I2.TEMPF_adt_net_855740__adt_net_855896__net_1\);
    
    \I3.VDBI_57_IV_0_0_O2_0_8_TZL0R_2271\ : AO21
      port map(A => EVRDY_c, B => \I3.N_2053\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_adt_net_146105_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_adt_net_146111_\);
    
    \I2.LEAD_FLAG6_7_i_0_o2l7r\ : OAI21FTF
      port map(A => \I2.NWPIPE5_net_1\, B => 
        \I2.PIPE5_DTL30R_622\, C => \I2.N_222_adt_net_63455_\, Y
         => \I2.N_222\);
    
    \I3.REG_1_214\ : MUX2L
      port map(A => VDB_inl1r, B => REGl407r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_214_0\);
    
    \I3.REG_1l149r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_197_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl149r\);
    
    \I1.sstate_tr18_0_a2_0_a2\ : NAND2FT
      port map(A => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854912__net_1\, B
         => \I1.N_598\, Y => \I1.N_604\);
    
    \I2.L2TYPEl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_592_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl3r_net_1\);
    
    \I2.TDCl2r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TDC_652_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TDCl2r_net_1\);
    
    \I1.REG_74l356r\ : NAND3FFT
      port map(A => \I1.N_41_9_adt_net_854784__net_1\, B => 
        \I1.REG_23_sqmuxa\, C => \I1.REG_74_0l348r\, Y => 
        \I1.N_225\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I163_Y\ : AND2FT
      port map(A => \I2.I163_un1_Y\, B => 
        \I2.N492_i_adt_net_89450_\, Y => \I2.N492_i\);
    
    \I2.LSRAM_IN_387\ : MUX2L
      port map(A => \I2.PIPE5_DTl3r_net_1\, B => 
        \I2.LSRAM_INl3r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_387_net_1\);
    
    \I5.SDANOE_8_0_915\ : NOR3FFT
      port map(A => \I5.SDAnoe_net_1\, B => 
        \I5.SDAnoe_8_adt_net_9736_\, C => \I5.sstate1l6r_net_1\, 
        Y => \I5.SDAnoe_8_adt_net_9738_\);
    
    \I2.PIPE10_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_611_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl6r_net_1\);
    
    \I2.CRC32_12_il4r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_118_i_i_0\, Y => 
        \I2.N_3921\);
    
    \I2.ROFFSET_n10\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\, B => 
        \I2.ROFFSET_n10_tz_i\, Y => \I2.ROFFSET_n10_net_1\);
    
    \I1.REG_74_0_IVL378R_1821\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l378r_adt_net_112657_\);
    
    \I2.DTE_21_1_IVL14R_1282\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l14r\, C
         => \I2.DTE_21_1l14r_adt_net_38070_\, Y => 
        \I2.DTE_21_1l14r_adt_net_38071_\);
    
    \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__3007\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854852__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__761\);
    
    \I3.PIPEBl31r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_110_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEB_i_0_il31r\);
    
    \I1.REG_74_0_ivl403r\ : AO21
      port map(A => \REGl403r\, B => \I1.N_273\, C => 
        \I1.REG_74l403r_adt_net_109842_\, Y => \I1.REG_74l403r\);
    
    \I5.sstate1se_6_i_0_m4\ : MUX2L
      port map(A => \I5.sstate1l7r_net_1\, B => 
        \I5.sstate1l6r_net_1\, S => TICKL0R_558, Y => \I5.N_98\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I62_Y_1678\ : AND2FT
      port map(A => \I2.LSRAM_OUTl8r\, B => \I2.PIPE7_DTL8R_697\, 
        Y => \I2.N312_0_adt_net_86450_\);
    
    \I2.RAMAD1_654\ : MUX2L
      port map(A => \I2.RAMAD1_12l0r_net_1\, B => 
        \I2.RAMAD1l0r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__169\, Y => 
        \I2.RAMAD1_654_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I177_Y_2680\ : OR3
      port map(A => \I2.N298_0\, B => 
        \I2.N477_adt_net_302175__net_1\, C => 
        \I2.N477_adt_net_302179__net_1\, Y => 
        \I2.N477_adt_net_371301_\);
    
    \I3.REG_1l55r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_156_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl55r);
    
    \I3.STATE1_ns_0_iv_0_0l7r\ : AO21
      port map(A => \I3.un1_REGMAP_34\, B => 
        \I3.STATE1_nsl7r_adt_net_136177_\, C => 
        \I3.STATE1_nsl7r_adt_net_136170_\, Y => \I3.STATE1_nsl7r\);
    
    \I3.VDBi_16_i_m2l5r\ : MUX2L
      port map(A => REGl37r, B => \I3.N_283\, S => 
        \I3.REGMAPl7r_net_1\, Y => \I3.N_282_i_i\);
    
    \I2.DTE_0_sqmuxa_i_0_m2_1\ : NOR2
      port map(A => \I2.WOFFSETl0r_adt_net_854640__net_1\, B => 
        \I2.N_223_156\, Y => \I2.DTE_0_sqmuxa_i_0_N_3_1\);
    
    \I3.un231_reg_ads_0_a2_4_a3\ : NOR3
      port map(A => \I3.N_547\, B => \I3.N_554\, C => 
        \I3.un231_reg_ads_1\, Y => 
        \I3.un231_reg_ads_0_a2_4_a3_net_1\);
    
    DTO_padl0r : IOB33PH
      port map(PAD => DTO(0), A => \I2.DTO_1l0r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl0r);
    
    \I2.un1_STATE3_0_sqmuxa_1\ : OR2
      port map(A => \I2.N_1170_adt_net_1217__net_1\, B => 
        \I2.L2SERVe_adt_net_26991_\, Y => \I2.L2SERVe\);
    
    \I5.REG_1_42\ : MUX2L
      port map(A => \I5.SENS_ADDRl1r_net_1\, B => REGl429r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_42_net_1\);
    
    \I1.REG_74_0_IV_I_A2L211R_2023\ : AND2
      port map(A => \REGl211r\, B => \I1.N_183_i_0\, Y => 
        \I1.N_144_adt_net_129587_\);
    
    \I2.OFFSET_37_22l6r\ : MUX2L
      port map(A => \REGl243r\, B => \REGl179r\, S => 
        \I2.PIPE7_DTL27R_77\, Y => \I2.N_809\);
    
    \I2.ADOl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl8r);
    
    \I1.REG_74_0_ivl378r\ : AO21
      port map(A => \REGl378r\, B => \I1.N_249\, C => 
        \I1.REG_74l378r_adt_net_112657_\, Y => \I1.REG_74l378r\);
    
    \I2.STATE1_1_sqmuxa_5_0_a2_0\ : NAND2FT
      port map(A => \I2.CHAINA_EN244_i_adt_net_855260__net_1\, B
         => \I2.N_3881\, Y => \I2.END_CHAINA1_1_sqmuxa_3\);
    
    \I2.CRC32l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_802_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l7r_net_1\);
    
    \I2.EVNT_NUM_80\ : NAND2FT
      port map(A => EV_RES_C_569, B => \I2.EVNT_NUMl0r_net_1\, Y
         => \I2.N_1211\);
    
    \I2.N_70_adt_net_54406_\ : AOI21
      port map(A => \I2.PIPE4_DTL10R_475\, B => 
        \I2.PIPE4_DTL9R_471\, C => \I2.RAMDT4L5R_137\, Y => 
        \I2.N_70_adt_net_54406__net_1\);
    
    VDB_padl2r : IOB33PH
      port map(PAD => VDB(2), A => \I3.VDBml2r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl2r);
    
    \I2.ROFFSETe_0_o3_i_a3\ : NOR2FT
      port map(A => \I2.FIFO_FULL_net_1\, B => 
        \I2.STATE3_0_sqmuxa_1_0\, Y => \I2.N_145\);
    
    NWRSRAME_pad : OB33PH
      port map(PAD => NWRSRAME, A => NWRSRAME_c);
    
    \I3.PIPEA_8_0l2r\ : MUX2L
      port map(A => DPR_cl2r, B => \I3.PIPEA1l2r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855364__net_1\, Y => \I3.N_211\);
    
    \I1.REG_74_0_IVL169R_2065\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l169r_adt_net_133321_\);
    
    \I2.un1_STATE1_23\ : NOR2
      port map(A => \I2.STATE1l11r_net_1\, B => 
        \I2.END_TDC1_0_sqmuxa_1_net_1\, Y => 
        \I2.un1_STATE1_23_net_1\);
    
    \I3.VDBml20r\ : MUX2L
      port map(A => \I3.VDBil20r_net_1\, B => \I3.N_162\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml20r_net_1\);
    
    \I3.VDBml19r\ : MUX2L
      port map(A => \I3.VDBil19r_net_1\, B => \I3.N_161\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml19r_net_1\);
    
    \I3.UN10_TCNT2_2105\ : OR2
      port map(A => \I3.TCNT2_i_0_il4r_net_1\, B => 
        \I3.TCNT2l3r_net_1\, Y => \I3.un10_tcnt2_adt_net_135286_\);
    
    \I2.END_EVNT9\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT8_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT9_net_1\);
    
    \I2.STATE1_ns_i_o3l9r\ : OR2FT
      port map(A => \I2.STATE1L10R_590\, B => \I2.N_3272_344\, Y
         => \I2.N_3288\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I70_Y\ : AOI21
      port map(A => \I2.N246_0\, B => \I2.N242\, C => \I2.N245\, 
        Y => \I2.N320\);
    
    \I2.NWPIPE9_0\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE8_i_0_i_0_0\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE9_0_net_1\);
    
    \I1.REG_74_0_IVL331R_1885\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l331r_adt_net_118002_\);
    
    \I3.STATE2l3r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.STATE2_ns_i_i_a5_0_a3l1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.STATE2l3r_net_1\);
    
    \I2.DTE_1_843\ : MUX2L
      port map(A => \I2.DTE_1l3r_net_1\, B => 
        \I2.DTE_21_1_iv_i_0l3r\, S => \I2.N_2868_1\, Y => 
        \I2.DTE_1_843_net_1\);
    
    \I2.NWPIPE4_1469\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE3_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE4_576\);
    
    \I2.PIPE5_DT_696\ : MUX2L
      port map(A => \I2.PIPE5_DTl20r_net_1\, B => 
        \I2.PIPE5_DT_6l20r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_696_net_1\);
    
    \I2.RAMAD_4_0l11r\ : MUX2H
      port map(A => \I2.RAMAD1l11r_net_1\, B => RAMAD_VMEl11r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_538\);
    
    FID_padl24r : OB33PH
      port map(PAD => FID(24), A => FID_cl24r);
    
    \I3.VDBi_31l9r\ : MUX2L
      port map(A => \I3.REGl142r\, B => \I3.VDBi_29l9r\, S => 
        \I3.REGMAPl17r_adt_net_854288__net_1\, Y => 
        \I3.VDBi_31l9r_net_1\);
    
    \I3.VDBI_57_0_IV_0L27R_2147\ : NOR2FT
      port map(A => \I3.REGl160r\, B => 
        \I3.N_1917_adt_net_855336__net_1\, Y => 
        \I3.VDBi_57l27r_adt_net_138431_\);
    
    \I2.I_1336_ca_0_and2\ : AND2FT
      port map(A => \I2.OFFSETL1R_680\, B => \I2.SUB8L4R_708\, Y
         => \I2.ca_0_and2\);
    
    \I1.REG_74_12_348_m9_i_o7\ : NOR2
      port map(A => \I1.PAGECNTL7R_525\, B => \I1.PAGECNTL6R_836\, 
        Y => \I1.REG_74_1_380_N_16\);
    
    \I3.PIPEA_8_0l4r\ : MUX2L
      port map(A => DPR_cl4r, B => \I3.PIPEA1l4r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855364__net_1\, Y => \I3.N_213\);
    
    TDCDA_padl0r : IB33
      port map(PAD => TDCDA(0), Y => TDCDA_cl0r);
    
    \I2.REG_1_c5_i\ : OAI21FTF
      port map(A => \I2.un8_evread_1_adt_net_855784__net_1\, B
         => \I2.N_124\, C => \I2.N_3834_i_0_adt_net_101432_\, Y
         => \I2.N_3834_i_0\);
    
    \I2.OFFSET_37_16l3r\ : MUX2L
      port map(A => \REGl264r\, B => \REGl200r\, S => 
        \I2.PIPE7_DTL27R_81\, Y => \I2.N_758\);
    
    \I2.N_4283_i_0_a2_m1_e_0_664\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__47\, B => 
        \I2.TEMPF_adt_net_855740__net_1\, Y => \I2.N_4283_I_0_42\);
    
    \I2.SUB9_1_ADD_18x18_fast_I59_Y\ : NAND2
      port map(A => \I2.N292\, B => \I2.N296\, Y => \I2.N327\);
    
    \I1.REG_74_0_iv_0_o2l253r\ : AND3
      port map(A => \I1.N_232_1\, B => \I1.N_395_adt_net_113232_\, 
        C => \I1.N_395_adt_net_113231_\, Y => \I1.N_395\);
    
    \I2.RAMDT4l13r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl13r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l13r_net_1\);
    
    \I3.REGMAPl9r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un41_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPl9r_net_1\);
    
    \I2.FCNTl2r_1493_1786\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_945_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.FCNTL2R_892\);
    
    \I3.LWORDS_3034\ : DFFC
      port map(CLK => CLK_c, D => \I3.LWORDS_61_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.LWORDS_788\);
    
    \I2.PIPE1_DT_42_1_IVL4R_1497\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855032__net_1\, 
        B => \I2.PIPE1_DT_12l4r_net_1\, Y => 
        \I2.PIPE1_DT_42l4r_adt_net_51418_\);
    
    \I2.BNCID_VECT_tile_0_DOUTl3r\ : MUX2L
      port map(A => \I2.DIN_REG1l3r\, B => \I2.DOUT_TMPl3r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl11r\);
    
    \I1.N_137_adt_net_854764_\ : BFR
      port map(A => \I1.N_137\, Y => 
        \I1.N_137_adt_net_854764__net_1\);
    
    \I2.PIPE9_DT_280\ : MUX2L
      port map(A => \I2.PIPE9_DTl11r_net_1\, B => 
        \I2.PIPE8_DTl11r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_280_net_1\);
    
    \I1.REG_74_0_iv_i_a2_il205r\ : AO21
      port map(A => \REGl205r\, B => \I1.N_183_i_0\, C => 
        \I1.N_280_adt_net_130103_\, Y => \I1.N_280\);
    
    \I2.resyn_0_I2_TRGCNT_c0_i\ : AOI21
      port map(A => \I2.N_3794\, B => \I2.un9_tdctrgi_i_0\, C => 
        \I2.TRGCNTl0r_net_1\, Y => \I2.N_3761\);
    
    \I5.BITCNTe_0_a2_0\ : OR2FT
      port map(A => \I5.N_130\, B => \I5.BITCNTe_adt_net_9456_\, 
        Y => \I5.BITCNTe\);
    
    \I3.REG_1_190\ : MUX2L
      port map(A => VDB_inl9r, B => \I3.REGl142r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, Y => 
        \I3.REG_1_190_0\);
    
    \I3.REGMAPl57r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un231_reg_ads_0_a2_4_a3_net_1\, Q => 
        \I3.REGMAPl57r_net_1\);
    
    \I2.CRC32_12_il15r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_113_i_i_0\, Y => 
        \I2.N_3932\);
    
    \I3.WRITES_1162\ : DFFC
      port map(CLK => CLK_c, D => \I3.WRITES_23_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.WRITES_424\);
    
    \I2.STATEel1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATEe_nsl3r_net_1\, CLR
         => \I2.STATEe_i_0l0r_net_1\, Q => \I2.STATEe_ipl1r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I110_Y\ : AND2FT
      port map(A => \I2.I110_un1_Y\, B => 
        \I2.N442_i_adt_net_71348_\, Y => \I2.N442_i\);
    
    \I2.PIPE9_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_295_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl26r_net_1\);
    
    \I2.WOFFSET_832\ : MUX2L
      port map(A => \I2.WOFFSETl5r_Rd1__net_1\, B => 
        \I2.N_4248_Rd1__net_1\, S => 
        \I2.N_2828_ADT_NET_1062__ADT_NET_835308_RD1__757\, Y => 
        \I2.WOFFSETl5r\);
    
    \I2.PIPE4_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl27r_net_1\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2518\ : AO21
      port map(A => \REGl195r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.N_2070_adt_net_163458_\, Y => 
        \I3.N_2070_adt_net_163499_\);
    
    TRM_BUSY_pad : OB33PH
      port map(PAD => TRM_BUSY, A => TRM_BUSY_c);
    
    \I1.REG_1_227\ : MUX2H
      port map(A => \REGl326r\, B => \I1.REG_74l326r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y => 
        \I1.REG_1_227_net_1\);
    
    \I2.PIPE1_DTl1r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_728_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl1r_net_1\);
    
    DTO_padl15r : IOB33PH
      port map(PAD => DTO(15), A => \I2.DTO_1l15r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl15r);
    
    \I2.SUB9_1_ADD_18x18_fast_I7_P0N\ : OR2FT
      port map(A => \I2.SUB8l11r_net_1\, B => \I2.N_3547_i_i\, Y
         => \I2.N247\);
    
    \I2.DTE_21_1l14r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l14r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l14r_Rd1__net_1\);
    
    FID_padl16r : OB33PH
      port map(PAD => FID(16), A => FID_cl16r);
    
    \I2.DTO_1l30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_904_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l30r_net_1\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__3052\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__806\);
    
    \I2.DT_SRAMl0r\ : MUX2L
      port map(A => \I2.N_868\, B => \I2.PIPE2_DTl0r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl0r_net_1\);
    
    \I2.CRC32_12_i_0_a2_1l6r_960\ : AND2
      port map(A => \I2.STATE2L0R_588\, B => 
        \I2.WR_SRAM_2_ADT_NET_748__39\, Y => \I2.N_2867_1_338\);
    
    \I3.REG3l3r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG3_128_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l3r_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I120_Y_0_1586\ : AO21
      port map(A => 
        \I2.PIPE4_DTl5r_adt_net_854412__adt_net_855600__net_1\, B
         => \I2.PIPE4_DTl6r_net_1\, C => \I2.RAMDT4L5R_821\, Y
         => \I2.N531_adt_net_59960_\);
    
    \I3.TCNT3_378\ : MUX2H
      port map(A => \I3.TCNT3l1r_net_1\, B => \I3.TCNT3_n1_net_1\, 
        S => \TICKl1r\, Y => \I3.TCNT3_378_net_1\);
    
    \I5.PULSE_FL_1465\ : DFFC
      port map(CLK => CLK_c, D => \I5.PULSE_FL_53_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.PULSE_FL_572\);
    
    \I3.TCNT1_n2\ : XOR2
      port map(A => \I3.TCNT1l2r_net_1\, B => \I3.TCNT1_c1_net_1\, 
        Y => \I3.TCNT1_n2_net_1\);
    
    \I3.VDBm_0l6r\ : MUX2L
      port map(A => \I3.PIPEAl6r_net_1\, B => \I3.PIPEBl6r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_148\);
    
    \I3.REG_1_206\ : MUX2L
      port map(A => VDB_inl25r, B => \I3.REGl158r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\, Y => 
        \I3.REG_1_206_0\);
    
    \I2.PIPE1_DT_42_1_iv_1l1r\ : NAND2FT
      port map(A => \I2.N_12169_i_adt_net_20407_\, B => 
        \I2.N_3254\, Y => \I2.N_12169_i\);
    
    \I2.un1_DTO_cl_0_sqmuxa_0_a2_1_a2_0_a2_0\ : NAND2FT
      port map(A => \I2.WOFFSETl0r_adt_net_854648__net_1\, B => 
        \I2.STATE2l2r_net_1\, Y => \I2.DTO_cl_0_sqmuxa_0\);
    
    \I3.VDBOFFA_31_IV_0L7R_2506\ : AO21
      port map(A => \REGl236r\, B => \I3.REGMAPl26r_net_1\, C => 
        \I3.VDBoffa_31l7r_adt_net_163308_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163315_\);
    
    \I2.MIC_ERR_REGS_360\ : MUX2H
      port map(A => \I2.MIC_ERR_REGSl31r_net_1\, B => 
        \I2.MIC_ERR_REGSl32r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_360_net_1\);
    
    \I2.DTE_21_1l12r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l12r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l12r_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2583\ : AND2
      port map(A => \REGl239r\, B => \I3.REGMAPl27r_net_1\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164218_\);
    
    \I2.OFFSET_37_17l4r\ : MUX2L
      port map(A => \I2.N_759\, B => \I2.N_751\, S => 
        \I2.PIPE7_DTL26R_353\, Y => \I2.N_767\);
    
    \I1.N_50_0_ADT_NET_1409__2884\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__200\, B => 
        \I1.N_50_0_adt_net_109751__net_1\, Y => 
        \I1.N_50_0_ADT_NET_1409__320\);
    
    \I2.PIPE1_DT_755\ : MUX2L
      port map(A => \I2.PIPE1_DTl28r_net_1\, B => 
        \I2.PIPE1_DT_42l28r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854560__net_1\, 
        Y => \I2.PIPE1_DT_755_net_1\);
    
    \I2.STATE1l7r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl11r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE1l7r_net_1\);
    
    \I3.RAMAD_VMEl8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_32_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl8r);
    
    \I1.REG_74_0_ivl341r\ : AO21
      port map(A => \REGl341r\, B => \I1.N_217\, C => 
        \I1.REG_74l341r_adt_net_116928_\, Y => \I1.REG_74l341r\);
    
    \I2.FID_7_0_ivl5r\ : OA21FTF
      port map(A => \I2.STATE3l2r_net_1\, B => \I2.DTOSl5r_net_1\, 
        C => \I2.FID_7_0_iv_0l5r_net_1\, Y => 
        \I2.FID_7_0_ivl5r_net_1\);
    
    \I2.DT_SRAM_0l14r\ : MUX2L
      port map(A => \I2.PIPE10_DTl14r_net_1\, B => 
        \I2.PIPE5_DTl14r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, Y => 
        \I2.N_882\);
    
    \I2.PIPE10_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_633_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl28r_net_1\);
    
    \I2.RAMDT4L12R_3045\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_799\);
    
    \I2.N_4667_1_ADT_NET_1046__2759\ : OAI21FTF
      port map(A => \I2.N_4261_302\, B => \I2.N_4283_I_0_45\, C
         => \I2.STATE2L2R_589\, Y => 
        \I2.N_4667_1_ADT_NET_1046__35\);
    
    \I1.PAGECNT_n8_i_i_o2\ : NAND2
      port map(A => \I1.PAGECNTl7r_net_1\, B => \I1.N_345\, Y => 
        \I1.N_369\);
    
    \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876_\ : BFR
      port map(A => \I5.REG_2_sqmuxa_0_adt_net_975__net_1\, Y => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\);
    
    \I2.STATE1l12r_adt_net_855184_\ : BFR
      port map(A => \I2.STATE1L12R_646\, Y => 
        \I2.STATE1l12r_adt_net_855184__net_1\);
    
    N_1_I3_TCNT3_373 : MUX2H
      port map(A => \I3.TCNT3_i_0_il6r_net_1\, B => 
        \N_1.I3.TCNT3_n6\, S => \TICKl1r\, Y => TCNT3_373);
    
    \I2.LSRAM_INl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_398_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl14r_net_1\);
    
    \I1.REG_74_0_IVL340R_1876\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l340r_adt_net_117228_\);
    
    REGl252r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_153_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl252r\);
    
    \I2.REG_1l33r_1127\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n1_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL33R_389);
    
    \I2.N_4251_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4251\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4251_Rd1__net_1\);
    
    \I5.COMMANDl2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_14_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl2r_net_1\);
    
    \I2.DT_SRAM_i_1_m2l2r\ : MUX2L
      port map(A => \I2.N_4191\, B => \I2.PIPE2_DTl2r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => \I2.N_4193\);
    
    \I2.TDCDASl18r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl18r, Q => 
        \I2.TDCDASl18r_net_1\);
    
    \I2.CRC32_12_i_m2l12r\ : MUX2H
      port map(A => \I2.DT_SRAMl12r_net_1\, B => 
        \I2.DT_TEMPl12r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854432__net_1\, Y => 
        \I2.N_3957_i_i\);
    
    \I2.CRC32_801\ : MUX2L
      port map(A => \I2.CRC32l6r_net_1\, B => \I2.N_3923\, S => 
        \I2.N_2826_1_ADT_NET_794__332\, Y => \I2.CRC32_801_net_1\);
    
    \I3.REG2_142\ : MUX2L
      port map(A => VDB_inl1r, B => \I3.REG2l1r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG2_142_net_1\);
    
    \I2.EVNT_REJ_2_SQMUXA_1058\ : AND2FT
      port map(A => \I2.FIFO_FULL_net_1\, B => \I3.N_203\, Y => 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26947_\);
    
    \I2.FID_7_0_IVL30R_976\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl78r, C => 
        \I2.FID_7l30r_adt_net_18551_\, Y => 
        \I2.FID_7l30r_adt_net_18559_\);
    
    \I2.TOKENA_CNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TOKENA_CNT_4l1r_net_1\, CLR
         => \I2.un6_clear_stat_i\, Q => \I2.TOKENA_CNTl1r_net_1\);
    
    \I1.NWRLUTI_0_SQMUXA_1_I_0_2070\ : OAI21TTF
      port map(A => \I1.sstatel0r_net_1\, B => \I1.N_380\, C => 
        \PULSE_0l0r_adt_net_834380_Rd1__net_1\, Y => 
        \I1.N_1192_adt_net_133761_\);
    
    \I5.SBYTEl5r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_70_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl5r_net_1\);
    
    \I4.un1_lead_flag_1_5_0\ : MUX2L
      port map(A => LEAD_FLAGl7r, B => LEAD_FLAGl3r, S => 
        \I4.bcnt_i_0_il2r_net_1\, Y => \I4.N_5\);
    
    VAD_padl5r : IOB33PH
      port map(PAD => VAD(5), A => \I3.VADml5r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl5r);
    
    RAMAD_padl13r : OB33PH
      port map(PAD => RAMAD(13), A => RAMAD_cl13r);
    
    \I2.REG_1_c6_i\ : AND2FT
      port map(A => \I2.N_126\, B => 
        \I2.N_3836_i_0_adt_net_2390__net_1\, Y => \I2.N_3835_i_0\);
    
    \I2.OFFSET_37_11l0r\ : MUX2L
      port map(A => \REGl373r\, B => \REGl309r\, S => 
        \I2.PIPE7_DTL27R_86\, Y => \I2.N_715\);
    
    \I2.PIPE1_DTl19r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_746_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl19r_net_1\);
    
    \I2.DTO_16_1_IV_0_0L25R_1086\ : AND2
      port map(A => \I2.N_4671_adt_net_854592__net_1\, B => 
        \I2.DT_TEMPl25r_net_1\, Y => 
        \I2.DTO_16_1l25r_adt_net_29612_\);
    
    \I1.PAGECNTL9R_2851\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854856__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL9R_245\);
    
    \I2.BNC_IDl7r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_38_0\, CLR => 
        \I2.N_4626_i_0\, SET => \I2.N_4609_i_0\, Q => 
        \I2.BNC_IDl7r_net_1\);
    
    DPR_padl24r : IB33
      port map(PAD => DPR(24), Y => DPR_cl24r);
    
    \I2.NWPIPE7\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE6_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE7_net_1\);
    
    \I3.VDBI_57_0_IVL30R_2142\ : AO21
      port map(A => \I3.VDBil30r_net_1\, B => 
        \I3.N_1910_0_adt_net_854340__net_1\, C => 
        \I3.VDBi_57l30r_adt_net_138033_\, Y => 
        \I3.VDBi_57l30r_adt_net_138039_\);
    
    \I3.REGMAPl8r_1633\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un37_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL8R_740\);
    
    \I2.DTESl30r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl30r, Q => 
        \I2.DTES_i_0_il30r\);
    
    \I3.VDBm_0l1r\ : MUX2L
      port map(A => \I3.PIPEAl1r_net_1\, B => \I3.PIPEBl1r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_143\);
    
    \I2.PIPE1_DT_42_1_IVL1R_1518\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855224__net_1\, B => 
        \I2.MIC_ERR_REGSl1r_net_1\, C => \I2.N_12169_i\, Y => 
        \I2.PIPE1_DT_42l1r_adt_net_52045_\);
    
    \I4.FLUSH_3\ : OAI21TTF
      port map(A => \I4.FLUSH_0_sqmuxa_net_1\, B => 
        \I4.STATE1_nsl2r_adt_net_15265_\, C => 
        \I4.FLUSH_3_adt_net_15593_\, Y => \I4.FLUSH_3_net_1\);
    
    \I1.REG_74_0_ivl328r\ : AO21
      port map(A => \REGl328r\, B => \I1.N_201\, C => 
        \I1.REG_74l328r_adt_net_118260_\, Y => \I1.REG_74l328r\);
    
    \I1.REG_1_219\ : MUX2H
      port map(A => \REGl318r\, B => \I1.REG_74l318r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_219_net_1\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3\ : AO21FTT
      port map(A => \I3.REG1l3r_net_1\, B => 
        \I2.DTE_0_sqmuxa_i_o2tt_N_8_Rd1__net_1\, C => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_adt_net_19883_Rd1__net_1\, 
        Y => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\);
    
    \I2.DT_SRAM_0l28r\ : MUX2L
      port map(A => \I2.PIPE10_DTl28r_net_1\, B => 
        \I2.PIPE5_DTl28r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, Y => 
        \I2.N_896\);
    
    \I2.PHASE_865_1727\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_C_834);
    
    \I3.VDBOFFA_31_IV_0L7R_2502\ : AO21
      port map(A => \REGl180r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        C => \I3.VDBoffa_31l7r_adt_net_163276_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163311_\);
    
    \I5.SENS_ADDRl0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SENS_ADDR_6l0r_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.SENS_ADDRl0r_net_1\);
    
    \I2.BNC_IDl0r_1133\ : DFFB
      port map(CLK => CLK_c, D => \I2.BNC_ID_i_0l0r\, CLR => 
        \I2.N_4621_i_0\, SET => \I2.N_4605_i_0\, Q => 
        \I2.BNC_IDL0R_395\);
    
    \I3.WRITES_0\ : DFFC
      port map(CLK => CLK_c, D => \I3.WRITES_23_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.WRITES_net_1\);
    
    \I3.VDBi_10_i_m2l5r\ : AO21
      port map(A => REG_i_il5r, B => \I3.N_283_adt_net_143533_\, 
        C => \I3.N_283_adt_net_143528_\, Y => \I3.N_283\);
    
    \I2.PIPE5_DT_6l9r\ : MUX2L
      port map(A => \I2.PIPE4_DTl9r_net_1\, B => \I2.N_1078\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\, Y
         => \I2.PIPE5_DT_6l9r_net_1\);
    
    \I1.REG_4_sqmuxa_0_a2_0_0_a4\ : OR2
      port map(A => \I1.PAGECNT_318_net_1\, B => \I1.N_299_Ra1_\, 
        Y => \I1.N_268_Ra1_\);
    
    \I1.REG_74_0_IVL315R_1901\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l315r_adt_net_119475_\);
    
    REGl359r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_260_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl359r\);
    
    \I2.ROFFSET_c3\ : NAND2
      port map(A => \I2.ROFFSETL3R_617\, B => 
        \I2.ROFFSET_c2_net_1\, Y => \I2.ROFFSET_c3_net_1\);
    
    \I3.un1_STATE2_15_1_adt_net_3723_\ : OAI21FTF
      port map(A => \I3.STATE2l1r_net_1\, B => \I3.N_297\, C => 
        \I3.un1_STATE2_15_1_adt_net_147708__net_1\, Y => 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\);
    
    DPR_padl30r : IB33
      port map(PAD => DPR(30), Y => DPR_cl30r);
    
    \I3.VDBOFFB_30_IV_0L6R_2373\ : AO21
      port map(A => \REGl403r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l6r_adt_net_161934_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161978_\);
    
    \I1.PAGECNTe_adt_net_854896_\ : BFR
      port map(A => \I1.PAGECNTe\, Y => 
        \I1.PAGECNTe_adt_net_854896__net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2607\ : AO21
      port map(A => \REGl198r\, B => \I3.REGMAPl22r_net_1\, C => 
        \I3.VDBoffa_31l1r_adt_net_164404_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164448_\);
    
    \I2.PIPE4_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl6r_net_1\);
    
    \I2.N_4547_1_adt_net_1209__adt_net_855612_\ : BFR
      port map(A => \I2.N_4547_1_adt_net_1209__net_1\, Y => 
        \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I154_Y_0\ : XOR2FT
      port map(A => \I2.N_3562_i\, B => \I2.N_3560_i_net_1\, Y
         => \I2.ADD_18x18_fast_I154_Y_0\);
    
    \I2.DTO_16_1_IV_1L30R_1069\ : OAI21FTF
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.DTO_9_ivl30r_net_1\, C => 
        \I2.DTO_16_1_iv_1l30r_adt_net_28466_\, Y => 
        \I2.DTO_16_1_iv_1l30r_adt_net_28472_\);
    
    \I5.SCL_1_i_o2_0\ : NOR2
      port map(A => \I5.sstate1l5r_net_1\, B => 
        \I5.sstate1l8r_net_1\, Y => \I5.N_81_i_0_i\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I179_Y\ : XOR2
      port map(A => \I2.N525\, B => \I2.ADD_21x21_fast_I179_Y_0\, 
        Y => \I2.un27_pipe5_dt0l9r\);
    
    \I2.PIPE4_DT_I_IL1R_3084\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DT_I_IL1R_848\);
    
    \I2.TDCDASl1r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl1r, Q => 
        \I2.TDCDASl1r_net_1\);
    
    \I2.STATE1l1r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1l0r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1l1r_net_1\);
    
    \I2.END_TDC3\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_TDC2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_TDC3_net_1\);
    
    \I1.sstate_ns_0_iv_0_0l2r\ : OR2FT
      port map(A => \I1.N_656\, B => 
        \I1.sstate_nsl2r_adt_net_107620_\, Y => \I1.sstate_nsl2r\);
    
    \I2.PIPE9_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_287_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl18r_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2398\ : AO21
      port map(A => \REGl394r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l5r_adt_net_162168_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162175_\);
    
    \I2.PIPE10_DT_17_I_A3_2L13R_1609\ : OR2
      port map(A => \I2.SUB9_i_0_il19r\, B => \I2.SUB9l18r_net_1\, 
        Y => \I2.N_3822_adt_net_64761_\);
    
    \I3.VDBoffbl7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_59_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl7r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL3R_1503\ : AND2FT
      port map(A => \I2.N_3279_0_adt_net_855232__net_1\, B => 
        \I2.MIC_ERR_REGSl3r_net_1\, Y => 
        \I2.PIPE1_DT_42l3r_adt_net_51627_\);
    
    \I3.REG_1_264\ : MUX2H
      port map(A => REGl83r, B => \I3.N_1629\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_264_0\);
    
    \I1.ISI_0_sqmuxa_1_0_i\ : OR3FTT
      port map(A => \I1.N_653\, B => \I1.N_1375_adt_net_134063_\, 
        C => \I1.N_1375_adt_net_134070_\, Y => \I1.N_1375\);
    
    \I2.un7_bnc_id_1_I_16\ : AND2
      port map(A => \I2.N_45\, B => \I2.BNC_IDL2R_711\, Y => 
        \I2.DWACT_FINC_El0r\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I138_Y_0_O2_1_1550\ : AND2
      port map(A => \I2.RAMDT4L5R_817\, B => 
        \I2.PIPE4_DTL11R_410\, Y => \I2.N_75_adt_net_54671_\);
    
    \I2.DTOSl12r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl12r, Q => 
        \I2.DTOSl12r_net_1\);
    
    \I5.sstate1se_0_0_0\ : AO21FTT
      port map(A => TICKl0r, B => \I5.sstate1l12r_net_1\, C => 
        \I5.sstate1_ns_el1r_adt_net_9243_\, Y => 
        \I5.sstate1_ns_el1r\);
    
    \I2.OFFSET_37_26l3r\ : MUX2L
      port map(A => \REGl224r\, B => \I2.N_830\, S => 
        \I2.PIPE7_DTl26r_net_1\, Y => \I2.N_838\);
    
    \I2.SUB9_1_ADD_18x18_fast_I156_Y_0\ : XOR2FT
      port map(A => \I2.SUB8l20r_net_1\, B => \I2.SUB8l19r_net_1\, 
        Y => \I2.ADD_18x18_fast_I156_Y_0\);
    
    \I2.UN1_STATE1_31_I_1592\ : OAI21TTF
      port map(A => \I2.N_3889\, B => 
        \I2.N_3887_adt_net_855068__net_1\, C => 
        \I2.N_3866_adt_net_61361_\, Y => 
        \I2.N_3866_adt_net_61369_\);
    
    \I2.PIPE10_DT_620\ : MUX2L
      port map(A => \I2.PIPE10_DTl15r_net_1\, B => \I2.N_3801\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_620_net_1\);
    
    \I2.N_3283_adt_net_855064_\ : BFR
      port map(A => \I2.N_3283\, Y => 
        \I2.N_3283_adt_net_855064__net_1\);
    
    \I2.SUB9l19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_587_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9_i_0_il19r\);
    
    \I2.OFFSET_37_6l4r\ : MUX2L
      port map(A => \I2.N_671\, B => \I2.N_663\, S => 
        \I2.PIPE7_DTL26R_353\, Y => \I2.N_679\);
    
    \I2.STATE2_NS_I_0_O2_0_0_M7_I_1002\ : MUX2L
      port map(A => \I2.END_EVNT5_839\, B => 
        \I2.END_EVNT10_net_1\, S => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\, Y => 
        \I2.N_4273_adt_net_20831_\);
    
    \I2.PIPE8_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_528_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl0r_net_1\);
    
    FID_padl5r : OB33PH
      port map(PAD => FID(5), A => FID_cl5r);
    
    \I1.REG_74_0_iv_0l394r\ : OAI21FTF
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, C => 
        \I1.REG_74l394r_adt_net_110698_\, Y => \I1.REG_74l394r\);
    
    \I1.REG_74_0_ivl312r\ : AO21
      port map(A => \REGl312r\, B => \I1.N_185\, C => 
        \I1.REG_74l312r_adt_net_119733_\, Y => \I1.REG_74l312r\);
    
    \I3.VDBm_0l30r\ : MUX2L
      port map(A => \I3.PIPEAl30r_net_1\, B => 
        \I3.PIPEBl30r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_172\);
    
    \I3.REG3_131\ : MUX2L
      port map(A => VDB_inl6r, B => \I3.REG3l6r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG3_131_net_1\);
    
    \I2.DTE_cl_63_870\ : MUX2L
      port map(A => \I2.DTE_cl_32l31r\, B => \I2.N_2822\, S => 
        \I2.un1_DTO_cl_1_sqmuxa_2\, Y => \I2.DTE_cl_63_870_net_1\);
    
    \I1.REG_74_0_IVL184R_2050\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l184r_adt_net_131957_\);
    
    \I2.PIPE1_DT_42_1_IVL15R_1432\ : AND2FT
      port map(A => \I2.N_3238\, B => \I2.BNCID_VECTror_net_1\, Y
         => \I2.PIPE1_DT_42l15r_adt_net_48714_\);
    
    REGl305r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_206_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl305r\);
    
    \I5.TEMPDATA_78\ : MUX2L
      port map(A => \I5.TEMPDATAl4r_net_1\, B => REGl129r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_78_net_1\);
    
    \I1.REG_1_216\ : MUX2H
      port map(A => \REGl315r\, B => \I1.REG_74l315r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_216_net_1\);
    
    \I2.RAMDT4L12R_2814\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_142\);
    
    \I1.REG_74l180r_889\ : OR3
      port map(A => \I1.N_41_8\, B => 
        \I1.N_113_ADT_NET_3714__271\, C => \I1.REG_1_sqmuxa\, Y
         => \I1.N_49_267\);
    
    \I2.un1_tdc_res_39_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl415r, Y => 
        \I2.N_4620_i_0\);
    
    \I1.SBYTE_8_0_a2_il4r\ : AND2
      port map(A => \I1.N_371_i\, B => \I1.N_1386\, Y => 
        \I1.N_192\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I186_Y\ : XOR2
      port map(A => \I2.N_82\, B => \I2.ADD_21x21_fast_I186_Y_0\, 
        Y => \I2.un27_pipe5_dt0l16r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I150_Y\ : XOR2FT
      port map(A => \I2.N454_i\, B => 
        \I2.ADD_18x18_fast_I150_Y_0\, Y => \I2.SUB9_1l13r\);
    
    \I2.L2TYPE_4_i_o2_0l14r\ : NAND2
      port map(A => \I2.L2ARRl3r_net_1\, B => \I2.L2ARRl2r_net_1\, 
        Y => \I2.N_4455\);
    
    \I3.PIPEAl10r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_241_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl10r_net_1\);
    
    \I1.N_300_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_300_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_300_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L3R_2578\ : AO21
      port map(A => \REGl184r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.VDBoffa_31l3r_adt_net_164068_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164075_\);
    
    \I2.OFFSET_37_9l7r\ : MUX2L
      port map(A => \REGl396r\, B => \REGl332r\, S => 
        \I2.PIPE7_DTL27R_75\, Y => \I2.N_706\);
    
    \I4.LSRAM_FL_RD_4\ : MUX2L
      port map(A => \I4.LSRAM_FL_RADDR_0_sqmuxa\, B => 
        LSRAM_FL_RD, S => \I4.STATE1l1r_net_1\, Y => 
        \I4.LSRAM_FL_RD_4_net_1\);
    
    \I3.VDBi_57_0_iv_0_a2_1l8r\ : NOR2
      port map(A => \I3.N_354_0\, B => \I3.REGMAPL55R_782\, Y => 
        \I3.N_2037\);
    
    DPR_padl11r : IB33
      port map(PAD => DPR(11), Y => DPR_cl11r);
    
    \I3.TCNT_n2_0_0\ : OR2
      port map(A => \I3.un1_STATE1_10_i_0\, B => 
        \I3.TCNT_n2_adt_net_137234_\, Y => \I3.TCNT_n2\);
    
    \I2.DTO_16_1_IV_0L9R_1173\ : AND2
      port map(A => \I2.N_4671_adt_net_854600__net_1\, B => 
        \I2.DT_TEMPl9r_net_1\, Y => 
        \I2.DTO_16_1l9r_adt_net_33240_\);
    
    \I1.REG_74_8_0_o4_a0_1l324r\ : NAND2
      port map(A => \I1.PAGECNTL9R_835\, B => \I1.PAGECNTL8R_456\, 
        Y => \I1.REG_74_12_220_m9_i_a6_0\);
    
    \I2.STATE1l12r_1538\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl6r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1L12R_645\);
    
    \I2.SUB8_515\ : MUX2H
      port map(A => \I2.SUB8l12r_adt_net_855576__net_1\, B => 
        \I2.SUB8_2l12r\, S => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855144__net_1\, Y => 
        \I2.SUB8_515_net_1\);
    
    \I2.PIPE10_DT_636\ : MUX2L
      port map(A => \I2.PIPE10_DTl31r_net_1\, B => 
        \I2.PIPE9_DTl31r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_636_net_1\);
    
    \I2.RAMDT4L12R_3069\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_823\);
    
    \I2.un7_bnc_id_1_I_31\ : XOR2
      port map(A => \I2.BNC_IDl6r_net_1\, B => \I2.N_29_0\, Y => 
        \I2.I_31_0\);
    
    \I1.REG_74_0_iv_0_0l256r\ : AO21
      port map(A => \REGl256r\, B => \I1.N_658\, C => 
        \I1.REG_74l256r_adt_net_125142_\, Y => \I1.REG_74l256r\);
    
    \I3.RAMAD_VMEl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_28_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl4r);
    
    \I3.PIPEB_99_2324\ : NOR2FT
      port map(A => \I3.PIPEBl20r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_99_adt_net_159873_\);
    
    \I2.MIC_ERR_REGSl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_339_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl10r_net_1\);
    
    \I2.STATE4_ns_i_0l1r\ : AND2
      port map(A => \I2.STATE4l2r_net_1\, B => \I2.N_3376_1\, Y
         => \I2.STATE4_ns_i_0l1r_net_1\);
    
    \I2.DTE_cl_0_sqmuxa_2_adt_net_20049_\ : AND2FT
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__148\, B => 
        \I2.NWPIPE2_578\, Y => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20049__net_1\);
    
    \I2.RAMAD_4_0l7r\ : MUX2H
      port map(A => \I2.RAMAD1l7r_net_1\, B => RAMAD_VMEl7r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_534\);
    
    \I2.DTO_16_1_IV_0L17R_1131\ : AND2
      port map(A => \I2.DTO_1l17r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l17r_adt_net_31522_\);
    
    \I2.STATE5l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE5_nsl2r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.STATE5l1r_net_1\);
    
    \I3.VDBI_57_0_IV_0L9R_2217\ : AO21
      port map(A => \I3.PIPEAl9r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l9r_adt_net_142322_\, Y => 
        \I3.VDBi_57l9r_adt_net_142331_\);
    
    \I1.REG_74_0_ivl395r\ : AO21
      port map(A => \REGl395r\, B => \I1.N_265\, C => 
        \I1.REG_74l395r_adt_net_110612_\, Y => \I1.REG_74l395r\);
    
    \I3.VDBOFFB_30_IV_0L2R_2439\ : AND2
      port map(A => \REGl319r\, B => \I3.REGMAPl37r_net_1\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162698_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I178_Y_2732\ : OR2
      port map(A => \I2.N296_0\, B => \I2.N479_adt_net_538261_\, 
        Y => \I2.N479_adt_net_649015_\);
    
    \I2.END_TDC1_1_SQMUXA_I_O2_1014\ : NOR2
      port map(A => \I2.un6_tdcgdb1_1_net_1\, B => 
        \I2.un6_tdcgdb1_0_net_1\, Y => \I2.N_3887_adt_net_21862_\);
    
    DPR_padl26r : IB33
      port map(PAD => DPR(26), Y => DPR_cl26r);
    
    \I3.un1_REGMAP_30_adt_net_855008_\ : BFR
      port map(A => \I3.un1_REGMAP_30\, Y => 
        \I3.un1_REGMAP_30_adt_net_855008__net_1\);
    
    \I2.CRC32_824\ : MUX2L
      port map(A => \I2.CRC32l29r_net_1\, B => \I2.N_3946\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_824_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0_a2_0_0\ : AO21
      port map(A => \I2.PIPE4_DTL10R_850\, B => 
        \I2.PIPE4_DTL9R_845\, C => \I2.RAMDT4L12R_145\, Y => 
        \I2.ADD_21x21_fast_I140_Y_0_a2_0_0_0\);
    
    \I2.PIPE7_DTL27R_2773\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_66\);
    
    \I2.PIPE5_DT_685\ : MUX2L
      port map(A => \I2.PIPE5_DTl9r_net_1\, B => 
        \I2.PIPE5_DT_6l9r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_685_net_1\);
    
    N_1_I3_TCNT3_c1 : AND2
      port map(A => \I3.TCNT3_i_0_il0r_net_1\, B => 
        \I3.TCNT3l1r_net_1\, Y => \I3.TCNT3_c1\);
    
    \I2.STATE1_ns_0l5r_adt_net_855816_\ : BFR
      port map(A => \I2.STATE1_ns_0l5r\, Y => 
        \I2.STATE1_ns_0l5r_adt_net_855816__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I178_Y\ : NOR3FFT
      port map(A => \I2.N297_0\, B => \I2.N301_2\, C => \I2.N348\, 
        Y => \I2.N479_adt_net_538167_\);
    
    \I3.VDBI_57_IV_0_0L7R_2228\ : NOR2FT
      port map(A => \I1.FBOUTl7r_net_1\, B => \I3.N_2047\, Y => 
        \I3.VDBi_57l7r_adt_net_143099_\);
    
    \I3.ASBS\ : DFFS
      port map(CLK => CLK_c, D => \I3.ASBSF1_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.ASBS_net_1\);
    
    \I3.VDBOFFB_30_IV_0L0R_2476\ : AND2
      port map(A => \REGl373r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163082_\);
    
    \I2.DT_SRAMl16r\ : MUX2L
      port map(A => \I2.N_884\, B => \I2.PIPE2_DTl16r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.DT_SRAMl16r_net_1\);
    
    \I3.REGMAPl26r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un111_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl26r_net_1\);
    
    \I2.L2SERVl3r_1253\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_515\);
    
    \I1.PAGECNT_318_adt_net_854852_\ : BFR
      port map(A => \I1.PAGECNT_318_net_1\, Y => 
        \I1.PAGECNT_318_adt_net_854852__net_1\);
    
    \I2.INT_ERRBF1_495_1705\ : AND2
      port map(A => \I2.N_3876_adt_net_855256__net_1\, B => 
        \I2.INT_ERRBF1_net_1\, Y => 
        \I2.INT_ERRBF1_495_adt_net_90378_\);
    
    \I3.VDBOFFB_30_IV_0L7R_2359\ : AO21
      port map(A => \REGl332r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l7r_adt_net_161760_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161792_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2713\ : 
        NOR3FFT
      port map(A => \I2.N_152_i_0_adt_net_502544_\, B => 
        \I2.N_2358_tz_tz_adt_net_854952__net_1\, C => 
        \I2.N_74_adt_net_55281_\, Y => 
        \I2.N_152_i_0_adt_net_610537_\);
    
    \I2.PIPE1_DT_42_1_IVL0R_1522\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl32r_net_1\, C => 
        \I2.PIPE1_DT_42l0r_adt_net_52231_\, Y => 
        \I2.PIPE1_DT_42l0r_adt_net_52246_\);
    
    \I1.REG_74_8_0_o4_a0_0l324r_722\ : OR2
      port map(A => \I1.PAGECNTL5R_311\, B => 
        \I1.PAGECNTl6r_adt_net_854932__net_1\, Y => 
        \I1.REG_74_1_A0_0L228R_100\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I57_Y_1758\ : NAND2
      port map(A => \I2.N267_0_869\, B => \I2.N264_0_867\, Y => 
        \I2.N307_2_865\);
    
    \I2.OFFSET_37_27l4r\ : MUX2L
      port map(A => \I2.N_839\, B => \I2.N_823\, S => 
        \I2.PIPE7_DTL25R_687\, Y => \I2.N_847\);
    
    \I2.SUB8l15r_adt_net_855572_\ : BFR
      port map(A => \I2.SUB8l15r_net_1\, Y => 
        \I2.SUB8l15r_adt_net_855572__net_1\);
    
    TDCDB_padl14r : IB33
      port map(PAD => TDCDB(14), Y => TDCDB_cl14r);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854236_\ : BFR
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854248__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854236__net_1\);
    
    \I2.MIC_ERR_REGSl44r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_373_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl44r_net_1\);
    
    \I2.DTE_21_1_IV_0L19R_1265\ : AND2
      port map(A => \I2.DTE_1l19r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1l19r_adt_net_37715_\);
    
    \I2.FCNTE_I_1053\ : NOR3FTT
      port map(A => FLUSH, B => \I2.FCNT_c1\, C => 
        \I2.FCNTL2R_600\, Y => \I2.N_3267_adt_net_25763_\);
    
    \I3.PIPEB_101\ : AO21
      port map(A => DPR_cl22r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\, 
        C => \I3.PIPEB_101_adt_net_159789_\, Y => 
        \I3.PIPEB_101_net_1\);
    
    \I2.STATE2_ns_0_a2l4r\ : NAND2
      port map(A => NOESRAME_C_834, B => 
        \I2.STATE2l1r_adt_net_855132__net_1\, Y => \I2.N_4293\);
    
    \I2.N477_adt_net_302175_\ : AND3
      port map(A => \I2.N510\, B => \I2.N498_1_adt_net_88035_\, C
         => \I2.N477_adt_net_301898__net_1\, Y => 
        \I2.N477_adt_net_302175__net_1\);
    
    \I1.REG_13_sqmuxa_adt_net_855440_\ : BFR
      port map(A => \I1.REG_13_sqmuxa\, Y => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\);
    
    \I1.REG_1_205\ : MUX2H
      port map(A => \REGl304r\, B => \I1.REG_74l304r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_205_net_1\);
    
    \I2.L2SERVl0r_1501\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_922_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL12R_608\);
    
    \I2.PIPE1_DT_42_1_IVL14R_1436\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl30r_net_1\, Y => 
        \I2.PIPE1_DT_42l14r_adt_net_48944_\);
    
    \I2.END_EVNT10\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT9_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT10_net_1\);
    
    \I2.PIPE2_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl24r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl24r_net_1\);
    
    \I2.PIPE10_DT_17_il18r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l5r_net_1\, C => \I2.PIPE10_DT_17_i_0l18r_net_1\, 
        Y => \I2.N_3804\);
    
    \I2.CRC32_811\ : MUX2L
      port map(A => \I2.CRC32l16r_net_1\, B => \I2.N_3933\, S => 
        \I2.N_2826_1_ADT_NET_794__331\, Y => \I2.CRC32_811_net_1\);
    
    \I2.resyn_0_I2_BITCNT_n5_i_x2\ : XOR2FT
      port map(A => \I2.N_4330\, B => \I2.BITCNTl5r_net_1\, Y => 
        \I2.N_28_i_0\);
    
    \I3.REGMAPl11r_1636\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un47_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL11R_743\);
    
    \I1.REG_16_sqmuxa_0_a2_m3_e\ : NAND3FFT
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536__net_1\, 
        B => \I1.N_253_96\, C => \I1.REG_74_1_i_a2_a0_2l404r\, Y
         => \I1.REG_16_sqmuxa\);
    
    \I2.RESYN_0_I2_UN1_TRGCNT14_I_940\ : NOR3FTT
      port map(A => \I2.N_3760_adt_net_15913_\, B => 
        \I2.TRGCNT_i_0_il1r\, C => \I2.TRGCNTl4r_net_1\, Y => 
        \I2.N_3760_adt_net_15916_\);
    
    \I3.ADACKCYC_1620\ : DFFC
      port map(CLK => CLK_c, D => \I3.ADACKCYC_112_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => \I3.ADACKCYC_727\);
    
    TDCDA_padl5r : IB33
      port map(PAD => TDCDA(5), Y => TDCDA_cl5r);
    
    \I3.VDBOFFA_31_IV_0L3R_2580\ : OR3
      port map(A => \I3.VDBoffa_31l3r_adt_net_164075_\, B => 
        \I3.VDBoffa_31l3r_adt_net_164069_\, C => 
        \I3.VDBoffa_31l3r_adt_net_164070_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164079_\);
    
    \I2.CHAIN_RDY_490\ : MUX2H
      port map(A => \I2.N_3510\, B => \I2.CHAIN_RDY_net_1\, S => 
        \I2.N_3494\, Y => \I2.CHAIN_RDY_490_net_1\);
    
    \I1.REG_1_218\ : MUX2H
      port map(A => \REGl317r\, B => \I1.REG_74l317r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_218_net_1\);
    
    REGl290r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_191_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl290r\);
    
    \I3.REG_1_177\ : MUX2L
      port map(A => VDB_inl28r, B => REGl76r, S => 
        \I3.N_1935_adt_net_855316__net_1\, Y => \I3.REG_1_177_0\);
    
    \I3.VASl5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_67_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl5r_net_1\);
    
    \I3.REG2_145\ : MUX2L
      port map(A => VDB_inl4r, B => \I3.REG2l4r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG2_145_net_1\);
    
    \I2.MIC_ERR_REGSl33r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_362_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl33r_net_1\);
    
    \I2.OFFSET_37_21l0r\ : MUX2L
      port map(A => \I2.N_787\, B => \I2.N_763\, S => 
        \I2.PIPE7_DTL25R_686\, Y => \I2.N_795\);
    
    \I5.sstate2se_1_0\ : MUX2L
      port map(A => \I5.sstate2l2r_net_1\, B => \I5.N_463\, S => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\, Y => 
        \I5.sstate2_ns_el2r\);
    
    \I3.PIPEA_254\ : MUX2L
      port map(A => \I3.PIPEAl23r_net_1\, B => 
        \I3.PIPEA_8l23r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854660__net_1\, Y
         => \I3.PIPEA_254_net_1\);
    
    \I2.SRAM_EVNTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SRAM_EVNT_n2_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.SRAM_EVNTl2r_net_1\);
    
    \I3.VDBoff_4_i_il2r\ : MUX2L
      port map(A => \I3.VDBoffbl2r_net_1\, B => 
        \I3.VDBoffal2r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_2066\);
    
    \I3.PIPEB_103_2320\ : NOR2FT
      port map(A => \I3.PIPEBl24r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_103_adt_net_159705_\);
    
    \I2.STATE2l1r_adt_net_855128_\ : BFR
      port map(A => \I2.STATE2l1r_adt_net_855132__net_1\, Y => 
        \I2.STATE2l1r_adt_net_855128__net_1\);
    
    \I2.REG_1l41r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n9_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl41r);
    
    REGl203r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_104_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl203r\);
    
    \I3.VDBi_55l1r\ : MUX2H
      port map(A => \I3.VDBil1r_net_1\, B => \I3.RAMDTSl1r_net_1\, 
        S => \I3.N_57_i_0_0_adt_net_854688__net_1\, Y => 
        \I3.VDBi_55l1r_net_1\);
    
    \I1.REG_74_0_ivl321r\ : AO21
      port map(A => \REGl321r\, B => \I1.N_193\, C => 
        \I1.REG_74l321r_adt_net_118959_\, Y => \I1.REG_74l321r\);
    
    \I2.PIPE1_DT_30l12r\ : MUX2L
      port map(A => \I2.TDCDBSl12r_net_1\, B => 
        \I2.TDCDBSl10r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, Y
         => \I2.PIPE1_DT_30l12r_net_1\);
    
    \I2.CRC32_12_0_0_m2l22r\ : MUX2H
      port map(A => \I2.DT_SRAMl22r_net_1\, B => 
        \I2.DT_TEMPl22r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854428__net_1\, Y => 
        \I2.N_4268_i_i\);
    
    NOE32R_pad : OB33PH
      port map(PAD => NOE32R, A => NOE32R_c);
    
    \I4.END_FLUSH_2_933\ : AND2
      port map(A => \I4.STATE1l1r_net_1\, B => END_FLUSH_560, Y
         => \I4.END_FLUSH_2_adt_net_15635_\);
    
    \I2.N_3560_i\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_520_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_3560_i_net_1\);
    
    \I0.BNC_RESF1\ : DFFC
      port map(CLK => CLK_c, D => BNC_RESIN_c, CLR => 
        \I0.un4_hwresi_i\, Q => \I0.BNC_RESF1_net_1\);
    
    \I2.TDCDASl29r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl29r, Q => 
        \I2.TDCDASl29r_net_1\);
    
    \I2.PIPE6_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_465_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl11r_net_1\);
    
    \I3.VDBi_57_0_ivl17r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l17r_net_1\, C
         => \I3.VDBi_57l17r_adt_net_139631_\, Y => 
        \I3.VDBi_57l17r\);
    
    \I2.PIPE9_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_276_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl7r_net_1\);
    
    \I2.DTO_16_1_IV_0L7R_1189\ : AO21
      port map(A => \I2.DTO_1l7r\, B => \I2.N_196\, C => 
        \I2.DTO_16_1l7r_adt_net_33720_\, Y => 
        \I2.DTO_16_1l7r_adt_net_33736_\);
    
    \I3.REG_1_183\ : MUX2L
      port map(A => VDB_inl2r, B => \I3.REGl135r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, Y => 
        \I3.REG_1_183_0\);
    
    \I2.ROFFSET_n9_tz\ : XOR2FT
      port map(A => \I2.ROFFSETl9r_net_1\, B => 
        \I2.ROFFSET_c8_net_1\, Y => \I2.ROFFSET_n9_tz_i\);
    
    \I1.REG_74_10l356r\ : NAND3FFT
      port map(A => \I1.N_1370_278\, B => 
        \I1.N_41_9_adt_net_3739__net_1\, C => \I1.N_273_9_274\, Y
         => \I1.N_41_9\);
    
    VDB_padl13r : IOB33PH
      port map(PAD => VDB(13), A => \I3.VDBml13r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl13r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I178_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_800\, B => 
        \I2.PIPE4_DTl8r_adt_net_854556__adt_net_855024__net_1\, Y
         => \I2.ADD_21x21_fast_I178_Y_0_0\);
    
    \I2.EVNT_NUMl9r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_954_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl9r_net_1\);
    
    \I3.PIPEA1_307\ : MUX2L
      port map(A => \I3.PIPEA1l9r_net_1\, B => 
        \I3.PIPEA1_12l9r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__254\, Y => 
        \I3.PIPEA1_307_net_1\);
    
    \I1.sstatel4r_1156\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl6r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL4R_418\);
    
    \I0.BNC_RESF3\ : DFFC
      port map(CLK => CLK_c, D => BNC_RES_E, CLR => 
        \I0.un4_hwresi_i\, Q => \I0.BNC_RESF3_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2617\ : OR3
      port map(A => \I3.VDBoffa_31l1r_adt_net_164457_\, B => 
        \I3.VDBoffa_31l1r_adt_net_164453_\, C => 
        \I3.VDBoffa_31l1r_adt_net_164454_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164460_\);
    
    ADE_padl8r : OB33PH
      port map(PAD => ADE(8), A => ADE_cl8r);
    
    \I2.SUB9_1_ADD_18x18_fast_I19_Y\ : OA21FTT
      port map(A => \I2.SUB8l20r_net_1\, B => \I2.SUB8l19r_net_1\, 
        C => \I2.N271\, Y => \I2.N284\);
    
    \I1.PAGECNTL6R_2853\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_321_adt_net_854880__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL6R_247\);
    
    FID_padl17r : OB33PH
      port map(PAD => FID(17), A => FID_cl17r);
    
    \I2.DTE_1_867\ : MUX2L
      port map(A => \I2.DTE_1l29r_net_1\, B => \I2.DTE_21_1l29r\, 
        S => \I2.N_2868_1\, Y => \I2.DTE_1_867_net_1\);
    
    \I4.resyn_0_I4_LSRAM_FL_RADDR_9\ : MUX2L
      port map(A => \I4.bcntl0r_net_1\, B => \LSRAM_FL_RADDRl0r\, 
        S => \I4.LSRAM_FL_RADDR_0_sqmuxa_1\, Y => 
        \I4.LSRAM_FL_RADDR_9\);
    
    \I3.VDBOFFA_31_IV_0L7R_2497\ : AND2
      port map(A => \REGl276r\, B => \I3.REGMAPl31r_net_1\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163284_\);
    
    \I0.EV_RESi_1\ : AND2FT
      port map(A => \I0.EV_RESF2_net_1\, B => \I0.EV_RESF1_net_1\, 
        Y => \I0.EV_RESi_1_net_1\);
    
    AMB_padl4r : IB33
      port map(PAD => AMB(4), Y => AMB_cl4r);
    
    \I3.PIPEB_96\ : AO21
      port map(A => DPR_cl17r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\, 
        C => \I3.PIPEB_96_adt_net_159999_\, Y => 
        \I3.PIPEB_96_net_1\);
    
    \I3.VDBOFFB_30_IV_0L2R_2451\ : AO21
      port map(A => \REGl303r\, B => \I3.REGMAPl35r_net_1\, C => 
        \I3.VDBoffb_30l2r_adt_net_162718_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162744_\);
    
    \I2.PIPE1_DT_42_1_IVL17R_1405\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040__net_1\, 
        B => \I2.PIPE1_DT_12l17r_net_1\, Y => 
        \I2.PIPE1_DT_42l17r_adt_net_47635_\);
    
    \I3.RAMDTSl8r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl8r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl8r_net_1\);
    
    \I2.ADO_3l1r\ : MUX2L
      port map(A => \I2.WOFFSETl2r_adt_net_854984__net_1\, B => 
        \I2.ROFFSETl2r_net_1\, S => NOESRAME_c, Y => 
        \I2.ADO_3l1r_net_1\);
    
    \I2.TRGSERVL1R_2952\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l1r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVL1R_469\);
    
    \I1.REG_74_0_iv_0_0_o2_245_m6_i_0_tz_i_adt_net_1555_\ : OR3
      port map(A => \I1.PAGECNTl5r_adt_net_855548__net_1\, B => 
        \I1.PAGECNTl7r_net_1\, C => \I1.PAGECNTl9r_net_1\, Y => 
        \I1.REG_74_0_iv_0_0_o2_245_m6_i_0_tz_i_adt_net_1555__net_1\);
    
    \I2.DTE_21_1_IV_0L6R_1324\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.DTE_2_1l6r_net_1\, C
         => \I2.DTE_21_1l6r_adt_net_38971_\, Y => 
        \I2.DTE_21_1l6r_adt_net_38982_\);
    
    \I3.VDBi_57l7r_adt_net_142961_\ : AO21FTT
      port map(A => \I2.N_4431\, B => \I3.N_2040\, C => 
        \I3.VDBi_57l7r_adt_net_142952__net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_142961__net_1\);
    
    \I2.PIPE7_DTL26R_2903\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_357\);
    
    \I2.CRC32_12_i_0l30r\ : NOR2
      port map(A => \I2.N_2867_1_adt_net_854964__net_1\, B => 
        \I2.N_245_i_i_0\, Y => \I2.N_3947\);
    
    \I1.REG_24_sqmuxa_adt_net_854776_\ : BFR
      port map(A => \I1.REG_24_sqmuxa\, Y => 
        \I1.REG_24_sqmuxa_adt_net_854776__net_1\);
    
    \I2.MIC_ERR_REGSl48r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_377_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl48r_net_1\);
    
    \I2.ADE_4l0r\ : MUX2H
      port map(A => \I2.WOFFSETl1r_adt_net_854992__net_1\, B => 
        \I2.ROFFSETl1r_net_1\, S => NOESRAME_c, Y => 
        \I2.ADE_4l0r_net_1\);
    
    \I3.PIPEBl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_83_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl4r_net_1\);
    
    \I3.un21_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.un60_reg_ads_3\, B => \I3.N_573\, Y => 
        \I3.un21_reg_ads_0_a2_0_a3_net_1\);
    
    \I3.RAMDTSl5r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl5r_net_1\);
    
    \I3.VDBI_57_0_IVL22R_2161\ : AND2
      port map(A => \I3.PIPEAl22r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l22r_adt_net_139083_\);
    
    \I2.PIPE2_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl31r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl31r_net_1\);
    
    \I2.TDCDASl17r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl17r, Q => 
        \I2.TDCDASl17r_net_1\);
    
    \I1.REG_74_0_ivl306r\ : AO21
      port map(A => \REGl306r\, B => \I1.N_177\, C => 
        \I1.REG_74l306r_adt_net_120352_\, Y => \I1.REG_74l306r\);
    
    \I3.VASl6r_1641\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_68_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASL6R_748\);
    
    \I1.REG_1_269\ : MUX2H
      port map(A => \REGl368r\, B => \I1.REG_74l368r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_269_net_1\);
    
    \I2.FID_7_0_ivl14r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl14r_net_1\, 
        C => \I2.FID_7l14r_adt_net_17995_\, Y => \I2.FID_7l14r\);
    
    \I2.resyn_0_I2_FID_436\ : MUX2H
      port map(A => FID_cl20r, B => \I2.FID_7l20r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\, 
        Y => \I2.FID_436\);
    
    \I2.RAMAD1_670\ : MUX2L
      port map(A => \I2.RAMAD1_12l16r_net_1\, B => 
        \I2.RAMAD1l16r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__170\, Y => 
        \I2.RAMAD1_670_net_1\);
    
    \I1.REG_74_2L340R_1875\ : NOR2FT
      port map(A => \I1.REG_74_12_300_N_15\, B => 
        \I1.REG_74_2_2_il340r\, Y => \I1.N_73_10_adt_net_117095_\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2388\ : AND2
      port map(A => \REGl362r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        Y => \I3.VDBoffb_30l5r_adt_net_162140_\);
    
    \I2.INT_ERRAS\ : DFFC
      port map(CLK => CLK_c, D => \I2.INT_ERRAS_526_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.INT_ERRAS_net_1\);
    
    \I1.REG_74_0_iv_0_0_o2_245_m6_i\ : AND2FT
      port map(A => \I1.N_1169_adt_net_854820__net_1\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0_adt_net_125522_\, Y => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\);
    
    \I2.DTE_21_1l26r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l26r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l26r_Rd1__net_1\);
    
    \I2.MIC_REG1_1_sqmuxa_0_adt_net_855860_\ : BFR
      port map(A => \I2.MIC_REG1_1_sqmuxa_0\, Y => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855860__net_1\);
    
    \I3.PIPEBl21r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_100_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl21r_net_1\);
    
    \I2.PIPE10_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_629_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl24r_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I153_Y_I_A4_0_1573\ : OR3
      port map(A => \I2.N_152_i_adt_net_4109__net_1\, B => 
        \I2.N_163_adt_net_1241__net_1\, C => \I2.N307\, Y => 
        \I2.N_86_i_adt_net_57123_\);
    
    \I2.STATEe_illegal\ : OR2
      port map(A => \I2.N_3457_ip_adt_net_23080_\, B => 
        \I2.N_3457_ip_adt_net_23081_\, Y => \I2.N_3457_ip\);
    
    \I2.BNCID_VECT_TILE_I_7_1416\ : NOR3
      port map(A => \I2.I_6_3_i_0_i\, B => \I2.N_11\, C => 
        \I2.I_6_0_i_0_i\, Y => \I2.N_13_adt_net_47925_\);
    
    \I2.PIPE4_DTl12r_1250_1751\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL12R_858\);
    
    RAMAD_padl14r : OB33PH
      port map(PAD => RAMAD(14), A => RAMAD_cl14r);
    
    \I5.AIR_WDATA_61\ : MUX2L
      port map(A => \I5.AIR_WDATAl11r_net_1\, B => 
        \I5.AIR_WDATA_9l11r_net_1\, S => \I5.N_461\, Y => 
        \I5.AIR_WDATA_61_net_1\);
    
    \I3.STATE1_ILLEGAL_2128\ : AO21
      port map(A => \I3.STATE1_ipl6r\, B => \I3.N_1168\, C => 
        \I3.N_1193_ip_adt_net_136550_\, Y => 
        \I3.N_1193_ip_adt_net_136551_\);
    
    \I2.STATE2l2r_1482\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl3r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L2R_589\);
    
    \I2.FIDl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_423_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl7r);
    
    \I2.UN1_END_CHAINA1_0_SQMUXA_I_A2_1_1016\ : AND2
      port map(A => \I2.N_3883_adt_net_854632__net_1\, B => 
        \I2.un1_STATE1_24\, Y => \I2.N_3347_1_adt_net_21905_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I205_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl9r\, B => 
        \I2.PIPE7_DTl9r_net_1\, Y => \I2.SUB_21x21_fast_I205_Y_0\);
    
    \I2.N_2867_1_adt_net_854960_\ : BFR
      port map(A => \I2.N_2867_1_338\, Y => 
        \I2.N_2867_1_adt_net_854960__net_1\);
    
    \I1.sstatel1r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl9r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel1r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL3R_1507\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, B => 
        \I2.PIPE1_DT_30l3r_net_1\, C => 
        \I2.PIPE1_DT_42l3r_adt_net_51635_\, Y => 
        \I2.PIPE1_DT_42l3r_adt_net_51637_\);
    
    \I1.REG_74_0_ivl243r\ : AO21
      port map(A => \REGl243r\, B => \I1.N_113\, C => 
        \I1.REG_74l243r_adt_net_126469_\, Y => \I1.REG_74l243r\);
    
    \I2.DTE_0_sqmuxa_i_o2tt_m2\ : XOR2
      port map(A => \I3.REG2_144_net_1\, B => \I3.REG3_128_net_1\, 
        Y => \I2.DTE_0_sqmuxa_i_o2tt_N_8_Ra1_\);
    
    \I1.N_113_adt_net_126301_\ : AND3FFT
      port map(A => \I1.N_1169_adt_net_854824__net_1\, B => 
        \I1.REG_74_12_220_m9_i_a6_0\, C => 
        \I1.REG_74_8_0_o4_372_N_9_i\, Y => 
        \I1.N_113_adt_net_126301__net_1\);
    
    \I3.REG_44_IL90R_2301\ : MUX2H
      port map(A => VDB_inl7r, B => REGl90r, S => \I3.N_98_0\, Y
         => \I3.N_1636_adt_net_150083_\);
    
    \I3.STATE2l0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE2_nsl4r\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.STATE2l0r_net_1\);
    
    RAMDT_padl0r : IOB33PH
      port map(PAD => RAMDT(0), A => \I1.RAMDT_SPI_1l0r_net_1\, 
        EN => \I1.RAMDT_SPI_E_0\, Y => RAMDT_inl0r);
    
    \I2.DTE_21_1_IVL11R_1294\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855128__net_1\, B => 
        \I2.EVNT_WORDl7r_net_1\, Y => 
        \I2.DTE_21_1l11r_adt_net_38399_\);
    
    \I3.VDBoff_4_i_il6r\ : MUX2L
      port map(A => \I3.VDBoffbl6r_net_1\, B => 
        \I3.VDBoffal6r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_79\);
    
    \I1.REG_74_0_ivl393r\ : AO21
      port map(A => \REGl393r\, B => \I1.N_265\, C => 
        \I1.REG_74l393r_adt_net_110784_\, Y => \I1.REG_74l393r\);
    
    \I2.CRC32_803\ : MUX2L
      port map(A => \I2.CRC32l8r_net_1\, B => \I2.N_3925\, S => 
        \I2.N_2826_1_ADT_NET_794__332\, Y => \I2.CRC32_803_net_1\);
    
    \I2.DTE_1l20r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l20r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l20r_Rd1__net_1\);
    
    \I1.BYTECNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_314_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTl0r_net_1\);
    
    \I2.FID_7_0_ivl12r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl12r_net_1\, 
        C => \I2.FID_7l12r_adt_net_18183_\, Y => \I2.FID_7l12r\);
    
    REGl385r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_286_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl385r\);
    
    \I2.OFFSET_37_18l7r\ : MUX2L
      port map(A => \REGl252r\, B => \REGl188r\, S => 
        \I2.PIPE7_DTL27R_75\, Y => \I2.N_778\);
    
    \I1.REG_74_0_IVL373R_1826\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l373r_adt_net_113087_\);
    
    \I2.DTE_21_1_IV_0L26R_1242\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.G_EVNT_NUMl10r_net_1\, 
        C => \I2.DTE_21_1l26r_adt_net_36962_\, Y => 
        \I2.DTE_21_1l26r_adt_net_36963_\);
    
    \I2.MIC_ERR_REGSl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_354_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl25r_net_1\);
    
    \I5.AIR_CHAIN_15\ : XOR2
      port map(A => \I5.AIR_CHAIN_net_1\, B => 
        \I5.sstate2_5_sqmuxa\, Y => \I5.AIR_CHAIN_15_net_1\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_adt_net_19883_Rd1_\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_adt_net_19883_Ra1_\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_adt_net_19883_Rd1__net_1\);
    
    \I1.REG_1_266\ : MUX2H
      port map(A => \REGl365r\, B => \I1.REG_74l365r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_266_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I5_P0N_i_a4_733\ : OR2
      port map(A => \I2.RAMDT4L12R_143\, B => 
        \I2.PIPE4_DTl5r_adt_net_854416__net_1\, Y => 
        \I2.N_89_0_111\);
    
    \I3.REG2_1_sqmuxa_i_0\ : AO21TTF
      port map(A => \I3.REGMAPl50r_net_1\, B => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        C => HWCLEAR, Y => \I3.N_1563\);
    
    \I3.PIPEA1_319\ : MUX2L
      port map(A => \I3.PIPEA1l21r_net_1\, B => 
        \I3.PIPEA1_12l21r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__251\, Y => 
        \I3.PIPEA1_319_net_1\);
    
    \I2.PIPE6_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_466_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl12r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I120_Y_0_78_tz_tz\ : AO21
      port map(A => \I2.N_52\, B => \I2.N357\, C => 
        \I2.N_2360_tz_tz_adt_net_54584_\, Y => \I2.N_2360_tz_tz\);
    
    \I2.L2ARR_943\ : MUX2L
      port map(A => \I2.L2ARRl1r_net_1\, B => \I2.L2ARR_n1_net_1\, 
        S => \I2.N_4482_0\, Y => \I2.L2ARR_943_net_1\);
    
    \I2.PIPE2_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl9r_net_1\);
    
    \I0.BNC_RESF2\ : DFFC
      port map(CLK => CLK_c, D => \I0.BNC_RESF1_net_1\, CLR => 
        \I0.un4_hwresi_i\, Q => \I0.BNC_RESF2_net_1\);
    
    \I5.REG_1l442r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_25_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl442r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I141_Y_0_o4\ : AOI21
      port map(A => \I2.N_107_0_adt_net_320361_\, B => 
        \I2.N525_0_adt_net_318530_\, C => 
        \I2.N_107_0_adt_net_320362_\, Y => 
        \I2.N522_0_adt_net_329169_\);
    
    REGl354r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_255_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl354r\);
    
    \I2.STATEE_ILLEGAL_1028\ : AO21
      port map(A => \I2.N_3496_adt_net_926__net_1\, B => 
        \I2.STATEel4r_net_1\, C => \I2.N_3457_ip_adt_net_23071_\, 
        Y => \I2.N_3457_ip_adt_net_23079_\);
    
    \I2.DTESl19r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl19r, Q => 
        \I2.DTESl19r_net_1\);
    
    \I1.BITCNTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BITCNT_315_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BITCNTl2r_net_1\);
    
    \I5.SBYTE_9_il1r\ : MUX2L
      port map(A => \I5.COMMANDl9r_net_1\, B => 
        \I5.SBYTEl0r_net_1\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.N_16\);
    
    \I2.FIDl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_445\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl29r);
    
    \I3.VASl7r_1640\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_69_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VAS_I_0_IL7R_747\);
    
    \I3.PIPEA_8l14r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854476__net_1\, B => 
        \I3.N_223\, Y => \I3.PIPEA_8l14r_net_1\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854512_\ : BFR
      port map(A => \I3.N_243_4_adt_net_1290__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854512__net_1\);
    
    RAMAD_padl17r : OB33PH
      port map(PAD => RAMAD(17), A => RAMAD_cl17r);
    
    \I2.LSRAM_OUTl14r_adt_net_854944_\ : BFR
      port map(A => \I2.LSRAM_OUTl14r\, Y => 
        \I2.LSRAM_OUTl14r_adt_net_854944__net_1\);
    
    \I2.BNCID_VECTROR_1424\ : OA21
      port map(A => \I2.BNCID_VECTror_9_tz_adt_net_48098_\, B => 
        \I2.BNCID_VECTror_9_tz_adt_net_48099_\, C => 
        \I2.TRGSERVL2R_581\, Y => 
        \I2.BNCID_VECTror_adt_net_48367_\);
    
    \I3.REGMAPl44r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un201_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl44r_net_1\);
    
    \I2.PIPE5_DT_6_0l0r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l0r\, B => 
        \I2.un27_pipe5_dt0l0r\, S => 
        \I2.dataout_0_adt_net_855800__net_1\, Y => \I2.N_1069\);
    
    VDB_padl19r : IOB33PH
      port map(PAD => VDB(19), A => \I3.VDBml19r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl19r);
    
    \I2.EVNT_WORD_722\ : MUX2H
      port map(A => \I2.EVNT_WORDl9r_net_1\, B => \I2.I_52\, S
         => \I2.N_2864_0_adt_net_854272__net_1\, Y => 
        \I2.EVNT_WORD_722_net_1\);
    
    \I0.CLEAR_935\ : NAND2FT
      port map(A => \HWRES_3_ADT_NET_738__17\, B => HWCLEAR, Y
         => \I0.CLEAR_adt_net_15816_\);
    
    \I2.DTO_16_1_IVL10R_1171\ : AO21
      port map(A => \I2.N_457\, B => \I2.DTE_2_1l10r_net_1\, C
         => \I2.DTO_16_1l10r_adt_net_33056_\, Y => 
        \I2.DTO_16_1l10r_adt_net_33065_\);
    
    \I2.REG_1_C10_I_1739\ : AND2
      port map(A => REG_i_0_il42r, B => \I2.N_3853\, Y => 
        \I2.N_3839_i_0_adt_net_101262_\);
    
    \I2.DTOSl10r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl10r, Q => 
        \I2.DTOSl10r_net_1\);
    
    \I2.TRGARR_3_I_1\ : AND2
      port map(A => TDCTRG_c, B => \I2.TRGARRl0r_net_1\, Y => 
        \I2.DWACT_ADD_CI_0_TMPl0r\);
    
    \I2.PIPE6_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_458_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl4r_net_1\);
    
    \I3.REGMAP_I_0_A2L52R_2094\ : AND3FFT
      port map(A => \I3.N_2018\, B => \I3.N_1907_264\, C => 
        \I3.N_638_adt_net_134642_\, Y => 
        \I3.N_638_adt_net_134645_\);
    
    \I2.PIPE4_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl14r_net_1\);
    
    \I1.REG_16_sqmuxa_0_a2_m3_e_717\ : NAND3FFT
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__net_1\, 
        B => \I1.N_253_98\, C => \I1.REG_74_1_i_a2_a0_2l404r\, Y
         => \I1.REG_16_SQMUXA_95\);
    
    \I2.OFFSET_37_5l1r\ : MUX2L
      port map(A => \REGl398r\, B => \REGl334r\, S => 
        \I2.PIPE7_DTL27R_84\, Y => \I2.N_668\);
    
    \I1.REG_1_255\ : MUX2H
      port map(A => \REGl354r\, B => \I1.REG_74l354r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_255_net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__2843\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__201\);
    
    \I2.MIC_ERR_REGSl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_345_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl16r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2550\ : AND2
      port map(A => \REGl249r\, B => \I3.REGMAPl28r_net_1\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163850_\);
    
    \I0.un12_clear\ : OR2
      port map(A => COM_SER_c, B => \I0.CLEAR_net_1\, Y => 
        \I0.un12_clear_i\);
    
    \I3.VDBoff_118\ : MUX2L
      port map(A => \I3.VDBoffl2r_net_1\, B => \I3.N_2066\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_118_net_1\);
    
    \I2.PIPE10_DT_17_i_0l19r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855592__net_1\, B => 
        \I2.PIPE9_DTl19r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l19r_net_1\);
    
    \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m3\ : MUX2H
      port map(A => \I2.MIC_REG2L3R_ADT_NET_834020_RD1__215\, B
         => \I2.MIC_REG3L3R_484\, S => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Rd1__net_1\, Y => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m3_net_1\);
    
    \I2.LSRAM_INl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_408_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl24r_net_1\);
    
    \I2.DTE_2_1_0l8r\ : XOR2
      port map(A => \I2.CRC32l16r_net_1\, B => 
        \I2.CRC32l4r_net_1\, Y => \I2.DTE_2_1_0l8r_net_1\);
    
    \I1.N_65_ADT_NET_1433__2848\ : OR3
      port map(A => \I1.N_65_12_273\, B => 
        \I1.N_193_adt_net_118653__net_1\, C => \I1.N_97_6\, Y => 
        \I1.N_65_ADT_NET_1433__218\);
    
    \I3.SINGCYC_956\ : DFFC
      port map(CLK => CLK_c, D => \I3.SINGCYC_115_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.SINGCYC_334\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I210_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl14r_adt_net_854944__net_1\, B
         => \I2.PIPE7_DTl14r_net_1\, Y => 
        \I2.SUB_21x21_fast_I210_Y_0\);
    
    \I2.END_CHAINB1\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.END_CHAINB1_709_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.END_CHAINB1_net_1\);
    
    \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834768_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_0_sqmuxa_i_0_N_3_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834768_Rd1__net_1\);
    
    \I3.VDBil27r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_367_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil27r_net_1\);
    
    \I2.FIDl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_437\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl21r);
    
    \I2.un1_tdc_res_33_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl407r, Y => 
        \I2.N_4614_i_0\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I216_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl20r\, B => 
        \I2.PIPE7_DTl20r_net_1\, Y => 
        \I2.SUB_21x21_fast_I216_Y_0\);
    
    \I2.REG_1_c4_i_a2_0\ : NOR3
      port map(A => REGL35R_564, B => REGL36R_565, C => 
        \I2.N_122\, Y => \I2.N_124\);
    
    \I2.PIPE7_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl4r_net_1\);
    
    \I3.VDBoffa_31_iv_i_a2_il6r\ : AND2
      port map(A => \REGl179r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        Y => \I3.N_2070_adt_net_163454_\);
    
    \I2.SUB9l13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_581_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9_i_0_il13r\);
    
    RAMDT_padl3r : IOB33PH
      port map(PAD => RAMDT(3), A => \I1.RAMDT_SPI_1l3r_net_1\, 
        EN => \I1.RAMDT_SPI_e_net_1\, Y => RAMDT_inl3r);
    
    \I2.PIPE1_DTl0r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_727_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl0r_net_1\);
    
    \I2.DTO_16_1_iv_0_a2_2l21r_673\ : AND3
      port map(A => \I2.N_223_54\, B => \I2.N_4182\, C => 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_888__net_1\, Y => 
        \I2.N_196_51\);
    
    \I2.un3_tdcgda1_1_adt_net_21664_\ : OR2
      port map(A => \I2.TDCDASl31r_net_1\, B => 
        \I2.TDCDASl29r_net_1\, Y => 
        \I2.un3_tdcgda1_1_adt_net_21664__net_1\);
    
    \I1.REG_74_12_220_m9_i_o6\ : NOR3
      port map(A => \I1.PAGECNTl6r_adt_net_854924__net_1\, B => 
        \I1.PAGECNTl5r_net_1\, C => 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__adt_net_855516__net_1\, 
        Y => \I1.REG_74_12_220_N_13\);
    
    \I5.sstate2_5_sqmuxa_0_a3\ : AND2FT
      port map(A => \I5.SENS_ADDR_1_sqmuxa_1_0_net_1\, B => 
        \I5.sstate2l0r_net_1\, Y => \I5.sstate2_5_sqmuxa\);
    
    \I5.SSTATE1SE_0_0_0_910\ : AND2
      port map(A => TICKL0R_557, B => \I5.COMMANDl1r_net_1\, Y
         => \I5.sstate1_ns_el1r_adt_net_9246_\);
    
    \I3.VDBOFFA_31_IV_0L5R_2542\ : AO21
      port map(A => \REGl194r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.VDBoffa_31l5r_adt_net_163688_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163695_\);
    
    \I3.VDBOFFA_31_IV_0L0R_2619\ : AND2
      port map(A => \REGl237r\, B => \I3.REGMAPl27r_net_1\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164598_\);
    
    \I2.EVNT_WORDl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_719_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl6r_net_1\);
    
    \I2.resyn_0_I2_FID_433\ : MUX2H
      port map(A => FID_cl17r, B => \I2.FID_7l17r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\, 
        Y => \I2.FID_433\);
    
    \I1.REG_1_268\ : MUX2H
      port map(A => \REGl367r\, B => \I1.REG_74l367r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_268_net_1\);
    
    \I3.REG_1_293\ : MUX2L
      port map(A => VDB_inl11r, B => REGl112r, S => 
        \I3.N_318_adt_net_855884__net_1\, Y => \I3.REG_1_293_0\);
    
    \I5.SBYTE_9_il6r\ : MUX2L
      port map(A => \I5.COMMANDl14r_net_1\, B => 
        \I5.SBYTEl5r_net_1\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.N_26\);
    
    \I2.PIPE2_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl22r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl22r_net_1\);
    
    REGl207r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_108_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl207r\);
    
    ADO_padl0r : OB33PH
      port map(PAD => ADO(0), A => ADO_cl0r);
    
    \I2.un1_TOKENA_CNT_I_8\ : XOR2
      port map(A => TICKL0R_557, B => \I2.TOKENA_CNTl0r_net_1\, Y
         => \I2.DWACT_ADD_CI_0_partial_sum_0l0r\);
    
    \I2.ADE_4l5r\ : MUX2H
      port map(A => \I2.WOFFSETl6r\, B => \I2.ROFFSETl6r_net_1\, 
        S => NOESRAME_c, Y => \I2.ADE_4l5r_net_1\);
    
    REGl283r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_184_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl283r\);
    
    \I3.VDBi_16_m_i_m2l11r\ : MUX2H
      port map(A => REGl27r, B => REGl43r, S => 
        \I3.REGMAPl7r_net_1\, Y => \I3.N_278\);
    
    REGl336r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_237_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl336r\);
    
    TDCDB_padl10r : IB33
      port map(PAD => TDCDB(10), Y => TDCDB_cl10r);
    
    \I2.PIPE1_DT_42_1_IVL14R_1438\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl10r\, Y => 
        \I2.PIPE1_DT_42l14r_adt_net_48954_\);
    
    \I2.DT_TEMPl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_768_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl7r_net_1\);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854240_\ : BFR
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854248__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854240__net_1\);
    
    \I5.DATA_12l11r\ : MUX2L
      port map(A => REGl128r, B => \I5.SBYTEl3r_net_1\, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l11r_net_1\);
    
    \I2.DTO_16_1_ivl22r\ : OR2
      port map(A => \I2.DTO_16_1l22r_adt_net_30361_\, B => 
        \I2.DTO_16_1l22r_adt_net_30362_\, Y => \I2.DTO_16_1l22r\);
    
    \I2.MIC_ERR_REGS_370\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl42r_net_1\, B => 
        \I2.MIC_ERR_REGSl41r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_370_net_1\);
    
    \I2.FID_7_0_IVL9R_1715\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl57r, C => 
        \I2.FID_7l9r_adt_net_92645_\, Y => 
        \I2.FID_7l9r_adt_net_92653_\);
    
    \I3.VDBI_57_IVL3R_2257\ : AO21
      port map(A => \I3.PIPEAl3r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l3r_adt_net_145062_\, Y => 
        \I3.VDBi_57l3r_adt_net_145072_\);
    
    \I2.PIPE1_DT_42_1_IVL12R_1453\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\, B => 
        \I2.PIPE1_DT_30l12r_net_1\, C => 
        \I2.PIPE1_DT_42l12r_adt_net_49442_\, Y => 
        \I2.PIPE1_DT_42l12r_adt_net_49458_\);
    
    \I2.N_3558_i_adt_net_855584_\ : BFR
      port map(A => \I2.N_3558_i_net_1\, Y => 
        \I2.N_3558_i_adt_net_855584__net_1\);
    
    \I2.BNC_IDl1r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_5_1\, CLR => 
        \I2.N_4628_i_0\, SET => \I2.N_4614_i_0\, Q => 
        \I2.BNC_IDl1r_net_1\);
    
    VAD_padl12r : IOB33PH
      port map(PAD => VAD(12), A => \I3.VADml12r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl12r);
    
    \I2.SUB9_1_ADD_18X18_FAST_I115_Y_1649\ : AND3
      port map(A => \I2.N469\, B => \I2.N300\, C => \I2.N304\, Y
         => \I2.N457_adt_net_69532_\);
    
    \I3.REG2l1r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG2_142_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l1r_net_1\);
    
    \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__2837\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854852__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__186\);
    
    \I2.un21_sram_empty_NE\ : NOR3FTT
      port map(A => \I2.un21_sram_empty_NE_adt_net_24173_\, B => 
        \I2.un21_sram_empty_1_net_1\, C => 
        \I2.un21_sram_empty_0_net_1\, Y => 
        \I2.un21_sram_empty_NE_net_1\);
    
    ADO_padl3r : OB33PH
      port map(PAD => ADO(3), A => ADO_cl3r);
    
    \I2.L2TYPE_4_il7r\ : OAI21FTF
      port map(A => \I2.L2TYPEl7r_net_1\, B => \I2.N_4466\, C => 
        \I2.N_4445_adt_net_67839_\, Y => \I2.N_4445\);
    
    \I2.DTE_2_1_0l5r\ : XOR2
      port map(A => \I2.CRC32l25r_net_1\, B => 
        \I2.CRC32l13r_net_1\, Y => \I2.DTE_2_1_0l5r_net_1\);
    
    \I0.REG_1l27r\ : DFFC
      port map(CLK => CLK_c, D => \I0.REG_1_3_net_1\, CLR => 
        NPWON_c_i_0, Q => REGl27r);
    
    \I3.VDBI_31L1R_2716\ : MUX2L
      port map(A => \I3.REGl134r\, B => 
        \I3.VDBi_29l1r_adt_net_411517_\, S => 
        \I3.REGMAPl17r_adt_net_854292__net_1\, Y => 
        \I3.VDBi_31l1r_adt_net_614331_\);
    
    \I2.BNCID_VECTrff_8\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_8_257_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_8\);
    
    \I2.PIPE8_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_542_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl14r_net_1\);
    
    \I2.DTO_16_1_iv_0_0l25r\ : OR2
      port map(A => \I2.DTO_16_1l25r_adt_net_29623_\, B => 
        \I2.DTO_16_1l25r_adt_net_29624_\, Y => \I2.DTO_16_1l25r\);
    
    \I2.N_1170_adt_net_1217__adt_net_855704_\ : BFR
      port map(A => \I2.N_1170_adt_net_1217__net_1\, Y => 
        \I2.N_1170_adt_net_1217__adt_net_855704__net_1\);
    
    \I2.TDCDASl26r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl26r, Q => 
        \I2.TDCDASl26r_net_1\);
    
    \I2.DTE_21_1_IV_0L16R_1272\ : AO21
      port map(A => \I2.N_3965_0\, B => 
        \I2.G_EVNT_NUM_i_0_il0r_net_1\, C => 
        \I2.DTE_21_1l16r_adt_net_37825_\, Y => 
        \I2.DTE_21_1l16r_adt_net_37834_\);
    
    \I2.N_3558_i\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_519_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_3558_i_net_1\);
    
    \I5.sstate2l3r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate2_ns_el1r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate2l3r_net_1\);
    
    \I3.REG_1l138r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_186_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl138r\);
    
    \I2.ADO_3l7r\ : MUX2L
      port map(A => \I2.WOFFSETl8r\, B => \I2.ROFFSETl8r_net_1\, 
        S => NOESRAME_C_243, Y => \I2.ADO_3l7r_net_1\);
    
    \I3.VDBoffal6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_50_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal6r_net_1\);
    
    \I3.TCNT4_387\ : MUX2H
      port map(A => \I3.TCNT4l1r_net_1\, B => \I3.TCNT4_n1_net_1\, 
        S => \I3.TICKl2r_net_1\, Y => \I3.TCNT4_387_net_1\);
    
    \I1.REG_74_0_IV_I_A2L207R_2027\ : AND2
      port map(A => \REGl207r\, B => \I1.N_183_i_0\, Y => 
        \I1.N_1346_adt_net_129931_\);
    
    DTO_padl14r : IOB33PH
      port map(PAD => DTO(14), A => \I2.DTO_1l14r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl14r);
    
    \I1.REG_1_97\ : MUX2H
      port map(A => \REGl196r\, B => \I1.REG_74l196r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\, Y
         => \I1.REG_1_97_net_1\);
    
    NOESRAME_pad : OB33PH
      port map(PAD => NOESRAME, A => NOESRAME_c);
    
    \I3.PIPEAl22r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_253_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl22r_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl9r\ : OR3
      port map(A => \I2.PIPE1_DT_42l9r_adt_net_50189_\, B => 
        \I2.PIPE1_DT_42l9r_adt_net_50198_\, C => 
        \I2.PIPE1_DT_42l9r_adt_net_50199_\, Y => 
        \I2.PIPE1_DT_42l9r\);
    
    \I2.CRC32_813\ : MUX2L
      port map(A => \I2.CRC32l18r_net_1\, B => \I2.N_3935\, S => 
        \I2.N_2826_1_ADT_NET_794__330\, Y => \I2.CRC32_813_net_1\);
    
    \I1.REG_74_i_o2_0_0_364_m9_i_a7_0\ : NAND2
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854400__net_1\, 
        B => \I1.PAGECNTl5r_net_1\, Y => 
        \I1.REG_74_1_396_m7_i_a5_0\);
    
    \I2.MIC_REG1_305\ : MUX2L
      port map(A => \I2.MIC_REG1l5r_net_1\, B => 
        \I2.MIC_REG1l4r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG1_305_net_1\);
    
    \I2.OFFSET_37_8l6r\ : MUX2L
      port map(A => \REGl363r\, B => \REGl299r\, S => 
        \I2.PIPE7_DTL27R_68\, Y => \I2.N_697\);
    
    \I3.VDBm_0l16r\ : MUX2L
      port map(A => \I3.PIPEAl16r_net_1\, B => 
        \I3.PIPEBl16r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_158\);
    
    \I2.L2TYPE_4_il8r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855716__net_1\, B => 
        \I2.N_4444_adt_net_67711_\, C => 
        \I2.N_4444_adt_net_67754_\, Y => \I2.N_4444\);
    
    \I1.sstate_ns_i_0_o2l0r\ : NOR3
      port map(A => \I1.SSTATEL9R_433\, B => \I1.SSTATEL7R_754\, 
        C => \I1.SSTATEL8R_524\, Y => \I1.N_355\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_A2_1_2662\ : OR2
      port map(A => \I2.N_107_adt_net_256839_\, B => 
        \I2.N_107_ADT_NET_256840__384\, Y => \I2.N_107\);
    
    \I2.SUB9_1_ADD_18x18_fast_I114_un1_Y\ : AND3
      port map(A => \I2.N313_0\, B => \I2.N466_adt_net_71184_\, C
         => \I2.N333\, Y => \I2.I114_un1_Y\);
    
    \I2.BNCID_VECTror\ : MUX2L
      port map(A => \I2.BNCID_VECTror_adt_net_48326_\, B => 
        \I2.BNCID_VECTror_adt_net_48422_\, S => 
        \I2.TRGSERVl3r_net_1\, Y => \I2.BNCID_VECTror_net_1\);
    
    \I3.un106_reg_ads_0_a2_0_a2_0_990\ : NOR2FT
      port map(A => \I3.VASl12r_net_1\, B => \I3.N_547_372\, Y
         => \I3.N_548_368\);
    
    \I2.N_4547_1_adt_net_1209__adt_net_855620_\ : BFR
      port map(A => \I2.N_4547_1_adt_net_1209__net_1\, Y => 
        \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\);
    
    \I2.EVNT_WORD_720\ : MUX2H
      port map(A => \I2.EVNT_WORDl7r_net_1\, B => \I2.I_38\, S
         => \I2.N_2864_0_adt_net_854272__net_1\, Y => 
        \I2.EVNT_WORD_720_net_1\);
    
    \I2.DTE_21_1_0_IV_1L30R_1230\ : OAI21TTF
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_289\, B => 
        \I2.DT_SRAMl30r_adt_net_854200__net_1\, C => 
        \I2.DTE_21_1_0_iv_1l30r_adt_net_36505_\, Y => 
        \I2.DTE_21_1_0_iv_1l30r_adt_net_36511_\);
    
    \I1.PAGECNT_n5_0_0_x2\ : XOR2
      port map(A => \I1.PAGECNTl5r_adt_net_855548__net_1\, B => 
        \I1.N_310_Rd1__net_1\, Y => \I1.N_398_i_i_0_i\);
    
    \I2.TOKENA_CNT_4l0r\ : AND2
      port map(A => \I2.N_3899\, B => 
        \I2.DWACT_ADD_CI_0_partial_sum_0l0r\, Y => 
        \I2.TOKENA_CNT_4l0r_net_1\);
    
    \I2.OFFSET_37_28l7r\ : MUX2L
      port map(A => \I2.N_850\, B => \I2.N_802\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_858\);
    
    \I3.VDBm_i_m2l7r\ : MUX2L
      port map(A => \I3.PIPEAl7r_net_1\, B => \I3.PIPEBl7r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_129\);
    
    \I1.BYTECNTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_309_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTl5r_net_1\);
    
    \I3.VDBI_57_0_IVL10R_2213\ : AND2
      port map(A => \I3.VDBil10r_net_1\, B => 
        \I3.N_1764_adt_net_854352__net_1\, Y => 
        \I3.VDBi_57l10r_adt_net_141874_\);
    
    \I2.TOKENA_CNT_4l1r\ : AND2
      port map(A => \I2.N_3899\, B => \I2.I_10_0\, Y => 
        \I2.TOKENA_CNT_4l1r_net_1\);
    
    \I3.VDBI_57_0_IVL11R_2209\ : AND2
      port map(A => \I3.VDBil11r_net_1\, B => 
        \I3.N_1764_adt_net_854352__net_1\, Y => 
        \I3.VDBi_57l11r_adt_net_141431_\);
    
    \I2.STATE4l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE4_ns_i_0l1r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE4l1r_net_1\);
    
    \I1.BYTECNT_n5_i_0_o2_1\ : NAND2
      port map(A => \I1.BYTECNTl5r_net_1\, B => \I1.N_334\, Y => 
        \I1.N_335\);
    
    \I2.SUB9l17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_585_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9_i_0_il17r\);
    
    \I2.OFFSET_37_7l1r\ : MUX2L
      port map(A => \I2.N_676\, B => \I2.N_652\, S => 
        \I2.PIPE7_DTL25R_683\, Y => \I2.N_684\);
    
    \I2.DTO_16_1_IV_0L8R_1182\ : AO21
      port map(A => \I2.DTO_1l8r\, B => \I2.N_196\, C => 
        \I2.DTO_16_1l8r_adt_net_33488_\, Y => 
        \I2.DTO_16_1l8r_adt_net_33490_\);
    
    \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872_\ : BFR
      port map(A => \I5.REG_2_sqmuxa_0_adt_net_975__net_1\, Y => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\);
    
    \I2.OFFSET_37_18l5r\ : MUX2L
      port map(A => \REGl250r\, B => \REGl186r\, S => 
        \I2.PIPE7_DTL27R_79\, Y => \I2.N_776\);
    
    \I2.N_4671_adt_net_854592_\ : BFR
      port map(A => \I2.N_4671\, Y => 
        \I2.N_4671_adt_net_854592__net_1\);
    
    \I2.PHASE_864_1726\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_C_833);
    
    REGl376r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_277_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl376r\);
    
    \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276_\ : BFR
      port map(A => \I3.un1_STATE2_7_1_adt_net_1473__net_1\, Y
         => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I136_Y_0_o2_m4_e_i_1\ : 
        AO21
      port map(A => \I2.PIPE4_DTL10R_851\, B => 
        \I2.PIPE4_DTL11R_409\, C => \I2.RAMDT4L12R_825\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_i_1\);
    
    \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004_\ : 
        BFR
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__net_1\, Y => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\);
    
    DTE_padl21r : IOB33PH
      port map(PAD => DTE(21), A => \I2.DTE_1l21r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl21r);
    
    \I3.VDBi_57l7r_adt_net_142960_\ : AND2FT
      port map(A => \I3.N_2018\, B => \I3.N_2056\, Y => 
        \I3.VDBi_57l7r_adt_net_142960__net_1\);
    
    \I3.PIPEA1_12l15r\ : AND2
      port map(A => DPR_cl15r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854500__net_1\, Y => 
        \I3.PIPEA1_12l15r_net_1\);
    
    \I1.PAGECNT_n5_0_0\ : OAI21
      port map(A => \I1.N_398_i_i_0_i\, B => 
        \I1.un1_sbyte13_1_i_1_adt_net_854520__net_1\, C => 
        \I1.N_473_206\, Y => \I1.PAGECNT_n5\);
    
    REGl315r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_216_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl315r\);
    
    \I3.VDBOFFB_30_IV_0L0R_2490\ : OR3
      port map(A => \I3.VDBoffb_30l0r_adt_net_163125_\, B => 
        \I3.VDBoffb_30l0r_adt_net_163119_\, C => 
        \I3.VDBoffb_30l0r_adt_net_163120_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163129_\);
    
    \I1.REG_4_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_268_Rd1__adt_net_854800__net_1\, B => 
        \I1.N_242\, Y => \I1.REG_4_sqmuxa\);
    
    REGl189r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_90_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl189r\);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854664_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854664__net_1\);
    
    \I2.DTE_21_1_IV_2L1R_1341\ : AND2
      port map(A => GA_cl1r, B => 
        \I2.STATE2l1r_adt_net_855120__net_1\, Y => 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39583_\);
    
    \I2.FID_423\ : MUX2H
      port map(A => FID_cl7r, B => \I2.FID_7l7r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        Y => \I2.FID_423_net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2465\ : AO21
      port map(A => \REGl382r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l1r_adt_net_162892_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162930_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I63_Y\ : AND2
      port map(A => \I2.N255_0\, B => \I2.N258_0\, Y => 
        \I2.N313_1\);
    
    \I3.STATE1_tr24_i_0_a3_5\ : OAI21TTF
      port map(A => \I3.N_2083\, B => \I3.REGMAPl13r_net_1\, C
         => \I3.REGMAPl51r_net_1\, Y => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135544_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I119_Y_i_o4\ : OAI21FTF
      port map(A => \I2.N_128_adt_net_54290_\, B => \I2.N_31\, C
         => \I2.N_3_adt_net_59496_\, Y => \I2.N_3\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I138_Y_0_0\ : AO21FTT
      port map(A => \I2.N_74_i_0_i\, B => 
        \I2.ADD_21x21_fast_I138_Y_0_0_adt_net_58475_\, C => 
        \I2.N_75\, Y => \I2.ADD_21x21_fast_I138_Y_0_0\);
    
    \I3.RAMAD_VMEl7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_31_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl7r);
    
    \I2.DTO_16_1_IV_0L13R_1153\ : AND2
      port map(A => \I2.DTO_1l13r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l13r_adt_net_32386_\);
    
    \I3.N_354_0_adt_net_855368_\ : BFR
      port map(A => \I3.N_354_0\, Y => 
        \I3.N_354_0_adt_net_855368__net_1\);
    
    \I2.PIPE1_DT_42_1_IVL7R_1481\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl39r_net_1\, C => 
        \I2.PIPE1_DT_42l7r_adt_net_50673_\, Y => 
        \I2.PIPE1_DT_42l7r_adt_net_50691_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I112_un1_Y\ : NOR3FFT
      port map(A => \I2.N302\, B => \I2.N306\, C => \I2.N329\, Y
         => \I2.I112_un1_Y_adt_net_71518_\);
    
    \I2.BNCID_VECTROR_1426\ : AOI21FTF
      port map(A => \I2.BNCID_VECTror_10_tz_0_net_1\, B => 
        \I2.BNCID_VECTror_10_tz_adt_net_48171_\, C => 
        \I2.TRGSERVL2R_583\, Y => 
        \I2.BNCID_VECTror_adt_net_48461_\);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854244_\ : BFR
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854248__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854244__net_1\);
    
    \I2.DTO_16_1_iv_0_o2_2tt_21_m2\ : XOR2
      port map(A => \I2.MIC_REG2l3r_adt_net_834020_Rd1__net_1\, B
         => \I2.MIC_REG3L3R_804\, Y => 
        \I2.DTO_16_1_iv_0_o2_2tt_21_N_8\);
    
    \I2.DTO_16_1_iv_0_a2_4_18_m7_0_a5_1\ : AND3FTT
      port map(A => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, B => 
        \I2.END_EVNT2_net_1\, C => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        Y => \I2.DTO_16_1_iv_0_a2_4_18_N_14_i\);
    
    \I2.PIPE1_DT_42_1_IVL3R_1505\ : OAI21TTF
      port map(A => GA_cl3r, B => \I2.N_3238\, C => 
        \I2.PIPE1_DT_42l3r_adt_net_51634_\, Y => 
        \I2.PIPE1_DT_42l3r_adt_net_51635_\);
    
    \I2.DTE_1l14r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l14r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l14r_Rd1__net_1\);
    
    \I2.DTE_21_1_IV_0_IL25R_1245\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.G_EVNT_NUMl9r_net_1\, 
        C => \I2.N_4644_adt_net_37064_\, Y => 
        \I2.N_4644_adt_net_37065_\);
    
    \I1.REG_16_sqmuxa_0_a2_0\ : OR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835132_RD1__884\, B
         => \I1.REG_74_1_A0_0L228R_99\, Y => \I1.N_253\);
    
    RAMAD_padl4r : OB33PH
      port map(PAD => RAMAD(4), A => RAMAD_cl4r);
    
    \I5.TEMPDATA_74\ : MUX2L
      port map(A => \I5.TEMPDATAl0r_net_1\, B => REGl125r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_74_net_1\);
    
    \I2.PIPE10_DT_615\ : MUX2L
      port map(A => \I2.PIPE10_DTl10r_net_1\, B => 
        \I2.PIPE9_DTl10r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_615_net_1\);
    
    \I2.UN1_REG80_I_1702\ : NOR3FFT
      port map(A => \I2.N_3824_adt_net_90287_\, B => REGl32r, C
         => REGl44r, Y => \I2.N_3824_adt_net_90294_\);
    
    \I2.DTESl3r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl3r, Q => 
        \I2.DTESl3r_net_1\);
    
    \I2.un28_sram_empty_13_0\ : MUX2L
      port map(A => \I2.N_631\, B => \I2.N_630\, S => 
        \I2.RPAGEL14R_614\, Y => \I2.N_632\);
    
    \I3.VDBOFFB_30_IV_0L3R_2424\ : AND2
      port map(A => \REGl360r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        Y => \I3.VDBoffb_30l3r_adt_net_162520_\);
    
    \I3.VDBi_40_0_i_m2l9r\ : MUX2L
      port map(A => REGl427r, B => REGl443r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_1854\);
    
    \I2.DTE_1l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_841_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l1r_net_1\);
    
    \I2.SUB8_514\ : MUX2H
      port map(A => \I2.SUB8l11r_adt_net_855580__net_1\, B => 
        \I2.SUB8_2l11r\, S => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855144__net_1\, Y => 
        \I2.SUB8_514_net_1\);
    
    \I2.PIPE9_DT_299\ : MUX2H
      port map(A => \I2.PIPE8_DTl30r_net_1\, B => 
        \I2.PIPE9_DTl30r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_299_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL5R_1492\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl1r\, Y => 
        \I2.PIPE1_DT_42l5r_adt_net_51177_\);
    
    \I2.DTO_16_1_iv_0_0l18r\ : OR2
      port map(A => \I2.DTO_16_1l18r_adt_net_31345_\, B => 
        \I2.DTO_16_1l18r_adt_net_31346_\, Y => \I2.DTO_16_1l18r\);
    
    \I3.NRDMEBi_2_sqmuxa_i_0_o3\ : AND2FT
      port map(A => \I3.un15_anycyc_net_1\, B => 
        \I3.N_297_adt_net_147649_\, Y => \I3.N_297\);
    
    \I3.VDBI_57_0_IV_0_0L24R_2155\ : AND2FT
      port map(A => \I3.N_1917_adt_net_855336__net_1\, B => 
        \I3.REGl157r\, Y => \I3.VDBi_57l24r_adt_net_138805_\);
    
    \I3.VDBoffl0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_116_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl0r_net_1\);
    
    \I2.un28_sram_empty_11_0\ : MUX2L
      port map(A => \I2.L2TYPEL11R_662\, B => \I2.L2TYPEL3R_661\, 
        S => \I2.RPAGEL15R_520\, Y => \I2.N_630\);
    
    \I2.PIPE1_DT_42_1_IVL12R_1452\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855228__net_1\, B => 
        \I2.MIC_ERR_REGSl12r_net_1\, C => 
        \I2.PIPE1_DT_42l12r_adt_net_49456_\, Y => 
        \I2.PIPE1_DT_42l12r_adt_net_49457_\);
    
    \I2.REG_1_n2_0\ : XOR2
      port map(A => REGl34r, B => \I2.N_3830\, Y => 
        \I2.REG_1_n2_0_net_1\);
    
    \I2.EVNT_NUM_954\ : MUX2L
      port map(A => \I2.EVNT_NUMl9r_net_1\, B => 
        \I2.EVNT_NUM_n9_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_954_net_1\);
    
    \I3.PULSE_46_0_IV_0_0L6R_2291\ : OAI21FTF
      port map(A => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        B => \I3.N_98_0\, C => \I3.PULSE_46l6r_adt_net_147009_\, 
        Y => \I3.PULSE_46l6r_adt_net_147015_\);
    
    \I3.REG_1l50r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_151_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl50r);
    
    \I2.ADEl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l5r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl5r);
    
    \I2.SRAM_EVNT_c3_i\ : OAI21FTF
      port map(A => \I2.N_3860\, B => \I2.N_128_1\, C => 
        \I2.N_3828_adt_net_101749_\, Y => \I2.N_3828\);
    
    \I2.DTE_21_1l19r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l19r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l19r_Rd1__net_1\);
    
    \I1.SBYTE_8_0_IL3R_1752\ : OA21TTF
      port map(A => \FBOUTl2r\, B => \I1.N_603_i\, C => 
        \I1.N_337\, Y => \I1.N_202_adt_net_105770_\);
    
    REGl294r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_195_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl294r\);
    
    \I2.RAMDT4L3R_3011\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl3r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L3R_765\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854492_\ : BFR
      port map(A => \I3.N_243_4_adt_net_1290__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854492__net_1\);
    
    \I3.VDBi_57_0_iv_0_a2_3l13r\ : OR2
      port map(A => \I3.REGMAPl17r_adt_net_854296__net_1\, B => 
        \I3.N_2014_121\, Y => \I3.N_2015\);
    
    \I3.VDBi_57_iv_0_0_a2_11l7r_938\ : AND2FT
      port map(A => \I3.N_2017_317\, B => 
        \I3.REGMAPl9r_adt_net_854328__net_1\, Y => 
        \I3.N_2044_316\);
    
    \I2.BNCID_VECTra14_1\ : AND2FT
      port map(A => \I2.TRGSERVL0R_466\, B => \I2.TRGSERVL1R_469\, 
        Y => \I2.BNCID_VECTra14_1_net_1\);
    
    \I2.STATE1l7r_1526\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl11r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE1L7R_633\);
    
    \I1.REG_74_8_0_o4_a0_0l324r_724\ : OR2
      port map(A => \I1.PAGECNTL5R_310\, B => \I1.PAGECNTL6R_248\, 
        Y => \I1.REG_74_1_A0_0L228R_102\);
    
    ADE_padl3r : OB33PH
      port map(PAD => ADE(3), A => ADE_cl3r);
    
    \I2.PIPE4_DTl13r_1535\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl13r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL13R_642\);
    
    \I2.DTO_16_1l17r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l17r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l17r_Rd1__net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I137_Y_I_2708\ : AND2FT
      port map(A => \I2.N_20_i_0\, B => 
        \I2.N_40_0_adt_net_58199_\, Y => 
        \I2.N_40_0_adt_net_577293_\);
    
    \I3.VDBI_57_0_IVL17R_2179\ : AND2
      port map(A => \I3.PIPEAl17r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l17r_adt_net_139627_\);
    
    \I2.LSRAM_IN_410\ : MUX2L
      port map(A => \I2.PIPE5_DTl26r_net_1\, B => 
        \I2.LSRAM_INl26r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_410_net_1\);
    
    \I2.DTE_21_1_IV_0L21R_1255\ : AND2
      port map(A => \I2.DT_TEMPl21r_net_1\, B => \I2.N_4038_233\, 
        Y => \I2.DTE_21_1l21r_adt_net_37485_\);
    
    \I2.DTE_21_1_IV_0L21R_1257\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.G_EVNT_NUMl5r_net_1\, 
        C => \I2.DTE_21_1l21r_adt_net_37496_\, Y => 
        \I2.DTE_21_1l21r_adt_net_37497_\);
    
    \I5.SDAOUT_12_IV_0_O4_911\ : NOR2FT
      port map(A => \I5.sstate1l6r_net_1\, B => \I5.N_67\, Y => 
        \I5.N_71_adt_net_9287_\);
    
    MTDCRESA_pad : OB33PH
      port map(PAD => MTDCRESA, A => MTDCRESA_c);
    
    REGl242r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_143_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl242r\);
    
    \I2.SUB8_521\ : MUX2H
      port map(A => \I2.N_3562_i\, B => \I2.SUB8_2l18r\, S => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855140__net_1\, Y => 
        \I2.SUB8_521_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl26r\ : OA21TTF
      port map(A => \I2.PIPE1_DT_42_3_0l28r\, B => 
        \I2.EVNT_NUMl10r_net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_2_il26r\, Y => 
        \I2.PIPE1_DT_42_1_iv_i_0l26r\);
    
    \I2.WOFFSET_13_il5r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_24\, Y => \I2.N_4248\);
    
    \I2.PIPE1_DT_42_1_IVL19R_1398\ : OAI21FTF
      port map(A => REGl439r, B => 
        \I2.N_3234_adt_net_855648__net_1\, C => 
        \I2.PIPE1_DT_42l19r_adt_net_47255_\, Y => 
        \I2.PIPE1_DT_42l19r_adt_net_47261_\);
    
    \I2.DTOSl18r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl18r, Q => 
        \I2.DTOSl18r_net_1\);
    
    \I3.VDBi_40_0_i_m2l4r\ : MUX2L
      port map(A => REGl422r, B => REGl438r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_136\);
    
    \I2.un1_tdc_res_34_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl412r, Y => 
        \I2.N_4615_i_0\);
    
    \I2.majority_reg_i_il6r\ : AO21
      port map(A => \I2.MIC_REG3l6r_net_1\, B => 
        \I2.MIC_REG1_i_il6r_net_1\, C => \REGl28r_adt_net_36082_\, 
        Y => REGl28r);
    
    \I5.AIR_PULSE\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_PULSE_64_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_PULSE_net_1\);
    
    \I3.REG_1_204\ : MUX2L
      port map(A => VDB_inl23r, B => \I3.REGl156r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\, Y => 
        \I3.REG_1_204_0\);
    
    \I3.PIPEA1l1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_299_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l1r_net_1\);
    
    REGl213r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_114_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl213r\);
    
    \I3.REG_1_297\ : MUX2L
      port map(A => VDB_inl15r, B => REGl116r, S => 
        \I3.N_318_adt_net_855884__net_1\, Y => \I3.REG_1_297_0\);
    
    \I2.RAMADl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l9r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl9r);
    
    \I1.sstate_tr17_0_a2_0_a4\ : AND2FT
      port map(A => \I1.N_604\, B => \I1.COMMAND_net_1\, Y => 
        \I1.sstate_nsl4r\);
    
    \I3.PIPEA_8l24r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854460__net_1\, B => 
        \I3.N_233\, Y => \I3.PIPEA_8l24r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I151_Y_i_a2_2\ : OA21
      port map(A => \I2.RAMDT4L5R_820\, B => 
        \I2.PIPE4_DTl19r_net_1\, C => \I2.N519_131\, Y => 
        \I2.N_152_i_adt_net_54886_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I13_P0N_i_a4\ : OR2
      port map(A => \I2.RAMDT4L12R_145\, B => 
        \I2.PIPE4_DTL13R_641\, Y => \I2.N_92_0\);
    
    \I1.sstate_ns_1_iv_0_i_a4_2l8r\ : OAI21FTF
      port map(A => \I1.sstatel9r_net_1\, B => 
        \I1.N_321_adt_net_855540__net_1\, C => 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r_adt_net_107364_\, Y => 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r\);
    
    \I2.DTO_16_1_IV_0_O2_2TT_21_M3_1063\ : NOR2
      port map(A => \I2.MIC_REG2l3r_adt_net_834020_Rd1__net_1\, B
         => \I2.MIC_REG3l3r_net_1\, Y => 
        \I2.DTO_16_1_iv_0_o2_2tt_21_m3_adt_net_27978_\);
    
    \I2.N_2864_0_adt_net_854276_\ : BFR
      port map(A => \I2.N_2864_0\, Y => 
        \I2.N_2864_0_adt_net_854276__net_1\);
    
    \I2.CRC32_12_i_0l6r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_251_i_i_0\, Y => 
        \I2.N_3923\);
    
    \I2.PIPE1_DT_30l1r\ : MUX2H
      port map(A => \I2.TDCDBSl20r_net_1\, B => 
        \I2.TDCDBSl1r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, Y
         => \I2.PIPE1_DT_30l1r_net_1\);
    
    \I1.REG_74_0_IVL316R_1900\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l316r_adt_net_119389_\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855524_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__281\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\);
    
    \I2.OFFSET_37_13l2r\ : MUX2L
      port map(A => \I2.N_725\, B => \I2.N_709\, S => 
        \I2.PIPE7_DTL25R_685\, Y => \I2.N_733\);
    
    \I3.un44_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_634\, B => \I3.N_573\, Y => 
        \I3.un44_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.L2TYPE_4_i_o2_0l10r\ : OR2FT
      port map(A => \I2.L2ARRl3r_net_1\, B => \I2.L2ARRl2r_net_1\, 
        Y => \I2.N_4459\);
    
    REGl186r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_87_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl186r\);
    
    \I2.L2SERVl3r_1256\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_518\);
    
    \I3.REGMAP_i_il46r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un211_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_il46r_net_1\);
    
    \I2.TDCDASl7r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl7r, Q => 
        \I2.TDCDASl7r_net_1\);
    
    \I2.WOFFSETl5r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl5r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl5r_Rd1__net_1\);
    
    \I2.SUB9_579\ : MUX2H
      port map(A => \I2.SUB9_i_0_il11r\, B => \I2.SUB9_1l11r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_579_net_1\);
    
    REGl349r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_250_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl349r\);
    
    \I1.UN1_SBYTE13_2_I_I_A2_I_1775\ : OAI21TTF
      port map(A => \I1.N_321_232\, B => \I1.N_355\, C => 
        \PULSE_0L0R_ADT_NET_834380_RD1__830\, Y => 
        \I1.N_223_adt_net_108706_\);
    
    \I2.DT_TEMP_781\ : MUX2H
      port map(A => \I2.DT_TEMPl20r_net_1\, B => 
        \I2.DT_TEMP_7l20r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_781_net_1\);
    
    \I2.un8_evread_1_adt_net_855792_\ : BFR
      port map(A => \I2.un8_evread_1\, Y => 
        \I2.un8_evread_1_adt_net_855792__net_1\);
    
    \I2.PIPE5_DT_6l5r\ : MUX2L
      port map(A => 
        \I2.PIPE4_DTl5r_adt_net_854412__adt_net_855600__net_1\, B
         => \I2.N_1074\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, Y => 
        \I2.PIPE5_DT_6l5r_net_1\);
    
    \I3.VDBI_57_0_IVL16R_2181\ : AND2
      port map(A => \I3.PIPEAl16r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l16r_adt_net_139761_\);
    
    \I2.MIC_ERR_REGS_346\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl18r_net_1\, B => 
        \I2.MIC_ERR_REGSl17r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_346_net_1\);
    
    \I2.EVNT_NUM_c4\ : AND2
      port map(A => \I2.EVNT_NUML4R_598\, B => 
        \I2.EVNT_NUM_c3_net_1\, Y => \I2.EVNT_NUM_c4_net_1\);
    
    \I2.PIPE10_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_623_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl18r_net_1\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854464_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854472__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854464__net_1\);
    
    REGl287r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_188_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl287r\);
    
    \I2.MIC_ERR_REGS_350\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl22r_net_1\, B => 
        \I2.MIC_ERR_REGSl21r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_350_net_1\);
    
    \I3.VASl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_65_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl3r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I121_Y_i_o2\ : OA21FTT
      port map(A => \I2.N_17_0\, B => 
        \I2.N_2358_tz_tz_adt_net_854956__net_1\, C => 
        \I2.N_29_i_0_adt_net_59529_\, Y => \I2.N_29_i_0\);
    
    \I2.MIC_REG1_303\ : MUX2H
      port map(A => \I2.MIC_REG1l2r_net_1\, B => 
        \I2.MIC_REG1l3r_adt_net_834596_Rd1__net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG1_303_net_1\);
    
    \I3.PULSE_46_0_iv_0_0l8r\ : AO21
      port map(A => PULSEl8r, B => 
        \I3.N_311_adt_net_854748__net_1\, C => 
        \I3.PULSE_46l8r_adt_net_146836_\, Y => \I3.PULSE_46l8r\);
    
    \I3.VDBi_57_0_iv_0_0_a2l13r\ : NAND2FT
      port map(A => \I3.REGMAPL16R_444\, B => \I3.N_354_0_128\, Y
         => \I3.N_2014\);
    
    \I2.OFFSETl0r_1479\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_560_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL0R_586\);
    
    \I3.RAMDTSl12r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl12r_net_1\);
    
    \I2.BNC_IDl4r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_20_0\, CLR => 
        \I2.N_4627_i_0\, SET => \I2.N_4607_i_0\, Q => 
        \I2.BNC_IDl4r_net_1\);
    
    \I3.STATE1_NS_0_IV_0_0_A3_0_1_0L7R_2081\ : NOR2
      port map(A => \I3.REGMAPL27R_533\, B => \I3.REGMAPL26R_532\, 
        Y => \I3.N_58_i_0_adt_net_134395_\);
    
    \I2.OFFSET_37_28l5r\ : MUX2L
      port map(A => \I2.N_848\, B => \I2.N_800\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_856\);
    
    \I2.DTO_9_ivl14r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl14r_net_1\, 
        C => \I2.DTO_9l14r_adt_net_32142_\, Y => \I2.DTO_9l14r\);
    
    \I2.L2TYPE_4_il2r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4450_adt_net_68435_\, C => 
        \I2.N_4450_adt_net_68478_\, Y => \I2.N_4450\);
    
    \I0.CLEAR_STATi\ : DFFC
      port map(CLK => CLK_c, D => \I0.CLEAR_STATi_4_net_1\, CLR
         => \I0.un12_clear_i\, Q => CLEAR_STAT);
    
    DPR_padl6r : IB33
      port map(PAD => DPR(6), Y => DPR_cl6r);
    
    \I2.END_EVNT10_1145_1785\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT9_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT10_891\);
    
    \I2.TDC_651\ : MUX2H
      port map(A => \I2.TDCl1r_net_1\, B => 
        \I2.RAMAD1_12l14r_net_1\, S => 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_1038__net_1\, Y => 
        \I2.TDC_651_net_1\);
    
    \I2.FID_7_0_ivl1r\ : OA21FTF
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl1r_net_1\, 
        C => \I2.FID_7_0_iv_0l1r_net_1\, Y => 
        \I2.FID_7_0_ivl1r_net_1\);
    
    \I2.resyn_0_I2_BITCNT_n4_i_a5\ : NOR2
      port map(A => \I2.N_4329\, B => \I2.BITCNT_i_0_il4r\, Y => 
        \I2.N_4337\);
    
    \I2.RESYN_0_I2_LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_946\ : NOR2
      port map(A => \I2.PIPE4_DTl22r_net_1\, B => \I2.N_2328_tz\, 
        Y => \I2.N_4524_adt_net_16635_\);
    
    \I2.OFFSET_37_9l2r\ : MUX2L
      port map(A => \REGl391r\, B => \REGl327r\, S => 
        \I2.PIPE7_DTL27R_82\, Y => \I2.N_701\);
    
    \I2.L2TYPEl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_594_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_i_0_il5r\);
    
    \I3.RAMAD_VMEl14r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_38_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl14r);
    
    \I2.BNCID_VECTrff_13_252_0\ : AO21
      port map(A => \I2.BNCID_VECTwa13_1_net_1\, B => 
        \I2.BNCID_VECTrff_12_253_0_a2_0\, C => 
        \I2.BNCID_VECTro_13\, Y => 
        \I2.BNCID_VECTrff_13_252_0_net_1\);
    
    \I2.DTE_21_1_iv_0l19r\ : OR3
      port map(A => \I2.DTE_21_1l19r_adt_net_37715_\, B => 
        \I2.DTE_21_1l19r_adt_net_37723_\, C => 
        \I2.DTE_21_1l19r_adt_net_37724_\, Y => \I2.DTE_21_1l19r\);
    
    ADE_padl4r : OB33PH
      port map(PAD => ADE(4), A => ADE_cl4r);
    
    \I2.SUB9_1_ADD_18X18_FAST_I46_Y_1648\ : AND2
      port map(A => \I2.ca_0_and2\, B => \I2.G_1_4\, Y => 
        \I2.N311_adt_net_69399_\);
    
    \I3.REG2l4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG2_145_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l4r_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl7r\ : OR3
      port map(A => \I2.PIPE1_DT_42l7r_adt_net_50683_\, B => 
        \I2.PIPE1_DT_42l7r_adt_net_50692_\, C => 
        \I2.PIPE1_DT_42l7r_adt_net_50693_\, Y => 
        \I2.PIPE1_DT_42l7r\);
    
    FBOUTl2r : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_60_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \FBOUTl2r\);
    
    \I2.DTOSl7r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl7r, Q => 
        \I2.DTOSl7r_net_1\);
    
    TDCDA_padl14r : IB33
      port map(PAD => TDCDA(14), Y => TDCDA_cl14r);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I171_Y\ : XOR2
      port map(A => \I2.N_85\, B => \I2.ADD_21x21_fast_I171_Y_0\, 
        Y => \I2.un27_pipe5_dt0l1r\);
    
    \I2.DTESl6r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl6r, Q => 
        \I2.DTESl6r_net_1\);
    
    \I3.REGMAPl9r_adt_net_854308_\ : BFR
      port map(A => \I3.REGMAPl9r_adt_net_854320__net_1\, Y => 
        \I3.REGMAPl9r_adt_net_854308__net_1\);
    
    TICKl1r : DFFC
      port map(CLK => CLK_c, D => \I3.un10_tcnt2_i_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => \TICKl1r\);
    
    REGl262r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_163_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl262r\);
    
    \I5.SBYTE_9_il4r\ : MUX2L
      port map(A => \I5.COMMANDl12r_net_1\, B => 
        \I5.SBYTEl3r_net_1\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.N_22\);
    
    \I2.BNC_IDl1r_1132\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_5_1\, CLR => 
        \I2.N_4628_i_0\, SET => \I2.N_4614_i_0\, Q => 
        \I2.BNC_IDL1R_394\);
    
    \I1.REG_74_0_IV_0_0_O2_245_M6_I_1973\ : AO21FTF
      port map(A => \I1.REG_74_8_1_tzl340r_net_1\, B => 
        \I1.REG_74_0_iv_0_0_o2_245_m6_i_0_tz_i_adt_net_1555__net_1\, 
        C => \I1.REG_74_1_404_m7_i_a5_0_net_1\, Y => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0_adt_net_125522_\);
    
    \I3.VDBI_57_0_IV_0L9R_2218\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => \I3.N_92\, C
         => \I3.VDBi_57l9r_adt_net_142331_\, Y => 
        \I3.VDBi_57l9r_adt_net_142332_\);
    
    \I1.REG_74_0_ivl354r\ : AO21
      port map(A => \REGl354r\, B => \I1.N_225\, C => 
        \I1.REG_74l354r_adt_net_115773_\, Y => \I1.REG_74l354r\);
    
    \I2.MAJORITY_REG_I_0L2R_897\ : AOI21
      port map(A => \I2.MIC_REG3L2R_462\, B => 
        \I2.MIC_REG1L2R_464\, C => \I2.MIC_REG2L2R_463\, Y => 
        \I2.N_3876_adt_net_4861_\);
    
    \I2.PIPE9_DT_290\ : MUX2L
      port map(A => \I2.PIPE9_DTl21r_net_1\, B => 
        \I2.PIPE8_DTl21r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_290_net_1\);
    
    \I3.PIPEBl24r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_103_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl24r_net_1\);
    
    RAMDT_padl1r : IOB33PH
      port map(PAD => RAMDT(1), A => \I1.RAMDT_SPI_1l1r_net_1\, 
        EN => \I1.RAMDT_SPI_E_0\, Y => RAMDT_inl1r);
    
    \I5.SDAnoe_8_0_o4_0\ : OR2FT
      port map(A => \I5.sstate1l3r_net_1\, B => \I5.N_67\, Y => 
        \I5.N_70\);
    
    \I1.REG_74_0_iv_i_a2l202r\ : AO21
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_1341_adt_net_130361_\, Y => \I1.N_1341\);
    
    \I2.un1_STATE1_12_0_a2_i\ : OR2
      port map(A => \I2.STATE1L12R_645\, B => 
        \I2.STATE1l11r_net_1\, Y => \I2.N_3870\);
    
    \I2.RAMAD_4_0l5r\ : MUX2H
      port map(A => \I2.RAMAD1l5r_net_1\, B => RAMAD_VMEl5r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_532\);
    
    \I1.N_311_I_I_RD1__3008\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_311_i_i_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.N_311_I_I_RD1__762\);
    
    VAD_padl14r : IOB33PH
      port map(PAD => VAD(14), A => \I3.VADml14r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl14r);
    
    \I2.DTO_16_1_IV_0L17R_1133\ : AO21
      port map(A => \I2.N_197_152\, B => \I2.N_188\, C => 
        \I2.DTO_16_1l17r_adt_net_31522_\, Y => 
        \I2.DTO_16_1l17r_adt_net_31532_\);
    
    \I1.REG_6_sqmuxa_adt_net_854708_\ : BFR
      port map(A => \I1.REG_6_sqmuxa\, Y => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\);
    
    \I2.TDCDBSl1r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl1r, Q => 
        \I2.TDCDBSl1r_net_1\);
    
    \I1.REG_74_0_ivl188r\ : AO21
      port map(A => \REGl188r\, B => \I1.N_57_268\, C => 
        \I1.REG_74l188r_adt_net_131613_\, Y => 
        \I1.REG_74l188r_net_1\);
    
    \I1.REG_74_0_IVL263R_1960\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, Y => 
        \I1.REG_74l263r_adt_net_124457_\);
    
    \I2.PIPE1_DTl27r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_754_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl27r_net_1\);
    
    \I2.MIC_ERR_REGSl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_348_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl19r_net_1\);
    
    \I1.REG_1_79\ : MUX2H
      port map(A => \REGl178r\, B => \I1.REG_74l178r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\, Y => 
        \I1.REG_1_79_net_1\);
    
    \I2.PIPE7_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl30r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl30r_net_1\);
    
    \I2.DTO_16_1_iv_0_a2_4_18_m7_0_0\ : AO21TTF
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608__net_1\, 
        B => \I2.DTO_16_1_iv_0_a2_4tt_18_m2_0_a2_net_1\, C => 
        \I2.DT_TEMPl18r_net_1\, Y => 
        \I2.DTO_16_1_iv_0_a2_4_18_m7_0_0_i\);
    
    \I3.PIPEA_8_0l15r\ : MUX2L
      port map(A => DPR_cl15r, B => \I3.PIPEA1l15r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855348__net_1\, Y => \I3.N_224\);
    
    \I2.un7_bnc_id_1_I_5\ : XOR2
      port map(A => \I2.BNC_IDl1r_net_1\, B => 
        \I2.BNC_IDl0r_net_1\, Y => \I2.I_5_1\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855448_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__292\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\);
    
    \I2.DTO_16_1_iv_0l28r\ : AO21FTT
      port map(A => \I2.DTO_1l28r_net_1\, B => \I2.N_196_52\, C
         => \I2.DTO_16_1_iv_0l28r_adt_net_28950_\, Y => 
        \I2.DTO_16_1_iv_0l28r_net_1\);
    
    \I3.N_1910_0_adt_net_854348_\ : BFR
      port map(A => \I3.N_1910_0\, Y => 
        \I3.N_1910_0_adt_net_854348__net_1\);
    
    \I2.SUB8_523\ : AND2
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855160__net_1\, B
         => \I2.SUB_21x21_fast_I216_Y_0\, Y => 
        \I2.SUB8_523_adt_net_566364_\);
    
    \I2.PIPE6_DT_466\ : MUX2H
      port map(A => \I2.PIPE5_DTl12r_net_1\, B => 
        \I2.PIPE6_DTl12r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_466_net_1\);
    
    \I2.ROFFSET_n5_tz\ : XOR2FT
      port map(A => \I2.ROFFSETl5r_net_1\, B => 
        \I2.ROFFSET_c4_net_1\, Y => \I2.ROFFSET_n5_tz_i\);
    
    \I2.MIC_ERR_REGSl42r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_371_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl42r_net_1\);
    
    \I1.REG_15_sqmuxa_adt_net_109461_Ra1_\ : OR3FFT
      port map(A => \I1.PAGECNT_319_adt_net_854864__net_1\, B => 
        \I1.PAGECNT_320_adt_net_854872__net_1\, C => 
        \I3.PULSE_330_net_1\, Y => 
        \I1.REG_15_sqmuxa_adt_net_109461_Ra1__net_1\);
    
    \I2.MIC_REG1l3r_adt_net_834596_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_304_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1l3r_adt_net_834596_Rd1__net_1\);
    
    \I2.EVNT_NUM_n4\ : NOR2
      port map(A => EV_RES_c, B => \I2.EVNT_NUM_n4_tz_i\, Y => 
        \I2.EVNT_NUM_n4_net_1\);
    
    \I3.UN10_TCNT2_2106\ : OR2
      port map(A => \I3.TCNT2_i_0_il0r_net_1\, B => 
        \I3.TCNT2l7r_net_1\, Y => \I3.un10_tcnt2_adt_net_135288_\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__2770\ : NAND3FFT
      port map(A => \I2.ENDF_618\, B => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149__net_1\, C => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_63\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__59\);
    
    REGl369r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_270_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl369r\);
    
    \I2.DTO_1l29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_903_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l29r_net_1\);
    
    \I2.UN1_STATE3_12_I_1711\ : OR3
      port map(A => \I2.STATE3l1r_net_1\, B => \I2.N_4676\, C => 
        \I2.STATE3l13r_net_1\, Y => \I2.N_2989_adt_net_92424_\);
    
    \I1.REG_74l196r_714\ : OR2
      port map(A => \I1.REG_3_sqmuxa\, B => 
        \I1.N_65_ADT_NET_1433__218\, Y => \I1.N_65_92\);
    
    \I3.PIPEA1l16r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_314_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l16r_net_1\);
    
    \I2.N_70_adt_net_255802_\ : OAI21TTF
      port map(A => \I2.N_107_ADT_NET_256840__384\, B => 
        \I2.N_108_adt_net_54237_\, C => 
        \I2.N_70_adt_net_255801__net_1\, Y => 
        \I2.N_70_adt_net_255802__net_1\);
    
    \I3.REG_1_191\ : MUX2L
      port map(A => VDB_inl10r, B => \I3.REGl143r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, Y => 
        \I3.REG_1_191_0\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I50_Y\ : AO21
      port map(A => \I2.N276\, B => \I2.N300_0_adt_net_87051_\, C
         => \I2.N300_0_adt_net_87046_\, Y => \I2.N300_0\);
    
    \I2.DTE_2_1_0l7r\ : XOR2
      port map(A => \I2.CRC32l27r_net_1\, B => 
        \I2.CRC32l15r_net_1\, Y => \I2.DTE_2_1_0l7r_net_1\);
    
    \I2.BNCID_VECT_tile_0_WADDR_REG1l2r\ : DFF
      port map(CLK => CLK_c, D => \I2.TRGARRl2r_net_1\, Q => 
        \I2.WADDR_REG1l2r\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2275\ : AND2
      port map(A => REGl406r, B => \I3.REGMAPl55r_net_1\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146422_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I149_Y_0\ : XOR2FT
      port map(A => \I2.SUB8l12r_adt_net_855576__net_1\, B => 
        \I2.SUB8l13r_adt_net_855564__net_1\, Y => 
        \I2.ADD_18x18_fast_I149_Y_0\);
    
    \I2.PIPE3_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl10r_net_1\);
    
    \I2.PIPE10_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_607_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl2r_net_1\);
    
    \I1.REG_74_0_IV_I_A2L200R_2034\ : AND2
      port map(A => \REGl200r\, B => \I1.N_182_i\, Y => 
        \I1.N_1339_adt_net_130533_\);
    
    \I2.DT_TEMP_789\ : MUX2H
      port map(A => \I2.DT_TEMPl28r_net_1\, B => 
        \I2.DT_TEMP_7l28r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_789_net_1\);
    
    \I2.BNCID_VECTrff_10\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_10_255_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_10\);
    
    \I3.TCNT4l1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT4_387_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT4l1r_net_1\);
    
    \I2.LEAD_FLAG6l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_637_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl0r);
    
    \I2.DTE_2_1_0l9r\ : XOR2
      port map(A => \I2.CRC32l17r_net_1\, B => 
        \I2.CRC32l5r_net_1\, Y => \I2.DTE_2_1_0l9r_net_1\);
    
    \I2.WROi_10_0_0_1\ : NOR2
      port map(A => \I2.STATE2L3R_440\, B => 
        \I2.STATE2l1r_adt_net_855124__net_1\, Y => \I2.WROi_10_1\);
    
    \I2.OFFSET_37_3l6r\ : MUX2L
      port map(A => \I2.N_649\, B => \I2.N_641\, S => 
        \I2.PIPE7_DTL26R_349\, Y => \I2.N_657\);
    
    \I2.PIPE3_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl12r_net_1\);
    
    \I1.REG_74_I_O2L364R_1840\ : NOR2
      port map(A => \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_1_RD1__458\, 
        B => \I1.REG_74_i_o2_1_0_364_N_6\, Y => 
        \I1.N_661_adt_net_114476_\);
    
    \I2.STATE2_ns_i_0_o2_1l0r\ : NOR2FT
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996__net_1\, 
        B => \I2.STATE2l0r_net_1\, Y => \I2.N_4284\);
    
    \I2.LSRAM_OUTl13r_adt_net_854940_\ : BFR
      port map(A => \I2.LSRAM_OUTl13r\, Y => 
        \I2.LSRAM_OUTl13r_adt_net_854940__net_1\);
    
    \I2.L2TYPE_4_il12r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855716__net_1\, B => 
        \I2.N_4440_adt_net_67210_\, C => 
        \I2.N_4440_adt_net_67253_\, Y => \I2.N_4440\);
    
    \I1.REG_74_8_0_o4_0l380r_812\ : NAND2
      port map(A => \I1.N_1366\, B => 
        \I1.N_1367_i_adt_net_854516__net_1\, Y => \I1.N_396_190\);
    
    \I2.PIPE8_DT_21_i_1l28r_adt_net_1233_\ : OAI21
      port map(A => \I2.NWPIPE7_689\, B => \I2.PIPE7_DT_i_0l33r\, 
        C => \I2.LSRAM_OUTl28r\, Y => 
        \I2.PIPE8_DT_21_i_1l28r_adt_net_1233__net_1\);
    
    \I3.REGMAPl0r_1770\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un2_reg_ads_0_a2_0_a3_net_1\, Q => \I3.REGMAPL0R_876\);
    
    \I2.REG_1_n13\ : XOR2FT
      port map(A => \I2.N_3841_i_0\, B => \I2.REG_1_n13_0_net_1\, 
        Y => \I2.REG_1_n13_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_O2_2663\ : 
        AND3FFT
      port map(A => \I2.N_3_0_adt_net_1070__net_1\, B => 
        \I2.N_95_0\, C => \I2.N_45_1_adt_net_271427_\, Y => 
        \I2.N_45_1\);
    
    \I2.un1_tdc_res_30_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl411r, Y => 
        \I2.N_4611_i_0\);
    
    \I2.EVNT_NUMl5r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_958_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl5r_net_1\);
    
    L2A_pad : IB33
      port map(PAD => L2A, Y => L2A_c);
    
    \I2.L2ARRl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_941_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRl3r_net_1\);
    
    \I2.CRC32_12_il9r\ : OA21
      port map(A => 
        \I2.N_4667_1_adt_net_1046__adt_net_854424__net_1\, B => 
        \I2.N_56_i_0\, C => \I2.N_3926_adt_net_42578_\, Y => 
        \I2.N_3926\);
    
    TDCDB_padl15r : IB33
      port map(PAD => TDCDB(15), Y => TDCDB_cl15r);
    
    \I3.VDBOFFA_31_IV_0L0R_2629\ : AO21
      port map(A => \REGl261r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        C => \I3.VDBoffa_31l0r_adt_net_164610_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164642_\);
    
    \I2.END_CHAINA1_0_sqmuxa_i_o3\ : OAI21
      port map(A => \I2.CHAINA_EN244_i_adt_net_855260__net_1\, B
         => \I2.TOKOUTAS_net_1\, C => \I2.STATE1l11r_net_1\, Y
         => \I2.N_3273\);
    
    \I3.VDBI_13L4R_2668\ : AND3FFT
      port map(A => \I3.N_203_adt_net_24459_\, B => 
        \I3.N_203_adt_net_24461_\, C => 
        \I3.N_283_adt_net_143533_\, Y => 
        \I3.VDBi_13l4r_adt_net_284335_\);
    
    \I1.SBYTE_8_0_a2_i_m2l1r\ : MUX2L
      port map(A => \FBOUTl0r\, B => REGl84r, S => 
        \I1.sstatel2r_net_1\, Y => \I1.N_406\);
    
    \I2.OFFSET_37_23l2r\ : MUX2L
      port map(A => \REGl271r\, B => \REGl207r\, S => 
        \I2.PIPE7_DTL27R_91\, Y => \I2.N_813\);
    
    \I2.L2TYPEl10r_1547\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_599_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL10R_654\);
    
    \I4.bcnt_6\ : MUX2H
      port map(A => \I4.bcntl1r_net_1\, B => \I4.I_5\, S => 
        \I4.STATE1l1r_net_1\, Y => \I4.bcnt_6_net_1\);
    
    \I5.BITCNT_n0_i_o4\ : NOR3FTT
      port map(A => TICKL0R_555, B => \I5.N_67\, C => \I5.N_77\, 
        Y => \I5.N_73\);
    
    \I2.CRC32_12_i_0_x2l11r\ : XOR2FT
      port map(A => \I2.CRC32l11r_net_1\, B => \I2.N_228_i_i\, Y
         => \I2.N_248_i_i_0\);
    
    \I3.PIPEA1_12l10r\ : AND2
      port map(A => DPR_cl10r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854504__net_1\, Y => 
        \I3.PIPEA1_12l10r_net_1\);
    
    \I1.N_97_6_adt_net_854712_\ : BFR
      port map(A => \I1.N_97_6\, Y => 
        \I1.N_97_6_adt_net_854712__net_1\);
    
    \I2.PIPE5_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_707_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl31r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I12_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L12R_824\, B => 
        \I2.PIPE4_DTL12R_855\, Y => \I2.N_53_0\);
    
    \I1.REG_74_0_IV_I_A2L212R_2022\ : AND2
      port map(A => \REGl212r\, B => \I1.N_183_i_0\, Y => 
        \I1.N_1350_adt_net_129501_\);
    
    \I1.SBYTE_8_0_IL5R_1753\ : OA21TTF
      port map(A => \I1.N_603_i\, B => \FBOUTl4r\, C => 
        \I1.N_337\, Y => \I1.N_204_adt_net_105924_\);
    
    \I1.REG_1_209\ : MUX2H
      port map(A => \REGl308r\, B => \I1.REG_74l308r_net_1\, S
         => \I1.N_50_0_ADT_NET_1409__295\, Y => 
        \I1.REG_1_209_net_1\);
    
    \I2.SUB8_523_2742\ : AO21
      port map(A => \I2.N475_adt_net_87372_\, B => 
        \I2.SUB8_523_adt_net_566364_\, C => 
        \I2.SUB8_523_adt_net_670057_\, Y => 
        \I2.SUB8_523_adt_net_670064_\);
    
    \I2.N_3279_0_adt_net_855232_\ : BFR
      port map(A => \I2.N_3279_0_adt_net_855236__net_1\, Y => 
        \I2.N_3279_0_adt_net_855232__net_1\);
    
    \I2.DT_SRAM_0l15r\ : MUX2L
      port map(A => \I2.PIPE10_DTl15r_net_1\, B => 
        \I2.PIPE5_DTl15r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, Y => 
        \I2.N_883\);
    
    \I2.resyn_0_I2_FID_430\ : MUX2H
      port map(A => FID_cl14r, B => \I2.FID_7l14r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\, 
        Y => \I2.FID_430\);
    
    \I2.L2TYPE_4_il1r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4451_adt_net_68574_\, C => 
        \I2.N_4451_adt_net_68617_\, Y => \I2.N_4451\);
    
    \I2.CRC32_1_sqmuxa_0_a2_0_a2_0\ : OR2
      port map(A => \I2.WR_SRAM_2_ADT_NET_748__39\, B => 
        \I2.N_4273\, Y => \I2.CRC32_1_sqmuxa_0\);
    
    \I3.REGMAPl17r_adt_net_854288_\ : BFR
      port map(A => \I3.REGMAPl17r_adt_net_854300__net_1\, Y => 
        \I3.REGMAPl17r_adt_net_854288__net_1\);
    
    \I2.PIPE10_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_632_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl27r_net_1\);
    
    \I2.OFFSET_560\ : MUX2L
      port map(A => \I2.OFFSETl0r_net_1\, B => \I2.OFFSET_37l0r\, 
        S => \I2.un1_NWPIPE7_2_net_1\, Y => \I2.OFFSET_560_net_1\);
    
    \I1.REG_74_0_ivl280r\ : AO21
      port map(A => \REGl280r\, B => \I1.N_153\, C => 
        \I1.REG_74l280r_adt_net_122721_\, Y => \I1.REG_74l280r\);
    
    \I3.MBLTCYC_1160\ : DFFC
      port map(CLK => CLK_c, D => \I3.MBLTCYC_114_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.MBLTCYC_422\);
    
    \I3.STATE1_NS_0_IV_0_O2_0_I_A2_0_0_O2L7R_2086\ : NOR3
      port map(A => \I3.REGMAPL47R_448\, B => \I3.REGMAPL43R_445\, 
        C => \I3.REGMAP_I_IL46R_447\, Y => 
        \I3.N_2083_adt_net_134513_\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803_\ : OR2FT
      port map(A => \I2.TDCGDA1_net_1\, B => 
        \I2.NWPIPE1_4_SQMUXA_1_0_300\, Y => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__net_1\);
    
    \I2.ROFFSET_n7_tz\ : XOR2FT
      port map(A => \I2.ROFFSETl7r_net_1\, B => 
        \I2.ROFFSET_c6_net_1\, Y => \I2.ROFFSET_n7_tz_i\);
    
    \I3.VDBOFFB_30_IV_0L3R_2425\ : AND2
      port map(A => \REGl344r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        Y => \I3.VDBoffb_30l3r_adt_net_162524_\);
    
    \I3.REGMAPl4r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un21_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl4r_net_1\);
    
    \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__2825\ : OAI21TTF
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100__net_1\, B
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855036__net_1\, 
        C => \I2.FIRST_TDC_1_sqmuxa_net_1\, Y => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__169\);
    
    \I1.un1_sbyte13_i_i_i_a4_1_0\ : NOR2
      port map(A => \I1.sstatel9r_net_1\, B => 
        \I1.sstatel0r_net_1\, Y => \I1.N_463_1\);
    
    \I2.DTO_16_1_iv_0_x2l12r\ : XOR2
      port map(A => \I2.CRC32l8r_net_1\, B => 
        \I2.CRC32l20r_net_1\, Y => \I2.N_93_i_0\);
    
    \I1.REG_74_0_IVL312R_1904\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l312r_adt_net_119733_\);
    
    \I2.MIC_REG1L1R_2938\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_302_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1L1R_455\);
    
    \I3.STATE1_NS_0_IV_0L1R_2077\ : NOR2
      port map(A => \I3.SINGCYC_880\, B => 
        \I3.N_1905_1_adt_net_855376__net_1\, Y => 
        \I3.STATE1_nsl1r_adt_net_134330_\);
    
    \I1.REG_1_92\ : MUX2H
      port map(A => \REGl191r\, B => \I1.REG_74l191r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\, Y => 
        \I1.REG_1_92_net_1\);
    
    \I1.REG_74_0_IVL186R_2048\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l186r_adt_net_131785_\);
    
    \I3.REGMAP_i_0_il30r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un131_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il30r_net_1\);
    
    \I2.PIPE10_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_609_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl4r_net_1\);
    
    \I2.DTE_1_848\ : MUX2L
      port map(A => \I2.DTE_1l8r_Rd1__net_1\, B => 
        \I2.DTE_21_1l8r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, Y => 
        \I2.DTE_1l8r\);
    
    \I3.PULSE_331_2295\ : AND2
      port map(A => PULSEl1r, B => 
        \I3.N_1409_adt_net_854744__net_1\, Y => 
        \I3.PULSE_331_adt_net_147557_\);
    
    \I2.L2TYPE_4_IL8R_1628\ : AND2
      port map(A => \I2.L2TYPEl8r_net_1\, B => 
        \I2.N_4444_adt_net_67711_\, Y => 
        \I2.N_4444_adt_net_67754_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I161_un1_Y\ : AND3
      port map(A => \I2.N510\, B => \I2.N346_0\, C => 
        \I2.N498_1_adt_net_88035_\, Y => \I2.I161_un1_Y\);
    
    \I2.DTE_2_1l11r\ : XOR2
      port map(A => \I2.CRC32l31r_net_1\, B => 
        \I2.DTE_2_1_0l11r_net_1\, Y => \I2.DTE_2_1l11r_net_1\);
    
    \I1.PAGECNT_n9_i_i_x2\ : XOR2
      port map(A => \I1.N_325\, B => \I1.PAGECNTl9r_net_1\, Y => 
        \I1.N_404_i_i_0_i\);
    
    \I1.PAGECNTl5r_adt_net_855548_\ : BFR
      port map(A => \I1.PAGECNTl5r_net_1\, Y => 
        \I1.PAGECNTl5r_adt_net_855548__net_1\);
    
    \I3.VDBml25r\ : MUX2L
      port map(A => \I3.VDBil25r_net_1\, B => \I3.N_167\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml25r_net_1\);
    
    \I3.VDBi_57l6r_adt_net_143326_\ : AO21
      port map(A => \I3.N_2046\, B => \I3.REGl139r\, C => 
        \I3.VDBi_57l6r_adt_net_143325__net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143326__net_1\);
    
    REGl217r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_118_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl217r\);
    
    \I2.DTO_1_875\ : MUX2L
      port map(A => \I2.DTO_1l1r_net_1\, B => 
        \I2.DTO_16_1_ivl1r_net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => \I2.DTO_1_875_net_1\);
    
    \I3.REGMAPL55R_3028\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un224_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL55R_782\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2391\ : AO21
      port map(A => \REGl402r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l5r_adt_net_162124_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162168_\);
    
    TDCDB_padl16r : IB33
      port map(PAD => TDCDB(16), Y => TDCDB_cl16r);
    
    \HWRES_3_adt_net_738_\ : NAND2
      port map(A => NPWON_c, B => SYSRESB_c, Y => 
        \HWRES_3_adt_net_738__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I212_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl16r\, B => 
        \I2.PIPE7_DTl16r_net_1\, Y => 
        \I2.SUB_21x21_fast_I212_Y_0\);
    
    \I3.RAMAD_VMEl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_25_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl1r);
    
    \I3.VDBI_57_IV_0_0L2R_2262\ : OA21TTF
      port map(A => \I3.VDBi_57l2r_adt_net_145305__net_1\, B => 
        \I3.VDBi_57l2r_adt_net_145306__net_1\, C => 
        \I3.N_1905_1_adt_net_855384__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145372_\);
    
    \I1.RAMDT_SPI_e_i_0\ : INV
      port map(A => LOAD_RES, Y => \I1.LOAD_RES_i_0\);
    
    \I3.un227_reg_ads_0_a2_3_a3\ : NOR3
      port map(A => \I3.N_546\, B => \I3.N_558\, C => 
        \I3.un227_reg_ads_2\, Y => 
        \I3.un227_reg_ads_0_a2_3_a3_net_1\);
    
    \I3.N_2034_adt_net_854684_\ : BFR
      port map(A => \I3.N_2034\, Y => 
        \I3.N_2034_adt_net_854684__net_1\);
    
    \I2.sram_empty_0\ : XOR2
      port map(A => \I2.RPAGEL12R_607\, B => \I2.WPAGEL12R_752\, 
        Y => \I2.sram_empty_0_i_0_i\);
    
    \I2.TRGCNT_n0\ : XOR2
      port map(A => \I2.un9_tdctrgi_i_0\, B => 
        \I2.TRGCNT_n0_0_net_1\, Y => \I2.TRGCNT_n0_net_1\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2521\ : AO21
      port map(A => \REGl259r\, B => \I3.REGMAPl29r_net_1\, C => 
        \I3.N_2070_adt_net_163470_\, Y => 
        \I3.N_2070_adt_net_163502_\);
    
    \I2.STATE2l0r_1481\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.WPAGEe_adt_net_855056__net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.STATE2L0R_588\);
    
    \I2.LSRAM_IN_390\ : MUX2L
      port map(A => \I2.PIPE5_DTl6r_net_1\, B => 
        \I2.LSRAM_INl6r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_390_net_1\);
    
    \I2.DTO_9_ivl3r\ : OAI21TTF
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl3r_net_1\, C => 
        \I2.DTO_9_ivl3r_adt_net_34552_\, Y => 
        \I2.DTO_9_ivl3r_net_1\);
    
    \I2.BITCNT_n3_i\ : NOR3
      port map(A => \I2.ERR_WORDS_RDY_0_sqmuxa\, B => \I2.N_4336\, 
        C => \I2.N_4329\, Y => \I2.N_4324\);
    
    \I2.RAMAD_4l8r\ : MUX2L
      port map(A => \I2.N_535\, B => 
        \I1.PAGECNTl0r_adt_net_833884_Rd1__net_1\, S => LOAD_RES, 
        Y => \I2.RAMAD_4l8r_net_1\);
    
    \I2.DTESl15r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl15r, Q => 
        \I2.DTESl15r_net_1\);
    
    \I1.REG_74_2l404r_896\ : OR3FFT
      port map(A => \I1.REG_74_2_0l404r_Rd1__net_1\, B => 
        \I1.REG_74_11_a0l404r_net_1\, C => 
        \I1.N_1169_adt_net_854828__net_1\, Y => \I1.N_273_9_274\);
    
    \I3.RAMDTSl7r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl7r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl7r_net_1\);
    
    \I3.REG_1l69r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_170_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl69r);
    
    \I1.REG_17_sqmuxa_0_a2_0_a3_0_a2_842\ : NAND2
      port map(A => \I1.N_590_229\, B => 
        \I1.PAGECNTl9r_adt_net_854816__net_1\, Y => 
        \I1.N_260_220\);
    
    \I3.un37_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.un47_reg_ads_1\, B => \I3.N_637\, Y => 
        \I3.un37_reg_ads_0_a2_1_a3_net_1\);
    
    \I1.REG_1_149\ : MUX2H
      port map(A => \REGl248r\, B => \I1.REG_74l248r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_149_net_1\);
    
    \I2.PIPE3_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl3r_net_1\);
    
    \I1.REG_1_206\ : MUX2H
      port map(A => \REGl305r\, B => \I1.REG_74l305r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_206_net_1\);
    
    \I3.VDBOFFA_46_2600\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal2r_net_1\, Y => 
        \I3.VDBoffa_46_adt_net_164308_\);
    
    \I2.N_4646_1_adt_net_19635_\ : NOR2
      port map(A => \I2.MIC_REG1L3R_ADT_NET_834596_RD1__381\, B
         => \I2.MIC_REG2L3R_ADT_NET_834020_RD1__491\, Y => 
        \I2.N_4646_1_adt_net_19635__net_1\);
    
    \I2.ADEl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l10r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl10r);
    
    \I2.WOFFSET_830\ : MUX2L
      port map(A => \I2.WOFFSETl3r_Rd1__net_1\, B => 
        \I2.N_4246_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835312_Rd1__net_1\, Y
         => \I2.WOFFSETl3r\);
    
    \I2.PIPE7_DTL27R_2783\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_76\);
    
    \I2.BNCID_VECT_tile_DOUTl7r\ : MUX2L
      port map(A => \I2.DIN_REG1l7r\, B => \I2.DOUT_TMPl7r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl7r\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__3093\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__863\);
    
    \I2.DTO_16_1_IV_0L21R_1113\ : AO21
      port map(A => \I2.G_EVNT_NUMl5r_net_1\, B => \I2.N_457\, C
         => \I2.DTO_16_1l21r_adt_net_30536_\, Y => 
        \I2.DTO_16_1l21r_adt_net_30547_\);
    
    \I3.TCNT1_n4\ : XOR2
      port map(A => \I3.TCNT1l4r_net_1\, B => \I3.TCNT1_c3_net_1\, 
        Y => \I3.TCNT1_n4_net_1\);
    
    \I2.G_EVNT_NUM_n0_0_a2\ : NOR2
      port map(A => EV_RES_C_568, B => 
        \I2.G_EVNT_NUM_i_0_il0r_net_1\, Y => \I2.G_EVNT_NUM_n0\);
    
    \I1.SSTATEL8R_2977\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl2r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL8R_524\);
    
    \I2.PIPE2_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl16r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl16r_net_1\);
    
    \I1.REG_1_291\ : MUX2H
      port map(A => \REGl390r\, B => \I1.REG_74l390r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y => 
        \I1.REG_1_291_net_1\);
    
    \I3.VDBm_0l18r\ : MUX2L
      port map(A => \I3.PIPEAl18r_net_1\, B => 
        \I3.PIPEBl18r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_160\);
    
    \I1.REG_74_0_ivl404r\ : AO21
      port map(A => \REGl404r\, B => \I1.N_273\, C => 
        \I1.REG_74l404r_adt_net_109656_\, Y => 
        \I1.REG_74l404r_net_1\);
    
    \I2.END_TDC6\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_TDC6_268_net_1\, CLR
         => CLEAR_STAT_i_0, Q => END_TDC);
    
    \I3.PIPEBl16r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_95_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl16r_net_1\);
    
    \I1.N_50_0_adt_net_109756_\ : AND3FFT
      port map(A => \I1.BYTECNTl2r_adt_net_855020__net_1\, B => 
        \I1.BYTECNTl0r_net_1\, C => \I1.BYTECNTl8r_net_1\, Y => 
        \I1.N_50_0_adt_net_109756__net_1\);
    
    \I2.DTO_16_1_IVL15R_1144\ : AO21
      port map(A => \I2.DTO_1l15r\, B => \I2.N_196\, C => 
        \I2.DTO_16_1l15r_adt_net_31948_\, Y => 
        \I2.DTO_16_1l15r_adt_net_31964_\);
    
    \I3.REGMAPl23r_adt_net_855016_\ : BFR
      port map(A => \I3.REGMAPl23r_net_1\, Y => 
        \I3.REGMAPl23r_adt_net_855016__net_1\);
    
    \I2.L2TYPE_594\ : MUX2L
      port map(A => \I2.L2TYPE_i_0_il5r\, B => \I2.N_4447\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_594_net_1\);
    
    \I3.VDBi_23_0l1r\ : AND2
      port map(A => REGl81r, B => \I3.REGMAPl11r_net_1\, Y => 
        \I3.VDBi_23l1r_adt_net_145581_\);
    
    \I3.VDBoffb_30_iv_0l1r\ : AND2
      port map(A => \REGl366r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162884_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I58_Y_1680\ : AND2FT
      port map(A => \I2.LSRAM_OUTl10r\, B => 
        \I2.PIPE7_DTl10r_net_1\, Y => \I2.N308_0_adt_net_86497_\);
    
    DTO_padl23r : IOB33PH
      port map(PAD => DTO(23), A => \I2.DTO_1l23r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl23r);
    
    \I2.DT_TEMP_782\ : MUX2H
      port map(A => \I2.DT_TEMPl21r_net_1\, B => 
        \I2.DT_TEMP_7l21r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_782_net_1\);
    
    \I3.VADm_0_a3l4r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl4r_net_1\, Y => \I3.VADml4r\);
    
    \I2.PIPE9_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_292_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl23r_net_1\);
    
    \I1.REG_74_0_ivl342r\ : AO21
      port map(A => \REGl342r\, B => \I1.N_217\, C => 
        \I1.REG_74l342r_adt_net_116842_\, Y => \I1.REG_74l342r\);
    
    REGl222r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_123_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl222r\);
    
    \I2.DTO_16_1_IV_0_0L25R_1088\ : AO21
      port map(A => \I2.G_EVNT_NUMl9r_net_1\, B => \I2.N_457\, C
         => \I2.DTO_16_1l25r_adt_net_29612_\, Y => 
        \I2.DTO_16_1l25r_adt_net_29623_\);
    
    \I2.REG_1_n0_0\ : XOR2
      port map(A => REGl32r, B => \I2.N_119\, Y => 
        \I2.REG_1_n0_0_net_1\);
    
    \I2.PIPE1_DTl21r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_748_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl21r_net_1\);
    
    \I3.VDBOFFB_54_2456\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl2r_net_1\, Y => 
        \I3.VDBoffb_54_adt_net_162790_\);
    
    \I2.BITCNT_n1_i_a5\ : NOR2
      port map(A => \I2.BITCNT_c0\, B => \I2.BITCNTl1r_net_1\, Y
         => \I2.N_4334\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2396\ : AO21
      port map(A => \REGl314r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        C => \I3.VDBoffb_30l5r_adt_net_162144_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162173_\);
    
    \I2.L2TYPEl6r_1548\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_595_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL6R_655\);
    
    REGl201r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_102_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl201r\);
    
    \I2.MIC_ERR_REGS_334\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl6r_net_1\, B => 
        \I2.MIC_ERR_REGSl5r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_334_net_1\);
    
    \I1.REG_74_0_ivl355r\ : AO21
      port map(A => \REGl355r\, B => \I1.N_225\, C => 
        \I1.REG_74l355r_adt_net_115687_\, Y => \I1.REG_74l355r\);
    
    \I3.VDBOFFA_31_IV_0L5R_2534\ : AND2
      port map(A => \REGl258r\, B => \I3.REGMAPl29r_net_1\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163668_\);
    
    \I3.PIPEA_248\ : MUX2L
      port map(A => \I3.PIPEAl17r_net_1\, B => 
        \I3.PIPEA_8l17r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854664__net_1\, Y
         => \I3.PIPEA_248_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I214_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl18r\, B => 
        \I2.PIPE7_DTl18r_net_1\, Y => 
        \I2.SUB_21x21_fast_I214_Y_0\);
    
    \I2.DTO_1_877\ : MUX2L
      port map(A => \I2.DTO_1l3r_net_1\, B => 
        \I2.DTO_16_1_ivl3r_net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => \I2.DTO_1_877_net_1\);
    
    \I3.VDBi_57_ivl4r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855380__net_1\, B => 
        \I3.VDBi_43l4r_net_1\, C => 
        \I3.VDBi_57l4r_adt_net_144441_\, Y => \I3.VDBi_57l4r\);
    
    \I3.VDBI_57_IVL3R_2259\ : AO21
      port map(A => 
        \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344__net_1\, 
        B => \I3.VDBi_52l3r_net_1\, C => 
        \I3.VDBi_57l3r_adt_net_145073_\, Y => 
        \I3.VDBi_57l3r_adt_net_145074_\);
    
    MROK_pad : GL33
      port map(PAD => MROK, GL => MROK_c);
    
    \I1.REG_74l380r\ : OR3FFT
      port map(A => \I1.N_179\, B => \I1.N_185_9\, C => 
        \I1.N_249_adt_net_112440_\, Y => \I1.N_249\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I72_Y\ : AO21
      port map(A => \I2.N243_0\, B => \I2.N239\, C => \I2.N242\, 
        Y => \I2.N322\);
    
    \I2.DT_TEMP_7l18r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854240__net_1\, B => 
        \I2.DTO_16_1l18r_adt_net_756__net_1\, Y => 
        \I2.DT_TEMP_7l18r_net_1\);
    
    \I3.VDBm_0l0r\ : MUX2L
      port map(A => \I3.PIPEAl0r_net_1\, B => \I3.PIPEBl0r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_142\);
    
    \I2.TDCDASl23r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl23r, Q => 
        \I2.TDCDASl23r_net_1\);
    
    \I1.REG_74_3_i_a2l172r_900\ : NAND2FT
      port map(A => \I1.N_1370_adt_net_112317_\, B => 
        \I1.N_273_6_i_0\, Y => \I1.N_1370_278\);
    
    \I3.PIPEBl13r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_92_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl13r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I96_Y\ : NOR2
      port map(A => \I2.N307_2_865\, B => \I2.N311_0\, Y => 
        \I2.N350\);
    
    N_1_I3_TCNT3_n6 : XOR2
      port map(A => \I3.TCNT3_i_0_il6r_net_1\, B => 
        \N_1.I3.TCNT3_c5\, Y => \N_1.I3.TCNT3_n6\);
    
    REGl191r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_92_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl191r\);
    
    \I2.NWPIPE3\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE2_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE3_net_1\);
    
    \I2.PIPE10_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_619_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl14r_net_1\);
    
    \I2.LSRAM_INl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_403_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl19r_net_1\);
    
    REGl344r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_245_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl344r\);
    
    \I3.VDBI_57_0_IV_0_0L15R_2184\ : AND3FFT
      port map(A => \I3.N_2014\, B => \I3.N_1917\, C => 
        \I3.REGl148r\, Y => \I3.VDBi_57l15r_adt_net_139961_\);
    
    \I2.DTOSl31r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl31r, Q => 
        \I2.DTOS_i_il31r\);
    
    \I2.OFFSET_37_16l5r\ : MUX2L
      port map(A => \REGl266r\, B => \REGl202r\, S => 
        \I2.PIPE7_DTL27R_78\, Y => \I2.N_760\);
    
    \I5.AIR_WDATAl0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_55_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl0r_net_1\);
    
    \I3.REG_1_210\ : MUX2L
      port map(A => VDB_inl29r, B => \I3.REGl162r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\, Y => 
        \I3.REG_1_210_0\);
    
    \I1.REG_1_191\ : MUX2H
      port map(A => \REGl290r\, B => \I1.REG_74l290r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\, Y => 
        \I1.REG_1_191_net_1\);
    
    \I3.REGMAPl17r_adt_net_854284_\ : BFR
      port map(A => \I3.REGMAPl17r_adt_net_854288__net_1\, Y => 
        \I3.REGMAPl17r_adt_net_854284__net_1\);
    
    REGl329r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_230_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl329r\);
    
    \I3.VADm_0_a3l3r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl3r_net_1\, Y => \I3.VADml3r\);
    
    \I1.REG_1_208\ : MUX2H
      port map(A => \REGl307r\, B => \I1.REG_74l307r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_208_net_1\);
    
    \I3.REG3_0_sqmuxa_0_a2_0_a3_i_0\ : AND2FT
      port map(A => \I3.WRITES_net_1\, B => \I3.STATE1_IPL8R_420\, 
        Y => \I3.N_1906_i_0_0\);
    
    \I2.DTO_16_1_iv_0_o2_0_i_o2l21r_776\ : OAI21FTF
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.N_182_ADT_NET_1007__155\, Y => \I2.N_197_154\);
    
    \I3.un176_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_558\, B => \I3.N_585\, Y => 
        \I3.un176_reg_ads_0_a2_0_a3_net_1\);
    
    \I1.BYTECNT_n6_i_0\ : AND2FT
      port map(A => \I1.N_223_adt_net_854848__net_1\, B => 
        \I1.N_77_adt_net_109270_\, Y => \I1.N_77\);
    
    \I1.ISI_7_I_0_2073\ : OA21TTF
      port map(A => \I1.sstatel9r_net_1\, B => \I1.N_329\, C => 
        \I1.N_337\, Y => \I1.N_1193_adt_net_134015_\);
    
    \I3.REG_1l100r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_281_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl100r\);
    
    \I3.RAMDTSl13r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl13r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl13r_net_1\);
    
    \I3.PURGED_43\ : OA21
      port map(A => EVREAD, B => \I3.PURGED_net_1\, C => 
        \I3.un22_bltcyc\, Y => \I3.PURGED_43_net_1\);
    
    \I3.VASl15r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_77_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VAS_i_0_il15r\);
    
    \I2.WOFFSET_13_I_O2L1R_1347\ : AO21FTF
      port map(A => \I2.N_4261_304\, B => \I2.N_223_156\, C => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855000__net_1\, 
        Y => \I2.N_4262_adt_net_39852_\);
    
    \I2.TRGCNTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGCNT_n4\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGCNTl4r_net_1\);
    
    \I3.REGMAPL33R_2944\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un146_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL33R_461\);
    
    \I3.RAMDTSl1r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl1r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl1r_net_1\);
    
    \I3.VDBm_0l25r\ : MUX2L
      port map(A => \I3.PIPEAl25r_net_1\, B => 
        \I3.PIPEBl25r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_167\);
    
    \I2.PIPE8_DT_16_0l18r\ : MUX2H
      port map(A => \I2.PIPE8_DTl18r_net_1\, B => 
        \I2.PIPE7_DTl18r_net_1\, S => 
        \I2.N_565_0_adt_net_855736__net_1\, Y => \I2.N_584\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854508_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854512__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854508__net_1\);
    
    \I2.LSRAM_WR_380\ : MUX2H
      port map(A => \I2.LEAD_FLAG6_0_sqmuxa\, B => 
        \I2.LSRAM_WR_net_1\, S => END_FLUSH, Y => 
        \I2.LSRAM_WR_380_net_1\);
    
    \I2.CRC32_12_i_0l17r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_252_i_i_0\, Y => 
        \I2.N_3934\);
    
    \I1.REG_74_0_ivl298r\ : AO21
      port map(A => \REGl298r\, B => \I1.N_169\, C => 
        \I1.REG_74l298r_adt_net_121040_\, Y => \I1.REG_74l298r\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2194\ : NOR3FFT
      port map(A => REGl29r, B => \I3.N_2040\, C => \I3.N_2015\, 
        Y => \I3.VDBi_57l13r_adt_net_140499_\);
    
    \I2.L2SERV_c1\ : AND2
      port map(A => \I2.RPAGEL13R_611\, B => \I2.RPAGEL12R_608\, 
        Y => \I2.L2SERV_c1_net_1\);
    
    \I3.REGMAP_I_0_IL42R_2984\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un191_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL42R_531\);
    
    \I2.DTO_1_884\ : MUX2L
      port map(A => \I2.DTO_1l10r_Rd1__net_1\, B => 
        \I2.DTO_16_1l10r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834772_Rd1__net_1\, Y
         => \I2.DTO_1l10r\);
    
    \I2.TDCDASl5r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl5r, Q => 
        \I2.TDCDASl5r_net_1\);
    
    \I2.DT_TEMP_7l12r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854244__net_1\, B => 
        \I2.DT_SRAMl12r_net_1\, Y => \I2.DT_TEMP_7l12r_net_1\);
    
    TDCDA_padl10r : IB33
      port map(PAD => TDCDA(10), Y => TDCDA_cl10r);
    
    \I2.END_CHAINB1_709_1537\ : OAI21FTF
      port map(A => \I2.STATE1l7r_net_1\, B => 
        \I2.N_3883_adt_net_854632__net_1\, C => 
        \I2.END_CHAINB1_709_adt_net_53455_\, Y => 
        \I2.END_CHAINB1_709_adt_net_53463_\);
    
    \I3.PIPEA1_12l31r\ : AND2
      port map(A => DPR_cl31r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854484__net_1\, Y => 
        \I3.PIPEA1_12l31r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2539\ : AO21
      port map(A => \REGl282r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        C => \I3.VDBoffa_31l5r_adt_net_163660_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163692_\);
    
    \I1.REG_74_0_ivl285r\ : AO21
      port map(A => \REGl285r\, B => \I1.N_161\, C => 
        \I1.REG_74l285r_adt_net_122291_\, Y => \I1.REG_74l285r\);
    
    \I2.SUB9l11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_579_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9_i_0_il11r\);
    
    \I2.RAMAD1l6r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_660_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l6r_net_1\);
    
    \I2.L1AF3\ : DFFS
      port map(CLK => CLK_c, D => \I2.L1AF2_i_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L1AF3_i_0\);
    
    \I2.STATE3l2r_1150\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_ns_il11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3L2R_412\);
    
    \I3.REGMAP_I_0_A2L52R_2091\ : NOR3FTT
      port map(A => \I3.N_2042\, B => \I3.REGMAPl56r_net_1\, C
         => \I3.REGMAP_i_0_il5r\, Y => \I3.N_638_adt_net_134642_\);
    
    \I3.PIPEA1l23r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_321_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l23r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I33_P0N_1761\ : OR2FT
      port map(A => \I2.LSRAM_OUTl12r\, B => 
        \I2.PIPE7_DTL12R_693\, Y => \I2.N267_0_868\);
    
    \I2.PIPE5_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_679_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl3r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I166_Y\ : AND3FTT
      port map(A => \I2.N479_adt_net_296182__net_1\, B => 
        \I2.N501_i_adt_net_88539_\, C => \I2.N355_0\, Y => 
        \I2.N501_i\);
    
    \I5.COMMANDl9r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_46_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl9r_net_1\);
    
    \I3.REG_1l95r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_276_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl95r\);
    
    \I2.PIPE5_DT_6l20r\ : MUX2L
      port map(A => \I2.PIPE5_DT_6_dl20r_net_1\, B => 
        \I2.un27_pipe5_dt0l20r\, S => \I2.PIPE5_DT_6_sl19r_net_1\, 
        Y => \I2.PIPE5_DT_6l20r_net_1\);
    
    \I1.REG_74_I_O2_0_0_364_M9_I_1_1837\ : AO21
      port map(A => \I1.PAGECNTL7R_526\, B => 
        \I1.REG_74_1_a0_0l228r_adt_net_854832__net_1\, C => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854400__net_1\, 
        Y => \I1.REG_74_i_o2_0_0_364_m9_i_1_adt_net_114039_\);
    
    \I2.TDCDASl2r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl2r, Q => 
        \I2.TDCDASl2r_net_1\);
    
    \I3.VDBoffbl0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_52_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl0r_net_1\);
    
    \I3.LWORDS_3033\ : DFFC
      port map(CLK => CLK_c, D => \I3.LWORDS_61_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.LWORDS_787\);
    
    \I3.VDBil21r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_361_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil21r_net_1\);
    
    \I1.PAGECNT_323\ : MUX2H
      port map(A => \I1.PAGECNTl4r_adt_net_835120_Rd1__net_1\, B
         => \I1.PAGECNT_n4\, S => 
        \I1.PAGECNTe_adt_net_854896__net_1\, Y => 
        \I1.PAGECNT_323_net_1\);
    
    \I1.REG_1_73\ : MUX2H
      port map(A => \REGl172r\, B => \I1.REG_74l172r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\, Y
         => \I1.REG_1_73_net_1\);
    
    \I1.REG_74_0_IV_0L368R_1833\ : AND2
      port map(A => \FBOUTl3r\, B => \I1.N_593\, Y => 
        \I1.REG_74l368r_adt_net_113654_\);
    
    \I2.PIPE1_DT_42_1_IV_1L24R_1373\ : NOR2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855756__net_1\, B => 
        \I2.TDCDBSl24r_net_1\, Y => 
        \I2.PIPE1_DT_42_1_iv_1_il24r_adt_net_46469_\);
    
    \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1_\ : 
        OR3
      port map(A => \I1.PAGECNT_323_net_1\, B => 
        \I1.PAGECNT_324_net_1\, C => \I1.PAGECNT_327_net_1\, Y
         => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\);
    
    \I2.CHAINA_ERRS_524\ : MUX2L
      port map(A => \I2.CHAINA_ERRS_net_1\, B => 
        \I2.CHAINA_ERRF1_net_1\, S => 
        \I2.N_3877_adt_net_855268__net_1\, Y => 
        \I2.CHAINA_ERRS_524_net_1\);
    
    \I3.PULSEl4r_637\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_334_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEL4R_15);
    
    \I2.N_587_adt_net_1201__adt_net_855168_\ : BFR
      port map(A => \I2.N_587_adt_net_1201__net_1\, Y => 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_45387_\ : OA21FTT
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855244__net_1\, 
        B => \I2.N_3885\, C => \I2.STATE1L5R_591\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45387__net_1\);
    
    \I2.MIC_REG3_324\ : MUX2H
      port map(A => \I2.MIC_REG3l7r_net_1\, B => 
        \I2.MTDIAS_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768__net_1\, Y => 
        \I2.MIC_REG3_324_net_1\);
    
    \I1.REG_74_0_ivl177r\ : AO21
      port map(A => \REGl177r\, B => \I1.N_49\, C => 
        \I1.REG_74l177r_adt_net_132596_\, Y => \I1.REG_74l177r\);
    
    \I3.VDBOFFB_30_IV_0L3R_2428\ : AO21
      port map(A => \REGl320r\, B => \I3.REGMAPl37r_net_1\, C => 
        \I3.VDBoffb_30l3r_adt_net_162508_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162549_\);
    
    \I2.REG_1_c6_i_o2\ : OR3FFT
      port map(A => REGL37R_566, B => REGL38R_873, C => 
        \I2.N_3847\, Y => \I2.N_3849\);
    
    \I1.PAGECNTL5R_2878\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_322_adt_net_854384__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL5R_310\);
    
    \I1.REG_1_259\ : MUX2H
      port map(A => \REGl358r\, B => \I1.REG_74l358r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_259_net_1\);
    
    \I2.FID_7_0_IVL27R_981\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl27r_net_1\, 
        Y => \I2.FID_7l27r_adt_net_18833_\);
    
    \I0.BNC_RESi\ : DFFC
      port map(CLK => CLK_c, D => \I0.BNC_RESF3_net_1\, CLR => 
        \I0.un4_hwresi_i\, Q => BNC_RES_c);
    
    \I4.FLUSH_0_sqmuxa\ : NAND2
      port map(A => END_TDC, B => \I4.STATE1l2r_net_1\, Y => 
        \I4.FLUSH_0_sqmuxa_net_1\);
    
    \I2.DTO_16_1_IV_0_0L19R_1125\ : AO21
      port map(A => \I2.N_197_151\, B => \I2.DT_SRAMl19r_net_1\, 
        C => \I2.DTO_16_1l19r_adt_net_30970_\, Y => 
        \I2.DTO_16_1l19r_adt_net_30980_\);
    
    \I2.CRC32_12_i_0_m2l11r\ : MUX2H
      port map(A => \I2.DT_SRAMl11r_net_1\, B => 
        \I2.DT_TEMPl11r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854436__net_1\, Y => 
        \I2.N_228_i_i\);
    
    \I2.CRC32_1_sqmuxa_1_i_o2_924\ : OR2
      port map(A => \I2.STATE2L4R_291\, B => \I2.STATE2L3R_437\, 
        Y => \I2.N_4261_302\);
    
    \I3.PIPEBl8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_87_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl8r_net_1\);
    
    \I3.REG_1l410r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_217_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl410r);
    
    \I5.sstate1_0l13r\ : DFFS
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el0r\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l13r_net_1\);
    
    \I2.un1_PIPE1_DT_0_sqmuxa_i_0\ : OAI21
      port map(A => \I2.N_3351\, B => \I2.N_3891\, C => 
        \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\, Y => 
        \I2.N_3254\);
    
    \I1.REG_74_8_308_m6_e\ : OR2FT
      port map(A => \I1.N_299_adt_net_833868_Rd1__net_1\, B => 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__363\, Y => 
        \I1.REG_74_8_308_m6_e_net_1\);
    
    \I2.STATE3_nsl8r\ : AO21
      port map(A => \I2.N_3012\, B => 
        \I2.N_12254_i_adt_net_24491_\, C => 
        \I2.STATE3_nsl8r_adt_net_24815_\, Y => 
        \I2.STATE3_nsl8r_net_1\);
    
    \I2.PIPE9_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_291_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl22r_net_1\);
    
    \I2.PIPE7_DTL26R_2906\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_360\);
    
    \I3.REGMAP_i_0_a3l52r\ : NAND2FT
      port map(A => \I3.REGMAPl0r_net_1\, B => \I3.N_638\, Y => 
        \I3.N_437\);
    
    \I5.REG_1l419r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_32_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl419r);
    
    \I1.REG_74_0_IVL321R_1895\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l321r_adt_net_118959_\);
    
    \I1.un1_sbyte13_i_i_i\ : OA21FTF
      port map(A => \I1.N_329\, B => \I1.N_653\, C => 
        \I1.un1_sbyte13_i_i_i_1_net_1\, Y => \I1.N_1376_i_0\);
    
    N_1_I3_TCNT2_c4 : AND2
      port map(A => \I3.TCNT2_i_0_il4r_net_1\, B => \I3.TCNT2_c3\, 
        Y => \I3.TCNT2_c4\);
    
    \I1.REG_1_68\ : MUX2H
      port map(A => \REGl167r\, B => \I1.REG_74l167r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, Y => 
        \I1.REG_1_68_net_1\);
    
    REGl364r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_265_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl364r\);
    
    \I1.REG_74_12_348_M9_I_1856\ : AO21
      port map(A => \I1.REG_74_1_380_N_16\, B => 
        \I1.REG_74_12_348_m9_i_adt_net_115429_\, C => 
        \PULSE_0L0R_ADT_NET_834380_RD1__831\, Y => 
        \I1.REG_74_12_348_m9_i_adt_net_115430_\);
    
    \I1.REG_74_0_IVL337R_1879\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l337r_adt_net_117486_\);
    
    \I3.N_243_4_adt_net_1290_\ : NAND2
      port map(A => \I3.EVREAD_DS_net_1\, B => \I3.STATE2L0R_378\, 
        Y => \I3.N_243_4_adt_net_1290__net_1\);
    
    \I2.WOFFSETl7r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl7r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl7r_Rd1__net_1\);
    
    \I2.N_199_0_ADT_NET_1054__2760\ : OAI21FTT
      port map(A => \I2.STATE2L3R_440\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.DTE_CL_0_SQMUXA_2_0_286\, Y => 
        \I2.N_199_0_ADT_NET_1054__36\);
    
    \I1.REG_74_0_IVL174R_2060\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, Y => 
        \I1.REG_74l174r_adt_net_132854_\);
    
    \I2.un2_evnt_word_I_56\ : XOR2
      port map(A => \I2.WOFFSETl10r\, B => \I2.N_16_1\, Y => 
        \I2.I_56\);
    
    \I3.VDBOFFA_31_IV_0L7R_2498\ : AND2
      port map(A => \REGl284r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        Y => \I3.VDBoffa_31l7r_adt_net_163288_\);
    
    \I2.resyn_0_I2_MIC_REG1_1_sqmuxa_0_a5_0\ : AND2FT
      port map(A => COM_SERS_561, B => \I2.STATE5L2R_763\, Y => 
        \I2.MIC_REG1_1_sqmuxa_0\);
    
    \I3.UN1_NOEDTKI_0_SQMUXA_0_O3_2313\ : OA21
      port map(A => \I3.STATE1_ipl4r\, B => \I3.STATE1_ipl6r\, C
         => \I3.DSS_9\, Y => 
        \I3.un1_NOEDTKi_0_sqmuxa_adt_net_159270_\);
    
    \I2.G_EVNT_NUM_N11_0_A2_1056\ : NOR2FT
      port map(A => \I2.G_EVNT_NUMl10r_net_1\, B => 
        \I2.N_218_548\, Y => \I2.N_287_adt_net_26828_\);
    
    \I1.REG_74_0_IV_0L273R_1950\ : AND2
      port map(A => \REGl273r\, B => 
        \I1.N_145_adt_net_854772__net_1\, Y => 
        \I1.REG_74l273r_adt_net_123560_\);
    
    \I5.COMMANDl13r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_50_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl13r_net_1\);
    
    \I2.PIPE5_DT_678\ : MUX2L
      port map(A => \I2.PIPE5_DTl2r_net_1\, B => 
        \I2.PIPE5_DT_6l2r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_678_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I168_un1_Y\ : AND3FFT
      port map(A => \I2.N316_i_i\, B => \I2.N359_adt_net_86622_\, 
        C => \I2.N495_i_adt_net_202093_\, Y => \I2.I168_un1_Y\);
    
    \I2.STATE2l1r_adt_net_855120_\ : BFR
      port map(A => \I2.STATE2l1r\, Y => 
        \I2.STATE2l1r_adt_net_855120__net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_45408_\ : OAI21FTF
      port map(A => \I2.STATE1l10r_net_1\, B => \I2.N_3898_i\, C
         => \I2.STATE1_nsl11r_adt_net_23385_\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45408__net_1\);
    
    \I2.STATE2L3R_2922\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl2r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L3R_439\);
    
    \I2.DTO_16_1_iv_0_0l6r\ : OR2
      port map(A => \I2.DTO_16_1l6r_adt_net_33921_\, B => 
        \I2.DTO_16_1l6r_adt_net_33922_\, Y => \I2.DTO_16_1l6r\);
    
    \I2.DTE_1_861\ : MUX2L
      port map(A => \I2.DTE_1l23r_Rd1__net_1\, B => 
        \I2.DTE_21_1l23r_Rd1_\, S => 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\, Y => 
        \I2.DTE_1l23r\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855404_\ : BFR
      port map(A => \I1.N_50_0_adt_net_1409__net_1\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\);
    
    \I3.PIPEB_97\ : AO21
      port map(A => DPR_cl18r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\, 
        C => \I3.PIPEB_97_adt_net_159957_\, Y => 
        \I3.PIPEB_97_net_1\);
    
    \I1.REG_1_256\ : MUX2H
      port map(A => \REGl355r\, B => \I1.REG_74l355r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_256_net_1\);
    
    \I1.BYTECNT_n0_0_0\ : OAI21
      port map(A => \I1.BYTECNTl0r_net_1\, B => 
        \I1.N_223_adt_net_854844__net_1\, C => \I1.N_485\, Y => 
        \I1.BYTECNT_n0\);
    
    \I2.WOFFSET_13_il2r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_9_0\, Y => 
        \I2.N_4245\);
    
    \I1.REG_14_sqmuxa_0_a2\ : NOR2
      port map(A => 
        \I1.REG_15_sqmuxa_adt_net_1457__adt_net_854380__net_1\, B
         => \I1.N_259\, Y => \I1.REG_14_sqmuxa\);
    
    \I2.STATE1l16r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1l17r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1_i_0_il16r\);
    
    \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824_\ : BFR
      port map(A => \I2.un1_STATE3_10_1_adt_net_999__net_1\, Y
         => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\);
    
    \I3.VDBoffbl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_54_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl2r_net_1\);
    
    \I2.LEAD_FLAG6_7_i_0_a2_2l7r\ : AND2
      port map(A => \I2.PIPE5_DTL30R_622\, B => 
        \I2.PIPE5_DTl22r_net_1\, Y => \I2.N_484\);
    
    \I2.PIPE1_DT_42_1_ivl25r\ : OA21
      port map(A => \I2.PIPE1_DT_42_3_0l28r\, B => 
        \I2.EVNT_NUMl9r_net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_2l25r_net_1\, Y => 
        \I2.PIPE1_DT_42_1_iv_i_0l25r\);
    
    \I1.REG_74_0_iv_0l363r\ : AO21
      port map(A => \REGl363r\, B => \I1.N_661\, C => 
        \I1.REG_74l363r_adt_net_114611_\, Y => \I1.REG_74l363r\);
    
    \I2.WPAGEL13R_2997\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_950_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEL13R_751\);
    
    \I3.VDBi_40l10r\ : MUX2L
      port map(A => \I3.N_348\, B => \I3.N_1855\, S => 
        \I3.N_354_0_adt_net_855368__net_1\, Y => 
        \I3.VDBi_40l10r_net_1\);
    
    \I2.DTE_21_1l23r_adt_net_37285_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.DTE_21_1l23r_adt_net_37285_\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.DTE_21_1l23r_adt_net_37285_Rd1__net_1\);
    
    \I2.DTO_16_1_iv_0_o2_0_i_o2l21r_775\ : OAI21FTF
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.N_182_ADT_NET_1007__155\, Y => \I2.N_197_153\);
    
    \I5.sstate1l9r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1se_3_i_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.sstate1l9r_net_1\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855464_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__21\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\);
    
    \I2.OFFSET_37_26l5r\ : MUX2L
      port map(A => \REGl226r\, B => \I2.N_832\, S => 
        \I2.PIPE7_DTL26R_360\, Y => \I2.N_840\);
    
    \I1.REG_74_0_ivl322r\ : AO21
      port map(A => \REGl322r\, B => \I1.N_193\, C => 
        \I1.REG_74l322r_adt_net_118873_\, Y => \I1.REG_74l322r\);
    
    \I3.N_318_adt_net_855884_\ : BFR
      port map(A => \I3.N_318\, Y => 
        \I3.N_318_adt_net_855884__net_1\);
    
    \I2.PIPE8_DT_537\ : MUX2L
      port map(A => \I2.PIPE8_DTl9r_net_1\, B => 
        \I2.PIPE8_DT_21l9r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_537_net_1\);
    
    \I2.STATE2_NS_I_0_1L0R_1008\ : AND2
      port map(A => \I2.N_4261\, B => \I2.N_4273\, Y => 
        \I2.STATE2_ns_i_0_1_il0r_adt_net_21493_\);
    
    PULSEL0R_3002 : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854736__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEL0R_756);
    
    \I2.STATE5_ns_i_o2_0_o5l0r\ : AO21
      port map(A => \I2.MSERCLKS_net_1\, B => 
        \I2.STATE5l1r_net_1\, C => \I2.STATE5l2r_net_1\, Y => 
        \I2.STATE5_nsl2r\);
    
    \I1.REG_74_0_ivl353r\ : AO21
      port map(A => \REGl353r\, B => \I1.N_225\, C => 
        \I1.REG_74l353r_adt_net_115859_\, Y => \I1.REG_74l353r\);
    
    \I3.PIPEA1_12l29r\ : NAND2FT
      port map(A => DPR_cl29r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, Y => 
        \I3.PIPEA1_12l29r_net_1\);
    
    \I3.N_318_adt_net_855888_\ : BFR
      port map(A => \I3.N_318\, Y => 
        \I3.N_318_adt_net_855888__net_1\);
    
    \I1.un1_sbyte13_2_i_i_a2_i_848\ : OR2FT
      port map(A => \I1.N_436_i_i\, B => 
        \I1.N_223_adt_net_108707_\, Y => \I1.N_223_226\);
    
    \I3.REGMAPl27r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un116_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAPl27r_net_1\);
    
    \I2.FID_7_0_IVL14R_963\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl14r_net_1\, 
        Y => \I2.FID_7l14r_adt_net_17987_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I121_Y_i_o4\ : OAI21
      port map(A => \I2.N_29_i\, B => 
        \I2.ADD_21x21_fast_I121_Y_i_a3_0_i\, C => \I2.N_89\, Y
         => \I2.N_31\);
    
    \I2.LEADSRAM.M2\ : RAM256x9SST
      generic map(MEMORYFILE => "LEAD_SRAM_M2.mem")

      port map(DO8 => \I2.LSRAM_OUTl26r\, DO7 => 
        \I2.LSRAM_OUTl25r\, DO6 => \I2.LSRAM_OUTl24r\, DO5 => 
        \I2.LSRAM_OUTl23r\, DO4 => \I2.LSRAM_OUTl22r\, DO3 => 
        \I2.LSRAM_OUTl21r\, DO2 => \I2.LSRAM_OUTl20r\, DO1 => 
        \I2.LSRAM_OUTl19r\, DO0 => \I2.LSRAM_OUTl18r\, WPE => 
        OPEN, RPE => OPEN, DOS => OPEN, WADDR7 => \GND\, WADDR6
         => \GND\, WADDR5 => \GND\, WADDR4 => \GND\, WADDR3 => 
        \GND\, WADDR2 => \I2.LSRAM_WADDRl2r_net_1\, WADDR1 => 
        \I2.LSRAM_WADDRl1r_net_1\, WADDR0 => 
        \I2.LSRAM_WADDRl0r_net_1\, RADDR7 => \GND\, RADDR6 => 
        \GND\, RADDR5 => \GND\, RADDR4 => \GND\, RADDR3 => \GND\, 
        RADDR2 => \I2.LSRAM_RADDRl2r_net_1\, RADDR1 => 
        \I2.LSRAM_RADDRl1r_net_1\, RADDR0 => 
        \I2.LSRAM_RADDRl0r_net_1\, DI8 => \I2.LSRAM_INl26r_net_1\, 
        DI7 => \I2.LSRAM_INl25r_net_1\, DI6 => 
        \I2.LSRAM_INl24r_net_1\, DI5 => \I2.LSRAM_INl23r_net_1\, 
        DI4 => \I2.LSRAM_INl22r_net_1\, DI3 => 
        \I2.LSRAM_INl21r_net_1\, DI2 => \I2.LSRAM_INl20r_net_1\, 
        DI1 => \I2.LSRAM_INl19r_net_1\, DI0 => 
        \I2.LSRAM_INl18r_net_1\, WRB => \I2.LSRAM_WR_net_1\, RDB
         => \I2.LSRAM_RD_net_1\, WBLKB => \GND\, RBLKB => \GND\, 
        PARODD => \GND\, WCLKS => CLK_c, RCLKS => CLK_c, DIS => 
        \GND\);
    
    \I1.REG_74_0_iv_0_0_o2_245_m6_i_0_0\ : AND2
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        B => \I1.PAGECNTl6r_adt_net_854928__net_1\, Y => 
        \I1.REG_74_1_404_m7_i_a5_0_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2386\ : AND2
      port map(A => \REGl378r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162132_\);
    
    \I2.DTO_16_1_IVL14R_1151\ : AO21
      port map(A => \I2.DTO_1l14r\, B => \I2.N_196\, C => 
        \I2.DTO_16_1l14r_adt_net_32194_\, Y => 
        \I2.DTO_16_1l14r_adt_net_32210_\);
    
    \I2.SUB8_505\ : MUX2H
      port map(A => \I2.SUB8l2r_net_1\, B => \I2.SUB8_2l2r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855136__net_1\, Y => 
        \I2.SUB8_505_net_1\);
    
    \I1.REG_74_0_IV_0L366R_1835\ : AND2
      port map(A => \FBOUTl1r\, B => \I1.N_593\, Y => 
        \I1.REG_74l366r_adt_net_113826_\);
    
    FID_padl9r : OB33PH
      port map(PAD => FID(9), A => FID_cl9r);
    
    \I2.DTE_21_1_IVL14R_1281\ : OR3
      port map(A => \I2.DTO_16_1l14r_adt_net_32202_\, B => 
        \I2.DTE_21_1l14r_adt_net_38061_\, C => 
        \I2.DTE_21_1l14r_adt_net_38068_\, Y => 
        \I2.DTE_21_1l14r_adt_net_38070_\);
    
    \I1.REG_74L220R_2008\ : AND3
      port map(A => \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, 
        B => \I1.REG_74_1_a0_0l228r_adt_net_854832__net_1\, C => 
        \I1.REG_74_5_404_m1_e_0_net_1\, Y => 
        \I1.N_89_adt_net_128728_\);
    
    \I2.DTE_21_1l8r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l8r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l8r_Rd1__net_1\);
    
    \I2.STATE3l2r_1152\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_ns_il11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3L2R_414\);
    
    \I3.REG_1_291\ : MUX2L
      port map(A => VDB_inl9r, B => REGl110r, S => 
        \I3.N_318_adt_net_855888__net_1\, Y => \I3.REG_1_291_0\);
    
    \I2.G_EVNT_NUM_n11_0\ : NAND2FT
      port map(A => \I2.G_EVNT_NUM_n11_adt_net_26872_\, B => 
        \I2.N_287\, Y => \I2.G_EVNT_NUM_n11\);
    
    \I3.VDBi_43l5r\ : MUX2L
      port map(A => REGl411r, B => \I3.VDBi_40l5r\, S => 
        \I3.REGMAPl55r_net_1\, Y => \I3.VDBi_43l5r_net_1\);
    
    \I2.DTE_21_1_0_iv_0_0l29r\ : AO21
      port map(A => \I2.DTE_1l29r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\, C => 
        \I2.DTE_21_1l29r_adt_net_36651_\, Y => \I2.DTE_21_1l29r\);
    
    \I3.un1_STATE2_6_1_adt_net_1481_\ : NAND2FT
      port map(A => \I3.STATE2l2r_net_1\, B => \I3.N_1896\, Y => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\);
    
    \I2.MIC_ERR_REGS_341\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl13r_net_1\, B => 
        \I2.MIC_ERR_REGSl12r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\, Y => 
        \I2.MIC_ERR_REGS_341_net_1\);
    
    \I2.FIDl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_439\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl23r);
    
    \I2.MIC_ERR_REGS_349\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl21r_net_1\, B => 
        \I2.MIC_ERR_REGSl20r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_349_net_1\);
    
    \I3.VDBI_57_0_IV_0L20R_2168\ : AND2
      port map(A => \I3.PIPEAl20r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l20r_adt_net_139285_\);
    
    \I1.PAGECNT_n6_i_i_a2\ : AND2FT
      port map(A => \I1.PAGECNTl6r_adt_net_854924__net_1\, B => 
        \I1.PAGECNTl5r_net_1\, Y => \I1.N_590\);
    
    \I2.G_EVNT_NUM_n2_i_0\ : AND3FFT
      port map(A => EV_RES_C_569, B => \I2.N_316_i\, C => 
        \I2.N_187\, Y => \I2.N_4342\);
    
    \I2.un8_evread_1_adt_net_855788_\ : BFR
      port map(A => \I2.un8_evread_1_adt_net_855792__net_1\, Y
         => \I2.un8_evread_1_adt_net_855788__net_1\);
    
    \I2.PIPE1_DTl25r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_752_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl25r_net_1\);
    
    \I3.REG_1l144r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_192_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl144r\);
    
    \I1.REG_0_sqmuxa_i_0_a2_645\ : AND3
      port map(A => \I1.SSTATEL0R_307\, B => \I1.N_324_25\, C => 
        \I1.BITCNTL2R_753\, Y => \I1.N_598_23\);
    
    REGl281r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_182_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl281r\);
    
    \I5.REG_12l431r\ : AND2
      port map(A => \I5.TEMP_ACK_net_1\, B => REGl118r, Y => 
        \I5.REG_12l431r_net_1\);
    
    \I2.resyn_0_I2_FID_447\ : MUX2H
      port map(A => FID_cl31r, B => \I2.FID_7l31r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\, 
        Y => \I2.FID_447\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604_\ : BFR
      port map(A => \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\, Y
         => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\);
    
    \I2.DTE_cl_0_sqmuxa_2_0_a2_0_a2_0_911\ : OR2FT
      port map(A => \I2.N_4241_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, Y => 
        \I2.DTE_CL_0_SQMUXA_2_0_289\);
    
    \I3.REG3_130\ : MUX2L
      port map(A => VDB_inl5r, B => \I3.REG3l5r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855624__net_1\, Y => 
        \I3.REG3_130_net_1\);
    
    \I3.VAS_75\ : MUX2L
      port map(A => VAD_inl13r, B => \I3.VAS_i_0_il13r\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_75_net_1\);
    
    \I2.PIPE3_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl11r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I120_Y_0_1588\ : AND2
      port map(A => \I2.N_89_0\, B => \I2.N_84_0\, Y => 
        \I2.N531_0_adt_net_60100_\);
    
    \I2.PIPE7_DTl11r_1587\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL11R_694\);
    
    \I2.DTO_1_878\ : MUX2L
      port map(A => \I2.DTO_1l4r_Rd1__net_1\, B => 
        \I2.DTO_16_1l4r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834776_Rd1__net_1\, Y
         => \I2.DTO_1l4r\);
    
    \I3.VDBoffal2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_46_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal2r_net_1\);
    
    \I1.REG_1_258\ : MUX2H
      port map(A => \REGl357r\, B => \I1.REG_74l357r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_258_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I26_G0N\ : AND2FT
      port map(A => \I2.LSRAM_OUTl5r\, B => \I2.PIPE7_DTL5R_700\, 
        Y => \I2.N245\);
    
    \I2.NWRSRAME\ : OR2
      port map(A => \I2.CLK_sram\, B => \I2.WREi_net_1\, Y => 
        NWRSRAME_c);
    
    \I2.un1_STATE1_31_i\ : OR2
      port map(A => \I2.N_3875_i_0\, B => 
        \I2.N_3866_adt_net_61369_\, Y => \I2.N_3866\);
    
    \I2.RAMDT4L5R_3056\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_810\);
    
    \I2.END_TDC1_1_sqmuxa_i_o3_802\ : OR2
      port map(A => \I2.TOKOUT_FL_644\, B => \I2.TOKOUTBS_163\, Y
         => \I2.N_3879_180\);
    
    \I2.ADOl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l10r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl10r);
    
    \I5.TEMPDATA_80\ : MUX2L
      port map(A => \I5.TEMPDATAl6r_net_1\, B => REGl131r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_80_net_1\);
    
    \I5.SBYTE_9_1l0r\ : MUX2L
      port map(A => \I5.COMMANDl8r_net_1\, B => 
        \I5.SBYTE_9l0r_adt_net_11050_\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.SBYTE_9l0r\);
    
    \I3.ASBSF1\ : DFFS
      port map(CLK => CLK_c, D => ASB_c, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.ASBSF1_net_1\);
    
    \I2.N_4253_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4253\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4253_Rd1__net_1\);
    
    \I3.REG1l405r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG1_227_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l405r_net_1\);
    
    \I2.PIPE5_DT_6_0l3r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l3r\, B => 
        \I2.un27_pipe5_dt0l3r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1072\);
    
    \I1.REG_74_3L404R_1839\ : AO21FTT
      port map(A => \I1.PAGECNTL7R_526\, B => \I1.N_127_i\, C => 
        \I1.N_1169_adt_net_854828__net_1\, Y => 
        \I1.N_273_10_adt_net_114361_\);
    
    \I1.REG_1_231\ : MUX2H
      port map(A => \REGl330r\, B => \I1.REG_74l330r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y => 
        \I1.REG_1_231_net_1\);
    
    \I2.CHA_DATA8_502\ : MUX2L
      port map(A => \I2.CHA_DATA8_net_1\, B => \I2.N_4398\, S => 
        \I2.NWPIPE7_net_1\, Y => \I2.CHA_DATA8_502_net_1\);
    
    \I2.DTE_21_1_IVL14R_1279\ : AND2FT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_288\, B => 
        \I2.DT_SRAMl14r_net_1\, Y => 
        \I2.DTE_21_1l14r_adt_net_38061_\);
    
    \I5.PULSE_FL\ : DFFC
      port map(CLK => CLK_c, D => \I5.PULSE_FL_53_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.PULSE_FL_net_1\);
    
    \I2.N_4255_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4255\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4255_Rd1__net_1\);
    
    \I2.DTOSl23r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl23r, Q => 
        \I2.DTOSl23r_net_1\);
    
    \I2.STATE1_ns_o3_i_a2l1r\ : OAI21TTF
      port map(A => \I2.N_3279_0\, B => \I2.ERR_WORDS_RDY_net_1\, 
        C => \I2.STATE1l1r_net_1\, Y => \I2.N_3798\);
    
    \I2.DTE_21_1_IV_0L5R_1326\ : AND2FT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_287\, B => 
        \I2.DT_SRAMl5r_net_1\, Y => 
        \I2.DTE_21_1l5r_adt_net_39091_\);
    
    \I3.VDBOFFB_30_IV_0L4R_2403\ : AND2
      port map(A => \REGl353r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162318_\);
    
    \I3.REG_1l136r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_184_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl136r\);
    
    \I2.DTE_21_1_IV_0L19R_1267\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.G_EVNT_NUMl3r_net_1\, 
        C => \I2.DTE_21_1l19r_adt_net_37713_\, Y => 
        \I2.DTE_21_1l19r_adt_net_37724_\);
    
    N_1_I3_TCNT2_c6 : NAND2
      port map(A => \I3.TCNT2_i_0_il6r_net_1\, B => 
        \N_1.I3.TCNT2_c5\, Y => \N_1.I3.TCNT2_c6\);
    
    \I2.L1AF2\ : DFFC
      port map(CLK => CLK_c, D => \I2.L1AF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L1AF2_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I139_Y_i_a4\ : NAND3FFT
      port map(A => \I2.N_16\, B => \I2.N_75_adt_net_54671_\, C
         => \I2.N_66\, Y => \I2.N_96_adt_net_481750_\);
    
    \I2.PIPE6_DT_463\ : MUX2H
      port map(A => \I2.PIPE5_DTl9r_net_1\, B => 
        \I2.PIPE6_DTl9r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_463_net_1\);
    
    \I2.DTO_16_1_IV_0L20R_1118\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.G_EVNT_NUMl4r_net_1\, Y
         => \I2.DTO_16_1l20r_adt_net_30786_\);
    
    \I1.sstatel5r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_ns_il5r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel5r_net_1\);
    
    \I2.OFFSETl2r_1571\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_562_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL2R_678\);
    
    \I1.REG_74_0_IVL319R_1897\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l319r_adt_net_119131_\);
    
    \I2.MIC_REG1_306\ : MUX2H
      port map(A => \I2.MIC_REG1l5r_net_1\, B => 
        \I2.MIC_REG1_i_il6r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG1_306_net_1\);
    
    \I2.FID_7_0_ivl21r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl21r_net_1\, 
        C => \I2.FID_7l21r_adt_net_19405_\, Y => \I2.FID_7l21r\);
    
    \I2.RAMAD1_656\ : MUX2L
      port map(A => \I2.RAMAD1_12l2r_net_1\, B => 
        \I2.RAMAD1l2r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__173\, Y => 
        \I2.RAMAD1_656_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2394\ : AO21
      port map(A => \REGl298r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l5r_adt_net_162136_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162171_\);
    
    \I1.REG_74_0_ivl400r\ : AO21
      port map(A => \REGl400r\, B => \I1.N_273\, C => 
        \I1.REG_74l400r_adt_net_110100_\, Y => \I1.REG_74l400r\);
    
    TDCDA_padl8r : IB33
      port map(PAD => TDCDA(8), Y => TDCDA_cl8r);
    
    \I2.PIPE9_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_298_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl29r_net_1\);
    
    \I3.REGMAPl31r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un136_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAPl31r_net_1\);
    
    \I3.VDBi_29_0_a3_1l5r\ : AND3FFT
      port map(A => \I3.REGMAPl14r_net_1\, B => \I3.N_1907\, C
         => \I3.N_282_i_i\, Y => \I3.N_1948\);
    
    \I1.REG_74_0_IV_I_A2L197R_2037\ : AND2
      port map(A => \REGl197r\, B => \I1.N_182_i\, Y => 
        \I1.N_129_adt_net_130791_\);
    
    \I2.SRAM_EVNT_n0\ : XOR2FT
      port map(A => \I2.N_128_1\, B => \I2.SRAM_EVNT_n0_0_net_1\, 
        Y => \I2.SRAM_EVNT_n0_net_1\);
    
    \I1.REG_74_0_ivl237r\ : AO21
      port map(A => \REGl237r\, B => \I1.N_113\, C => 
        \I1.REG_74l237r_adt_net_126985_\, Y => \I1.REG_74l237r\);
    
    \I2.PIPE1_DT_42_1_IVL12R_1449\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044__net_1\, 
        B => \I2.PIPE1_DT_12l12r_net_1\, Y => 
        \I2.PIPE1_DT_42l12r_adt_net_49442_\);
    
    \I3.REG_1_sqmuxa_3_adt_net_855340_\ : BFR
      port map(A => \I3.REG_1_sqmuxa_3\, Y => 
        \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\);
    
    \I2.FID_7_0_IVL10R_972\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl58r, C => 
        \I2.FID_7l10r_adt_net_18363_\, Y => 
        \I2.FID_7l10r_adt_net_18371_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I105_Y\ : AND2FT
      port map(A => \I2.N320\, B => \I2.N317\, Y => 
        \I2.N359_adt_net_86622_\);
    
    \I2.SUB8l8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_511_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l8r_net_1\);
    
    \I2.PIPE4_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl13r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl13r_net_1\);
    
    \I2.PIPE1_DTl24r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_751_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl24r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2593\ : AO21
      port map(A => \REGl279r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        C => \I3.VDBoffa_31l2r_adt_net_164230_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164262_\);
    
    \I2.BNCID_VECTrff_13\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_13_252_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_13\);
    
    \I2.EVNT_WORD_723\ : MUX2H
      port map(A => \I2.EVNT_WORDl10r_net_1\, B => \I2.I_56\, S
         => \I2.N_2864_0_adt_net_854272__net_1\, Y => 
        \I2.EVNT_WORD_723_net_1\);
    
    \I2.sram_empty_2\ : XOR2
      port map(A => \I2.RPAGEL14R_615\, B => \I2.WPAGEL14R_750\, 
        Y => \I2.sram_empty_2_i_0_i\);
    
    \I1.sstate_tr29_0_a2_0_a4\ : AND2FT
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.sstatel1r_net_1\, Y => \I1.sstate_ns_il10r\);
    
    \I2.WOFFSET_13_il10r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_56\, Y => \I2.N_4253\);
    
    \I2.RAMAD1_664\ : MUX2L
      port map(A => \I2.RAMAD1_12l10r_net_1\, B => 
        \I2.RAMAD1l10r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__171\, Y => 
        \I2.RAMAD1_664_net_1\);
    
    DTO_padl1r : IOB33PH
      port map(PAD => DTO(1), A => \I2.DTO_1l1r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl1r);
    
    \I2.CRC32_12_i_0_x2l19r\ : XOR2FT
      port map(A => \I2.CRC32l19r_net_1\, B => \I2.N_229_i_i\, Y
         => \I2.N_247_i_i_0\);
    
    \I1.REG_1_131\ : MUX2H
      port map(A => \REGl230r\, B => \I1.REG_74l230r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\, Y => 
        \I1.REG_1_131_net_1\);
    
    \I1.REG_74_2_3l228r\ : OAI21TTF
      port map(A => \I1.N_253\, B => 
        \I1.REG_74_24_404_m3_e_net_1\, C => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536__net_1\, 
        Y => \I1.REG_74_2_3_il228r\);
    
    \I2.PIPE8_DT_535\ : MUX2L
      port map(A => \I2.PIPE8_DTl7r_net_1\, B => 
        \I2.PIPE8_DT_21l7r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_535_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2397\ : AO21
      port map(A => \REGl338r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l5r_adt_net_162148_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162174_\);
    
    \I3.TCNT1_n1\ : XOR2
      port map(A => \I3.TCNT1l0r_net_1\, B => 
        \I3.TCNT1_i_0_il1r_net_1\, Y => \I3.TCNT1_n1_net_1\);
    
    RAMDT_padl13r : IOB33PH
      port map(PAD => RAMDT(13), A => \I1.RAMDT_SPI_1l6r_net_1\, 
        EN => \I1.RAMDT_SPI_E_0\, Y => RAMDT_inl13r);
    
    \I2.FID_7_0_ivl16r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl16r_net_1\, 
        C => \I2.FID_7l16r_adt_net_17807_\, Y => \I2.FID_7l16r\);
    
    \I3.VDBil3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_343_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil3r_net_1\);
    
    \I2.NOESRAMO\ : DFFS
      port map(CLK => CLK_c, D => NOESRAME_c, SET => 
        CLEAR_STAT_i_0, Q => NOESRAMO_c);
    
    \I3.VDBOFFB_30_IV_0L0R_2481\ : AO21
      port map(A => \REGl397r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l0r_adt_net_163074_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163118_\);
    
    DTE_padl10r : IOB33PH
      port map(PAD => DTE(10), A => \I2.DTE_1l10r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl10r);
    
    \I1.REG_20_sqmuxa_adt_net_855484_\ : BFR
      port map(A => \I1.REG_20_sqmuxa\, Y => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\);
    
    \I1.PAGECNT_n6_i_i_a2_850\ : AND2FT
      port map(A => \I1.PAGECNTl6r_adt_net_854932__net_1\, B => 
        \I1.PAGECNTL5R_311\, Y => \I1.N_590_228\);
    
    DS1B_pad : IB33
      port map(PAD => DS1B, Y => DS1B_c);
    
    REGl324r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_225_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl324r\);
    
    \I2.CHAINA_EN244_i_adt_net_855264_\ : BFR
      port map(A => \I2.CHAINA_EN244_i\, Y => 
        \I2.CHAINA_EN244_i_adt_net_855264__net_1\);
    
    \I1.un1_sbyte13_1_i_0_s_831\ : AO21
      port map(A => \I1.N_370_adt_net_854904__net_1\, B => 
        \I1.un1_sbyte13_1_i_1_adt_net_106369__adt_net_854528__net_1\, 
        C => \PULSE_0L0R_ADT_NET_834380_RD1__199\, Y => 
        \I1.UN1_SBYTE13_1_I_1_209\);
    
    \I1.REG_74_0_IV_0_0L248R_1978\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l248r_adt_net_125949_\);
    
    \I2.PIPE3_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl16r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl16r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL21R_1385\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855032__net_1\, 
        B => \I2.TDCDASl21r_net_1\, Y => 
        \I2.PIPE1_DT_42l21r_adt_net_46859_\);
    
    \I2.PIPE1_DT_30l3r\ : MUX2L
      port map(A => \I2.TDCDBSl3r_net_1\, B => 
        \I2.TDCDBSl1r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, Y
         => \I2.PIPE1_DT_30l3r_net_1\);
    
    \I3.VDBi_43l4r\ : MUX2L
      port map(A => REGl410r, B => \I3.VDBi_40l4r_net_1\, S => 
        \I3.REGMAPl55r_net_1\, Y => \I3.VDBi_43l4r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I141_Y_0\ : XOR2
      port map(A => \I2.ca_0_and2\, B => \I2.G_1_4\, Y => 
        \I2.ADD_18x18_fast_I141_Y_0\);
    
    \I2.DTO_16_1_IVL11R_1166\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854624__net_1\, 
        B => \I2.DT_TEMPl11r_net_1\, C => 
        \I2.DTO_16_1l11r_adt_net_32872_\, Y => 
        \I2.DTO_16_1l11r_adt_net_32878_\);
    
    \I5.un1_BITCNT_1_sqmuxa_i_1_0_o4\ : NAND3FFT
      port map(A => \I5.N_75\, B => \I5.N_71\, C => \I5.N_70\, Y
         => \I5.N_94\);
    
    \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855280_\ : BFR
      port map(A => \I3.un1_STATE2_7_1_adt_net_1473__net_1\, Y
         => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855280__net_1\);
    
    \I2.un21_pipe5_dt_1\ : XOR2
      port map(A => \I2.RAMDT4l2r_net_1\, B => 
        \I2.RAMDT4l1r_net_1\, Y => \I2.un21_pipe5_dt_1_net_1\);
    
    \I2.DTO_1_902\ : MUX2L
      port map(A => \I2.DTO_1l28r_net_1\, B => 
        \I2.DTO_16_1_ivl28r_net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => \I2.DTO_1_902_net_1\);
    
    \I1.REG_74_3_4L380R_1943\ : OAI21FTF
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854404__net_1\, 
        B => \I1.PAGECNTl6r_net_1\, C => 
        \PULSE_0L0R_ADT_NET_834380_RD1__832\, Y => 
        \I1.REG_74_3_4_il380r_adt_net_123085_\);
    
    \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828_\ : BFR
      port map(A => \I2.un1_STATE3_10_1_adt_net_999__net_1\, Y
         => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\);
    
    \I2.L2ARRl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_942_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRl2r_net_1\);
    
    \I1.PAGECNT_n6_i_i_a4_0_828\ : OR2FT
      port map(A => \I1.UN1_SBYTE13_1_I_1_210\, B => 
        \I1.N_656_494\, Y => \I1.N_473_206\);
    
    \I3.REG_1_173\ : MUX2L
      port map(A => VDB_inl24r, B => REGl72r, S => 
        \I3.N_1935_adt_net_855320__net_1\, Y => \I3.REG_1_173_0\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I204_Y\ : XOR2
      port map(A => \I2.I168_un1_Y\, B => 
        \I2.SUB_21x21_fast_I204_Y_0\, Y => \I2.SUB8_2_i_i_0l8r\);
    
    \I2.PIPE1_DT_736\ : MUX2L
      port map(A => \I2.PIPE1_DTl9r_net_1\, B => 
        \I2.PIPE1_DT_42l9r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854580__net_1\, 
        Y => \I2.PIPE1_DT_736_net_1\);
    
    \I2.DTESl27r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl27r, Q => 
        \I2.DTESl27r_net_1\);
    
    \I2.BNCID_VECTrff_2\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_2_263_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_2\);
    
    \I1.REG_1_sqmuxa_0_a2_3_0_a4\ : OR2
      port map(A => \I1.PAGECNTL9R_492\, B => \I1.PAGECNTL6R_247\, 
        Y => \I1.N_237\);
    
    \I2.N_4646_1_adt_net_1645_Ra1_\ : OAI21TTF
      port map(A => \I2.MIC_REG1_304_net_1\, B => 
        \I2.MIC_REG2_312_net_1\, C => 
        \I2.N_4646_1_adt_net_19637_Ra1__net_1\, Y => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\);
    
    \I3.VDBi_346\ : MUX2L
      port map(A => \I3.VDBil6r_net_1\, B => \I3.VDBi_57l6r\, S
         => \I3.un1_STATE1_13_1_adt_net_1351__net_1\, Y => 
        \I3.VDBi_346_net_1\);
    
    \I2.dataout_0_adt_net_855800_\ : BFR
      port map(A => \I2.dataout_0\, Y => 
        \I2.dataout_0_adt_net_855800__net_1\);
    
    \I3.PIPEA1_299\ : MUX2L
      port map(A => \I3.PIPEA1l1r_net_1\, B => 
        \I3.PIPEA1_12l1r_net_1\, S => 
        \I3.un1_STATE2_15_1_adt_net_1342__net_1\, Y => 
        \I3.PIPEA1_299_net_1\);
    
    \I2.un1_STATE2_15_i_0_a2_1_i_678\ : NAND2
      port map(A => \I2.STATE2L5R_508\, B => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__59\, Y => 
        \I2.N_4641_56\);
    
    \I1.REG_74_0_iv_0_0l250r\ : AO21
      port map(A => \REGl250r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l250r_adt_net_125777_\, Y => \I1.REG_74l250r\);
    
    \I2.L2TYPE_4_i_o2_0l2r\ : NOR2
      port map(A => \I2.L2ARRl3r_net_1\, B => \I2.L2ARRl2r_net_1\, 
        Y => \I2.N_4461\);
    
    \I2.RAMAD_4l1r\ : MUX2L
      port map(A => \I2.N_528\, B => \I1.BYTECNT_i_0_il1r_net_1\, 
        S => LOAD_RES, Y => \I2.RAMAD_4l1r_net_1\);
    
    \I2.DTE_21_1_iv_0_0l17r\ : OR3
      port map(A => \I2.DTE_21_1l17r_adt_net_36142_\, B => 
        \I2.DTE_21_1l17r_adt_net_36153_\, C => 
        \I2.DTE_21_1l17r_adt_net_36154_\, Y => \I2.DTE_21_1l17r\);
    
    \I2.UN1_REG80_I_1697\ : NOR2
      port map(A => REGl45r, B => REGl43r, Y => 
        \I2.N_3824_adt_net_90287_\);
    
    \I2.STATE1l13r_1494\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_il5r_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.STATE1L13R_601\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I96_Y_1757\ : NOR2
      port map(A => \I2.N307_2_865\, B => \I2.N311_0\, Y => 
        \I2.N350_864\);
    
    \I2.PIPE8_DT_16_0l1r\ : MUX2H
      port map(A => \I2.PIPE8_DTl1r_net_1\, B => 
        \I2.PIPE7_DTl1r_net_1\, S => 
        \I2.N_565_0_adt_net_855728__net_1\, Y => \I2.N_567\);
    
    \I2.PIPE8_DT_21l7r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl7r\, B => \I2.N_573\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l7r_net_1\);
    
    \I2.PIPE4_DTl12r_1250_1750\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL12R_857\);
    
    \I1.REG_74_0_IVL374R_1825\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l374r_adt_net_113001_\);
    
    \I2.DTE_21_1_0_ivl30r\ : AOI21FTT
      port map(A => \I2.DTE_1l30r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, C => 
        \I2.DTE_21_1_0_iv_1l30r_net_1\, Y => 
        \I2.DTE_21_1_0_ivl30r_net_1\);
    
    \I1.PAGECNTlde_0_o2_2\ : NAND2FT
      port map(A => \I1.N_310_RD1__335\, B => 
        \I1.N_311_I_I_RD1__762\, Y => \I1.N_325\);
    
    \I5.REG_1_34\ : MUX2L
      port map(A => \I5.TEMPDATAl1r_net_1\, B => REGl421r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_34_net_1\);
    
    \I3.TCNTl0r_1166\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_384_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTL0R_428\);
    
    \I2.EVNT_NUM_961\ : MUX2L
      port map(A => \I2.EVNT_NUMl2r_net_1\, B => 
        \I2.EVNT_NUM_n2_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_961_net_1\);
    
    \I3.REGMAP_I_0_A2L52R_2090\ : NOR2
      port map(A => \I3.REGMAPL10R_719\, B => \I3.REGMAPL1R_724\, 
        Y => \I3.N_638_adt_net_134639_\);
    
    \I2.TDCDBSl7r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl7r, Q => 
        \I2.TDCDBSl7r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I152_Y_0_2710\ : NOR2FT
      port map(A => \I2.N498_0_adt_net_56939_\, B => 
        \I2.N502_i_0_adt_net_490392_\, Y => 
        \I2.N498_0_adt_net_598283_\);
    
    \I2.PIPE1_DT_734\ : MUX2L
      port map(A => \I2.PIPE1_DTl7r_net_1\, B => 
        \I2.PIPE1_DT_42l7r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854584__net_1\, 
        Y => \I2.PIPE1_DT_734_net_1\);
    
    \I2.EVNT_WORD_724\ : MUX2H
      port map(A => \I2.EVNT_WORDl11r_net_1\, B => \I2.I_66\, S
         => \I2.N_2864_0_adt_net_854268__net_1\, Y => 
        \I2.EVNT_WORD_724_net_1\);
    
    \I2.DTE_cl_5l31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4180_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_cll31r\);
    
    \I2.BNCID_VECT_tile_I_6_2\ : XOR2
      port map(A => \I2.TRGSERVl2r_net_1\, B => 
        \I2.WADDR_REG1l2r\, Y => \I2.I_6_2_i_0_i\);
    
    \I3.REG_1_199\ : MUX2L
      port map(A => VDB_inl18r, B => \I3.REGl151r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\, Y => 
        \I3.REG_1_199_0\);
    
    \I2.REG_1l80r\ : DFFC
      port map(CLK => MWOK_c, D => \VCC\, CLR => \I2.un8_hwres_i\, 
        Q => REGl80r);
    
    \I2.FIRST_TDC_1_sqmuxa_1_0_922\ : OR2FT
      port map(A => \I2.STATE1L12R_645\, B => 
        \I2.END_CHAINA1_1_sqmuxa_3\, Y => 
        \I2.NWPIPE1_4_SQMUXA_1_0_300\);
    
    \I2.OFFSET_37_14l7r\ : MUX2L
      port map(A => \I2.N_738\, B => \I2.N_690\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_746\);
    
    \I2.FID_7_0_IVL11R_970\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl59r, C => 
        \I2.FID_7l11r_adt_net_18269_\, Y => 
        \I2.FID_7l11r_adt_net_18277_\);
    
    \I2.LSRAM_INl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_393_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl9r_net_1\);
    
    \I3.VDBi_57_0_iv_0l9r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855380__net_1\, B => 
        \I3.VDBi_43l9r_net_1\, C => 
        \I3.VDBi_57l9r_adt_net_142332_\, Y => \I3.VDBi_57l9r\);
    
    \I2.ROFFSET_914\ : MUX2H
      port map(A => \I2.ROFFSETl4r_net_1\, B => 
        \I2.ROFFSET_n4_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_914_net_1\);
    
    \I2.WOFFSETl0r_adt_net_854648_\ : BFR
      port map(A => \I2.WOFFSETl0r_net_1\, Y => 
        \I2.WOFFSETl0r_adt_net_854648__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0_o2_1_947\ : 
        OR3FFT
      port map(A => \I2.N_107_0\, B => \I2.N_13_1\, C => 
        \I2.N_95_0\, Y => \I2.N_74_ADT_NET_55281__325\);
    
    \I1.REG_28_sqmuxa_0_a2\ : NOR2
      port map(A => 
        \I1.REG_15_sqmuxa_adt_net_1457__adt_net_854380__net_1\, B
         => \I1.N_253\, Y => \I1.REG_28_sqmuxa\);
    
    \I1.REG_74_0_IV_0L271R_1952\ : AND2
      port map(A => \REGl271r\, B => 
        \I1.N_145_adt_net_854772__net_1\, Y => 
        \I1.REG_74l271r_adt_net_123732_\);
    
    \I2.MIC_REG2_i_0_il5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_314_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2_i_0_il5r_net_1\);
    
    \I2.LSRAM_INl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_413_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl29r_net_1\);
    
    \I2.FID_7_0_ivl28r\ : AO21
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl28r_net_1\, 
        C => \I2.FID_7l28r_adt_net_18747_\, Y => \I2.FID_7l28r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I38_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl17r\, B => 
        \I2.PIPE7_DTl17r_net_1\, Y => \I2.N282\);
    
    \I2.DTE_21_1_IV_0_0L4R_1334\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.DTE_2_1l4r_net_1\, C
         => \I2.DTE_21_1l4r_adt_net_39199_\, Y => 
        \I2.DTE_21_1l4r_adt_net_39210_\);
    
    \I2.PIPE4_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl15r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl15r_net_1\);
    
    \I2.FID_7_0_ivl13r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl13r_net_1\, 
        C => \I2.FID_7l13r_adt_net_18089_\, Y => \I2.FID_7l13r\);
    
    \I4.un1_lead_flag_1_3_0\ : MUX2L
      port map(A => \I4.N_2\, B => \I4.N_1\, S => 
        \I4.bcntl1r_net_1\, Y => \I4.N_3\);
    
    \I2.RAMAD_4_0l14r\ : MUX2H
      port map(A => \I2.RAMAD1l14r_net_1\, B => RAMAD_VMEl14r, S
         => \REG_i_il5r_adt_net_855552__net_1\, Y => \I2.N_541\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I177_Y\ : XOR2
      port map(A => \I2.N531_0\, B => 
        \I2.ADD_21x21_fast_I177_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l7r\);
    
    \I2.PLL_tdc_del.Core\ : PLLCORE
      port map(SDOUT => OPEN, SCLK => \GND\, SDIN => \GND\, 
        SSHIFT => \GND\, SUPDATE => \GND\, GLB => \I2.CLK_tdc\, 
        CLK => CLK_c, GLA => OPEN, CLKA => \GND\, LOCK => 
        \I2.PLL_LOCK_tdc\, MODE => \GND\, FBDIV5 => \GND\, EXTFB
         => \GND\, FBSEL0 => \VCC\, FBSEL1 => \GND\, FINDIV0 => 
        \GND\, FINDIV1 => \GND\, FINDIV2 => \GND\, FINDIV3 => 
        \GND\, FINDIV4 => \GND\, FBDIV0 => \GND\, FBDIV1 => \GND\, 
        FBDIV2 => \GND\, FBDIV3 => \GND\, FBDIV4 => \GND\, 
        STATBSEL => \GND\, DLYB0 => \GND\, DLYB1 => \GND\, OBDIV0
         => \GND\, OBDIV1 => \GND\, STATASEL => \GND\, DLYA0 => 
        \GND\, DLYA1 => \GND\, OADIV0 => \GND\, OADIV1 => \GND\, 
        OAMUX0 => \GND\, OAMUX1 => \GND\, OBMUX0 => \GND\, OBMUX1
         => \VCC\, OBMUX2 => \GND\, FBDLY0 => \VCC\, FBDLY1 => 
        \VCC\, FBDLY2 => \VCC\, FBDLY3 => \VCC\, XDLYSEL => \VCC\);
    
    DTE_padl31r : IOB33PH
      port map(PAD => DTE(31), A => \I2.DTE_1l31r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl31r);
    
    \I2.OFFSET_37_10l4r\ : MUX2L
      port map(A => \I2.N_703\, B => \I2.N_695\, S => 
        \I2.PIPE7_DTL26R_353\, Y => \I2.N_711\);
    
    \I3.PIPEA_240\ : MUX2L
      port map(A => \I3.PIPEAl9r_net_1\, B => 
        \I3.PIPEA_8l9r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854672__net_1\, Y
         => \I3.PIPEA_240_net_1\);
    
    \I1.NOELUTi_51\ : OAI21FTF
      port map(A => NOELUT_c, B => \I1.sstatel3r_net_1\, C => 
        \PULSEl0r_adt_net_854532__adt_net_855544__net_1\, Y => 
        \I1.NOELUTi_51_net_1\);
    
    \I3.VDBil8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_348_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil8r_net_1\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2527\ : OR3
      port map(A => \I3.N_2070_adt_net_163507_\, B => 
        \I3.N_2070_adt_net_163503_\, C => 
        \I3.N_2070_adt_net_163504_\, Y => 
        \I3.N_2070_adt_net_163510_\);
    
    TDCDA_padl15r : IB33
      port map(PAD => TDCDA(15), Y => TDCDA_cl15r);
    
    \I2.un78_pipe5_dt_2\ : XOR2
      port map(A => \I2.RAMDT4l11r_net_1\, B => 
        \I2.RAMDT4l10r_net_1\, Y => \I2.un78_pipe5_dt_2_net_1\);
    
    \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_1_1_net_1\, Y => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\);
    
    REGl200r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_101_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl200r\);
    
    \I5.SDAout_12_iv_0_o4_0\ : OAI21TTF
      port map(A => \I5.N_64\, B => \I5.COMMANDl1r_net_1\, C => 
        \I5.sstate1l11r_net_1\, Y => \I5.N_75\);
    
    REGl211r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_112_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl211r\);
    
    \I3.VDBi_31l10r\ : MUX2L
      port map(A => \I3.REGl143r\, B => \I3.VDBi_20l10r\, S => 
        \I3.REGMAPl17r_adt_net_854288__net_1\, Y => 
        \I3.VDBi_31l10r_net_1\);
    
    \I2.PIPE8_DT_546\ : MUX2L
      port map(A => \I2.PIPE8_DTl18r_net_1\, B => 
        \I2.PIPE8_DT_21l18r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_546_net_1\);
    
    \I1.REG_74_0_ivl165r\ : AO21
      port map(A => \REGl165r\, B => \I1.N_41\, C => 
        \I1.REG_74l165r_adt_net_133665_\, Y => \I1.REG_74l165r\);
    
    \I5.COMMANDl10r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_47_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl10r_net_1\);
    
    \I3.VDBoffa_50\ : OR3
      port map(A => \I3.VDBoffa_50_adt_net_163548_\, B => 
        \I3.N_2070_adt_net_163509_\, C => 
        \I3.N_2070_adt_net_163510_\, Y => \I3.VDBoffa_50_net_1\);
    
    \I2.un1_STATE1_24_0\ : AND2FT
      port map(A => \I2.STATE1l6r_net_1\, B => \I2.N_3887\, Y => 
        \I2.un1_STATE1_24\);
    
    \I2.NWPIPE2_1471\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE1_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE2_578\);
    
    \I5.SDAOUT_12_IV_0_920\ : AO21
      port map(A => \I5.N_75\, B => \I5.COMMANDl15r_net_1\, C => 
        \I5.SDAout_12_adt_net_9914_\, Y => 
        \I5.SDAout_12_adt_net_9915_\);
    
    \I2.TOKENTOB_RES\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.TOKENTOB_RES_649_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.TOKENTOB_RES_net_1\);
    
    \I2.DTO_16_1l10r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l10r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l10r_Rd1__net_1\);
    
    \I3.VDBI_31L1R_2700\ : OR3
      port map(A => \I3.VDBi_23l1r_adt_net_145542__net_1\, B => 
        \I3.VDBi_23l1r_adt_net_145528__net_1\, C => 
        \I3.VDBi_23l1r_adt_net_145541__net_1\, Y => 
        \I3.VDBi_31l1r_adt_net_506164_\);
    
    \I3.PIPEA_251\ : MUX2L
      port map(A => \I3.PIPEAl20r_net_1\, B => 
        \I3.PIPEA_8l20r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854660__net_1\, Y
         => \I3.PIPEA_251_net_1\);
    
    \I2.PIPE8_DT_533\ : MUX2L
      port map(A => \I2.PIPE8_DTl5r_net_1\, B => 
        \I2.PIPE8_DT_21l5r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_533_net_1\);
    
    \I3.VDBil6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_346_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil6r_net_1\);
    
    \I3.BLTCYC_113\ : MUX2H
      port map(A => \I3.BLTCYC_net_1\, B => 
        \I3.un7_cycs_0_a3_0_a3_net_1\, S => \I3.N_1508\, Y => 
        \I3.BLTCYC_113_net_1\);
    
    \I2.PIPE6_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_483_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl29r_net_1\);
    
    \I2.TDCGDBi\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TDCGDBi_673_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => TDCGDB_c);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I0_CO1_i_o2\ : AND2
      port map(A => \I2.RAMDT4L0R_770\, B => \I2.PIPE4_DTL0R_643\, 
        Y => \I2.N_85\);
    
    \I3.N_1935_adt_net_855332_\ : BFR
      port map(A => \I3.N_1935\, Y => 
        \I3.N_1935_adt_net_855332__net_1\);
    
    \I2.PIPE7_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl29r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl29r_net_1\);
    
    \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284_\ : BFR
      port map(A => \I3.un1_STATE2_7_1_adt_net_1473__net_1\, Y
         => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\);
    
    \I1.REG_74_i_o2_1_0_364_m4\ : NAND3
      port map(A => \I1.N_238_Rd1__adt_net_854888__net_1\, B => 
        \I1.PAGECNTl8r_net_1\, C => 
        \I1.REG_74_i_o2_1_0tt_364_m2_e_net_1\, Y => 
        \I1.REG_74_i_o2_1_0_364_N_5\);
    
    \I2.CRC32_12_0_0_m2l2r\ : MUX2L
      port map(A => \I2.DT_TEMPl2r_net_1\, B => \I2.N_4193\, S
         => \I2.N_4667_1_adt_net_1046__adt_net_854440__net_1\, Y
         => \I2.N_4187_i_i\);
    
    \I2.DTE_1l25r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l25r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l25r_Rd1__net_1\);
    
    \I3.VDBi_16_m_i_o3l3r_885\ : OR2
      port map(A => \I3.REGMAPL8R_741\, B => \I3.REGMAPl9r_net_1\, 
        Y => \I3.N_1907_263\);
    
    \I2.MIC_REG3_317\ : MUX2L
      port map(A => \I2.MIC_REG3l1r_net_1\, B => 
        \I2.MIC_REG3l0r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG3_317_net_1\);
    
    \I3.LWORDS_61\ : MUX2H
      port map(A => \I3.LWORDS_net_1\, B => LWORDB_in, S => 
        \I3.VSEL_0\, Y => \I3.LWORDS_61_net_1\);
    
    \I2.N_4538_i_i_o2\ : AND2
      port map(A => \I2.PIPE5_DTL23R_623\, B => 
        \I2.PIPE5_DTL21R_625\, Y => \I2.N_219\);
    
    \I3.RAMAD_VME_41\ : MUX2H
      port map(A => RAMAD_VMEl17r, B => \I3.REGl100r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_41_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL23R_1377\ : NOR2FT
      port map(A => REGl427r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, Y => 
        \I2.PIPE1_DT_42l23r_adt_net_46647_\);
    
    \I5.sstate1l8r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el5r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l8r_net_1\);
    
    \I3.un5_noemic_0_a2_i_o3_0_o3\ : AND2
      port map(A => \I3.SINGCYC_334\, B => \I3.WRITES_424\, Y => 
        \I3.N_277\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0\ : OR2FT
      port map(A => \I2.N_45_0\, B => \I2.N525_adt_net_57834_\, Y
         => \I2.N525\);
    
    TDCDB_padl8r : IB33
      port map(PAD => TDCDB(8), Y => TDCDB_cl8r);
    
    \I5.CHAIN_SELECT_11\ : MUX2H
      port map(A => \I5.CHAIN_SELECT_net_1\, B => 
        \I5.CHAIN_SELECT_4_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.CHAIN_SELECT_11_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I92_un1_Y\ : AND2
      port map(A => \I2.N338\, B => \I2.N331\, Y => 
        \I2.I92_un1_Y\);
    
    \I2.G_EVNT_NUM_n4_i_0_o2\ : NAND2
      port map(A => \I2.N_189_554\, B => \I2.G_EVNT_NUML4R_606\, 
        Y => \I2.N_4669\);
    
    \I1.REG_74_0_IVL244R_1982\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_10_sqmuxa_adt_net_854716__net_1\, Y => 
        \I1.REG_74l244r_adt_net_126383_\);
    
    \I1.REG_74_0_iv_0_0l260r\ : AO21
      port map(A => \REGl260r\, B => \I1.N_658\, C => 
        \I1.REG_74l260r_adt_net_124798_\, Y => \I1.REG_74l260r\);
    
    \I2.majority_reg_il4r\ : OAI21TTF
      port map(A => \I2.MIC_REG2_i_0_il4r_net_1\, B => 
        \I2.MIC_REG1l4r_net_1\, C => \I2.N_4424_adt_net_22594_\, 
        Y => \I2.N_4424\);
    
    TDCDA_padl16r : IB33
      port map(PAD => TDCDA(16), Y => TDCDA_cl16r);
    
    \I2.PIPE1_DT_42_1_IVL17R_1408\ : OAI21FTF
      port map(A => REGl437r, B => 
        \I2.N_3234_adt_net_855652__net_1\, C => 
        \I2.PIPE1_DT_42l17r_adt_net_47643_\, Y => 
        \I2.PIPE1_DT_42l17r_adt_net_47649_\);
    
    \I2.G_EVNT_NUM_923\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl11r_net_1\, B => 
        \I2.G_EVNT_NUM_n11\, S => \I2.N_3769\, Y => 
        \I2.G_EVNT_NUM_923_net_1\);
    
    \I2.un1_tdc_res_24_i_a3_0\ : NOR2
      port map(A => BNC_RES_c, B => TDC_RES_c_c, Y => 
        \I2.N_4680_0\);
    
    \I2.CRC32_12_i_0_x2l7r\ : XOR2FT
      port map(A => \I2.CRC32l7r_net_1\, B => \I2.N_226_i_i\, Y
         => \I2.N_250_i_i_0\);
    
    \I2.PIPE1_DT_42_1_IVL5R_1493\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl37r_net_1\, C => 
        \I2.PIPE1_DT_42l5r_adt_net_51167_\, Y => 
        \I2.PIPE1_DT_42l5r_adt_net_51185_\);
    
    \I3.VDBOFFA_31_IV_0L3R_2573\ : AO21
      port map(A => \REGl224r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.VDBoffa_31l3r_adt_net_164032_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164070_\);
    
    \I3.REG1l1r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG1_134_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l1r_net_1\);
    
    \I3.UN1_MYBERRI_1_SQMUXA_0_0_2347\ : AND2FT
      port map(A => \I3.ASBS_net_1\, B => \I3.PURGED_net_1\, Y
         => \I3.un1_MYBERRi_1_sqmuxa_adt_net_161483_\);
    
    \I2.EVNT_NUM_958\ : MUX2L
      port map(A => \I2.EVNT_NUMl5r_net_1\, B => 
        \I2.EVNT_NUM_n5_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_958_net_1\);
    
    \I2.TRGARRl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGARR_3l1r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGARRl1r_net_1\);
    
    \I2.END_TDC1_711\ : AO21FTF
      port map(A => \I2.N_3277\, B => \I2.END_TDC1_net_1\, C => 
        \I2.N_3281\, Y => \I2.END_TDC1_711_net_1\);
    
    \I5.COMMAND_13\ : MUX2H
      port map(A => \I5.COMMANDl1r_net_1\, B => 
        \I5.COMMAND_4l1r_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.COMMAND_13_net_1\);
    
    \I1.REG_74_0_IVL345R_1868\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l345r_adt_net_116584_\);
    
    \I3.REGMAP_I_0_IL19R_2987\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un76_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL19R_534\);
    
    \I2.CRC32_12_il8r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_117_i_i_0\, Y => 
        \I2.N_3925\);
    
    TOKOUTB_pad : IB33
      port map(PAD => TOKOUTB, Y => TOKOUTB_c);
    
    \I2.PIPE4_DTl11r_1148\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL11R_410\);
    
    \I1.REG_74_0_IV_0L363R_1844\ : AND2
      port map(A => \FBOUTl6r\, B => \I1.REG_25_sqmuxa\, Y => 
        \I1.REG_74l363r_adt_net_114611_\);
    
    \I3.REGMAPl10r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un44_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl10r_net_1\);
    
    \I2.PIPE8_DT_16_0l16r\ : MUX2H
      port map(A => \I2.PIPE8_DTl16r_net_1\, B => 
        \I2.PIPE7_DTl16r_net_1\, S => 
        \I2.N_565_0_adt_net_855736__net_1\, Y => \I2.N_582\);
    
    \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848_\ : BFR
      port map(A => \I2.MIC_REG1_1_sqmuxa_0\, Y => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I111_Y_1666\ : OA21FTF
      port map(A => \I2.N334\, B => \I2.N327\, C => \I2.N326\, Y
         => \I2.N445_i_adt_net_71447_\);
    
    \I2.ROFFSET_918\ : MUX2H
      port map(A => \I2.ROFFSETl0r_net_1\, B => 
        \I2.ROFFSET_n0_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_918_net_1\);
    
    LSRAM_FL_RADDRl0r : DFFC
      port map(CLK => CLK_c, D => \I4.LSRAM_FL_RADDR_9\, CLR => 
        CLEAR_STAT_i_0, Q => \LSRAM_FL_RADDRl0r\);
    
    \I3.REG_1_165\ : MUX2L
      port map(A => VDB_inl16r, B => REGl64r, S => 
        \I3.N_1935_adt_net_855324__net_1\, Y => \I3.REG_1_165_0\);
    
    ADE_padl13r : OB33PH
      port map(PAD => ADE(13), A => ADE_cl13r);
    
    \I2.SUB9_1_ADD_18X18_FAST_I36_Y_1655\ : AO21
      port map(A => \I2.N_3545_i_i\, B => \I2.G_1\, C => 
        \I2.N_3547_i_i\, Y => \I2.N301_1_adt_net_70232_\);
    
    \I3.PIPEB_107\ : MUX2H
      port map(A => \I3.PIPEBl28r_net_1\, B => 
        \I3.PIPEB_4l28r_net_1\, S => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_107_net_1\);
    
    \I2.PIPE7_DTL26R_2901\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_355\);
    
    \I2.un1_STATE2_9_0_0\ : OAI21TTF
      port map(A => \I2.N_176_i_adt_net_855708__net_1\, B => 
        \I2.N_4641\, C => \I2.STATE2l2r_adt_net_855212__net_1\, Y
         => \I2.un1_STATE2_9\);
    
    \I2.PIPE6_DT_476\ : MUX2H
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => 
        \I2.PIPE6_DTl22r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_476_net_1\);
    
    \I2.FCNT_946\ : MUX2L
      port map(A => \I2.FCNTl1r_net_1\, B => \I2.FCNT_n1_net_1\, 
        S => \I2.N_3267\, Y => \I2.FCNT_946_net_1\);
    
    \I3.REG_1l416r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_223_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl416r);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2387\ : AND2
      port map(A => \REGl290r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162136_\);
    
    \I2.L2TYPE_4_il14r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855716__net_1\, B => 
        \I2.N_4438_adt_net_66932_\, C => 
        \I2.N_4438_adt_net_66975_\, Y => \I2.N_4438\);
    
    \I2.G_EVNT_NUM_m_1_i_0_o2l8r_778\ : OR2FT
      port map(A => \I2.N_176_I_157\, B => \I2.N_4641_55\, Y => 
        \I2.N_223_156\);
    
    \I2.BNCID_VECTrff_11_254_0\ : AO21
      port map(A => \I2.BNCID_VECTwa15_1_net_1\, B => 
        \I2.BNCID_VECTrff_8_257_0_a2_0\, C => 
        \I2.BNCID_VECTro_11\, Y => 
        \I2.BNCID_VECTrff_11_254_0_net_1\);
    
    \I2.DTO_1l27r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l27r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l27r_Rd1__net_1\);
    
    \I1.BYTECNT_n4_i_o2\ : AND2
      port map(A => \I1.BYTECNT_i_0_il4r_net_1\, B => \I1.N_327\, 
        Y => \I1.N_334\);
    
    \I2.RAMAD1_661\ : MUX2L
      port map(A => \I2.RAMAD1_12l7r_net_1\, B => 
        \I2.RAMAD1l7r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__172\, Y => 
        \I2.RAMAD1_661_net_1\);
    
    \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Rd1__net_1\);
    
    \I2.SUB8_520_2727\ : OR3
      port map(A => \I2.SUB8_520_adt_net_635607_\, B => 
        \I2.SUB8_520_adt_net_635612_\, C => 
        \I2.SUB8_520_adt_net_635603_\, Y => \I2.SUB8_520_net_1\);
    
    \I2.FID_7_0_ivl20r\ : AO21
      port map(A => \I2.DTESl20r_net_1\, B => 
        \I2.STATE3l3r_net_1\, C => \I2.FID_7l20r_adt_net_17388_\, 
        Y => \I2.FID_7l20r\);
    
    \I1.REG_74_12_284_M10_I_0_0_1926\ : NOR2
      port map(A => \I1.PAGECNTl9r_net_1\, B => 
        \I1.REG_74_12_284_m10_i_o6_net_1\, Y => 
        \I1.REG_74_12_284_m10_i_0_i_adt_net_121593_\);
    
    \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392_\ : BFR
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854396__net_1\, 
        Y => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\);
    
    \I2.OFFSET_37_24l7r\ : MUX2L
      port map(A => \I2.N_818\, B => \I2.N_810\, S => 
        \I2.PIPE7_DTL26R_355\, Y => \I2.N_826\);
    
    \I2.PIPE10_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_622_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl17r_net_1\);
    
    \I2.RAMAD1_657\ : MUX2L
      port map(A => \I2.RAMAD1_12l3r_net_1\, B => 
        \I2.RAMAD1l3r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__173\, Y => 
        \I2.RAMAD1_657_net_1\);
    
    \I2.resyn_0_I2_un9_tdctrgi_0_a2\ : OR2FT
      port map(A => TDCTRG_C_570, B => \I2.STATE1l17r_net_1\, Y
         => \I2.un9_tdctrgi_i_0\);
    
    \I2.RAMDT4L12R_2815\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_143\);
    
    \I1.BYTECNT_N7_I_0_1782\ : XOR2
      port map(A => \I1.BYTECNTl7r_net_1\, B => \I1.N_358\, Y => 
        \I1.N_79_adt_net_109340_\);
    
    \I2.WPAGE_949\ : MUX2H
      port map(A => \I2.WPAGEl14r_net_1\, B => 
        \I2.WPAGE_n2_net_1\, S => 
        \I2.WPAGEe_adt_net_855056__net_1\, Y => 
        \I2.WPAGE_949_net_1\);
    
    \I3.VDBI_57_0_IVL23R_2159\ : AND2
      port map(A => \I3.PIPEAl23r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l23r_adt_net_138945_\);
    
    \I2.TDCDBSl29r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl29r, Q => 
        \I2.TDCDBSl29r_net_1\);
    
    \I2.N_2826_1_ADT_NET_794__2891\ : OAI21FTF
      port map(A => \I2.N_4261_304\, B => \I2.N_4282\, C => 
        \I2.N_2826_1_adt_net_40744__net_1\, Y => 
        \I2.N_2826_1_ADT_NET_794__332\);
    
    \I2.DTE_1l7r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l7r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l7r_Rd1__net_1\);
    
    \I1.REG_1_115\ : MUX2H
      port map(A => \REGl214r\, B => \I1.REG_74l214r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_115_net_1\);
    
    \I3.PIPEB_93_2330\ : NOR2FT
      port map(A => \I3.PIPEBl14r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_93_adt_net_160125_\);
    
    \I3.un64_reg_ads_0_a2_3_a3\ : NOR3
      port map(A => \I3.N_547\, B => \I3.N_554\, C => \I3.N_578\, 
        Y => \I3.un64_reg_ads_0_a2_3_a3_net_1\);
    
    \I3.N_90_i_0_a2_1\ : AND2
      port map(A => \I3.STATE1_IPL9R_717\, B => 
        \I3.REGMAPL0R_876\, Y => \I3.N_90_i_0_1\);
    
    \I4.bcnt_8\ : MUX2H
      port map(A => \I4.bcntl3r_net_1\, B => \I4.bcnt_3l3r_net_1\, 
        S => \I4.STATE1l1r_net_1\, Y => \I4.bcnt_8_net_1\);
    
    \I3.VADm_0_a3l9r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl9r_net_1\, Y => \I3.VADml9r\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I152_Y_0_1571\ : AO21
      port map(A => \I2.PIPE4_DTl17r_net_1\, B => 
        \I2.PIPE4_DTl18r_net_1\, C => \I2.RAMDT4L12R_797\, Y => 
        \I2.N498_0_adt_net_56939_\);
    
    \I5.REG_1_54\ : OAI21FTF
      port map(A => REGl117r, B => \I5.PULSE_I2C_net_1\, C => 
        \I5.REG_1_54_adt_net_11847_\, Y => \I5.REG_1_54_net_1\);
    
    \I5.REG_1l430r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_43_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl430r);
    
    \I2.OFFSET_37_20l4r\ : MUX2L
      port map(A => \I2.N_783\, B => \I2.N_775\, S => 
        \I2.PIPE7_DTL26R_358\, Y => \I2.N_791\);
    
    \I2.SUB8_523_2740\ : AND2FT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855156__net_1\, B
         => \I2.SUB8l20r_net_1\, Y => 
        \I2.SUB8_523_adt_net_670057_\);
    
    \I2.PIPE4_DTl14r_1533\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL14R_640\);
    
    \I3.PIPEA_8_0l25r\ : MUX2L
      port map(A => DPR_cl25r, B => \I3.PIPEA1l25r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855360__net_1\, Y => \I3.N_234\);
    
    \I1.REG_1_117\ : MUX2H
      port map(A => \REGl216r\, B => \I1.REG_74l216r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_117_net_1\);
    
    \I3.NOEAD_c_i_635\ : NOR2FT
      port map(A => \I3.MBLTCYC_net_1\, B => \I3.ADACKCYC_net_1\, 
        Y => NOEAD_C_I_0_13);
    
    \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_44987_\ : NOR2
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096__net_1\, B
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        Y => \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_44987__net_1\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855508_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__294\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\);
    
    \I2.REG_1l43r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n11_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl43r);
    
    \I2.CRC32_804\ : MUX2L
      port map(A => \I2.CRC32l9r_net_1\, B => \I2.N_3926\, S => 
        \I2.N_2826_1_ADT_NET_794__332\, Y => \I2.CRC32_804_net_1\);
    
    \I1.REG_74_0_IV_0_0L257R_1968\ : AND2
      port map(A => \FBOUTl4r\, B => \I1.N_596\, Y => 
        \I1.REG_74l257r_adt_net_125056_\);
    
    \I2.SUB8_1_sqmuxa_0_adt_net_855140_\ : BFR
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855152__net_1\, Y
         => \I2.SUB8_1_sqmuxa_0_adt_net_855140__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I28_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl7r\, B => \I2.PIPE7_DTL7R_698\, 
        Y => \I2.N252_0\);
    
    \I2.PIPE4_DTl2r_1252\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL2R_514\);
    
    \I2.PIPE1_DT_727\ : MUX2L
      port map(A => \I2.PIPE1_DTl0r_net_1\, B => 
        \I2.PIPE1_DT_42l0r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854588__net_1\, 
        Y => \I2.PIPE1_DT_727_net_1\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040_\ : BFR
      port map(A => \I2.PIPE1_DT_2_SQMUXA_ADT_NET_803__299\, Y
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040__net_1\);
    
    \I3.PIPEB_80_2343\ : NOR2FT
      port map(A => \I3.PIPEBl1r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_80_adt_net_160671_\);
    
    \I3.PIPEAl17r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_248_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl17r_net_1\);
    
    \I2.DTEST_FIFO\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTEST_FIFO_645_net_1\, CLR
         => CLEAR_STAT_i_0, Q => DTEST_FIFO);
    
    \I3.VDBi_57_0_iv_0l18r\ : OR2
      port map(A => \I3.VDBi_57l18r_adt_net_139494_\, B => 
        \I3.VDBi_57l18r_adt_net_139495_\, Y => \I3.VDBi_57l18r\);
    
    \I2.DTE_21_1_iv_2l2r\ : AO21
      port map(A => \I2.STATE2L3R_440\, B => \I2.DTO_9_ivl2r\, C
         => \I2.DTE_21_1_iv_2_il2r_adt_net_39453_\, Y => 
        \I2.DTE_21_1_iv_2_il2r\);
    
    \I2.REG_1_c10_i\ : OAI21FTF
      port map(A => \I2.un8_evread_1_adt_net_855784__net_1\, B
         => \I2.N_131\, C => \I2.N_3839_i_0_adt_net_101262_\, Y
         => \I2.N_3839_i_0\);
    
    \I3.PIPEBl15r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_94_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl15r_net_1\);
    
    \I2.SUB8_520_2725\ : AOI21TTF
      port map(A => \I2.N299_0\, B => \I2.N481_adt_net_88982_\, C
         => \I2.SUB8_520_adt_net_531407_\, Y => 
        \I2.SUB8_520_adt_net_635607_\);
    
    \I2.DTE_21_1l6r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l6r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l6r_Rd1__net_1\);
    
    \I3.TCNT_382\ : MUX2H
      port map(A => \I3.TCNTl2r_net_1\, B => \I3.TCNT_n2\, S => 
        \I3.TCNTe\, Y => \I3.TCNT_382_net_1\);
    
    \I4.LSRAM_FL_RD\ : DFFS
      port map(CLK => CLK_c, D => \I4.LSRAM_FL_RD_4_net_1\, SET
         => CLEAR_STAT_i_0, Q => LSRAM_FL_RD);
    
    \I2.FIDl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_434\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl18r);
    
    \I2.BNCID_VECTROR_1423\ : AOI21FTT
      port map(A => \I2.BNCID_VECTror_8_tz_0_i\, B => 
        \I2.BNCID_VECTror_8_tz_i_adt_net_48039_\, C => 
        \I2.TRGSERVL2R_582\, Y => 
        \I2.BNCID_VECTror_adt_net_48365_\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I140_Y_0_1549\ : AND2
      port map(A => \I2.N_59\, B => \I2.N_2360_tz_tz\, Y => 
        \I2.N519_adt_net_54631_\);
    
    \I2.ADEl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl6r);
    
    \I1.PAGECNT_327\ : MUX2H
      port map(A => \I1.PAGECNTl0r_adt_net_833884_Rd1__net_1\, B
         => \I1.PAGECNT_n0\, S => 
        \I1.PAGECNTe_adt_net_854896__net_1\, Y => 
        \I1.PAGECNT_327_net_1\);
    
    \I2.PIPE7_DTL27R_2792\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_85\);
    
    \I4.resyn_0_I4_LSRAM_FL_RADDR_0_sqmuxa\ : NAND2
      port map(A => \I4.N_48_3\, B => \I4.un1_lead_flag_1\, Y => 
        \I4.LSRAM_FL_RADDR_0_sqmuxa\);
    
    \I2.SUB8_522_2736\ : AOI21TTF
      port map(A => \I2.N477_adt_net_371248_\, B => 
        \I2.N477_adt_net_371301_\, C => 
        \I2.SUB8_522_adt_net_552099_\, Y => 
        \I2.SUB8_522_adt_net_659164_\);
    
    \I5.DATA_12l15r\ : MUX2H
      port map(A => \I5.SBYTEl7r_net_1\, B => REGl132r, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l15r_net_1\);
    
    \I3.VDBoffa_31_iv_0l4r\ : AND2
      port map(A => \REGl177r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        Y => \I3.VDBoffa_31l4r_adt_net_163834_\);
    
    \I2.TRGCNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGCNT_n0_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGCNTl0r_net_1\);
    
    \I5.AIR_WDATAl2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_57_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl2r_net_1\);
    
    \I1.REG_74_0_iv_0_0_a2l253r\ : AND2FT
      port map(A => \I1.N_1169_adt_net_854820__net_1\, B => 
        \I1.N_596_adt_net_124704_\, Y => \I1.N_596\);
    
    \I2.DTE_1_857\ : MUX2L
      port map(A => \I2.DTE_1l19r_Rd1__net_1\, B => 
        \I2.DTE_21_1l19r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\, Y => 
        \I2.DTE_1l19r\);
    
    \I2.un2_evnt_word_I_37\ : AND2
      port map(A => \I2.WOFFSETl6r\, B => \I2.N_34\, Y => 
        \I2.N_29\);
    
    \I2.MIC_ERR_REGSl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_349_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl20r_net_1\);
    
    \I2.CRC32l25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_820_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l25r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL4R_1500\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855224__net_1\, B => 
        \I2.MIC_ERR_REGSl4r_net_1\, C => 
        \I2.PIPE1_DT_42l4r_adt_net_51432_\, Y => 
        \I2.PIPE1_DT_42l4r_adt_net_51433_\);
    
    \I1.REG_74_0_IVL188R_2046\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l188r_adt_net_131613_\);
    
    \I3.REGMAP_I_0_IL38R_2801\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un171_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL38R_113\);
    
    \I2.MIC_REG2_310\ : MUX2H
      port map(A => \I2.MIC_REG2l1r_net_1\, B => 
        \I2.MIC_REG2l2r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG2_310_net_1\);
    
    \I5.COMMAND_4l10r\ : MUX2L
      port map(A => \I5.AIR_WDATAl10r_net_1\, B => REGl111r, S
         => REGl7r, Y => \I5.COMMAND_4l10r_net_1\);
    
    \I2.REG_1l36r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl36r);
    
    \I2.MIC_REG3_318\ : MUX2H
      port map(A => \I2.MIC_REG3l1r_net_1\, B => 
        \I2.MIC_REG3l2r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG3_318_net_1\);
    
    \I2.PIPE1_DT_42_I_0L15R_1428\ : OAI21FTT
      port map(A => \I2.N_3876_adt_net_855252__net_1\, B => 
        \I2.STATE1L18R_628\, C => \I2.N_3888\, Y => 
        \I2.N_3238_adt_net_48555_\);
    
    \I3.VDBoffb_30_iv_0l0r\ : AND2
      port map(A => \REGl365r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163074_\);
    
    DTE_padl15r : IOB33PH
      port map(PAD => DTE(15), A => \I2.DTE_1l15r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl15r);
    
    \I3.TCNT1_n3\ : XOR2
      port map(A => \I3.TCNT1_i_0_il3r_net_1\, B => 
        \I3.TCNT1_c2_net_1\, Y => \I3.TCNT1_n3_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I64_Y\ : AO21
      port map(A => \I2.N255_0\, B => 
        \I2.N316_i_i_adt_net_86577_\, C => 
        \I2.N312_0_adt_net_86450_\, Y => \I2.N314\);
    
    \I3.REG2_228\ : OAI21FTF
      port map(A => \I3.REG2l405r_net_1\, B => \I3.N_1563\, C => 
        \I3.REG2_15l405r\, Y => \I3.REG2_228_net_1\);
    
    \I2.resyn_0_I2_BITCNT_n4_i\ : NOR3
      port map(A => \I2.ERR_WORDS_RDY_0_sqmuxa\, B => \I2.N_4337\, 
        C => \I2.N_4330\, Y => \I2.N_4325\);
    
    \I3.REGMAPL27R_2986\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un116_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAPL27R_533\);
    
    \I3.VDBi_16l8r\ : MUX2L
      port map(A => REGl40r, B => \I3.VDBi_10l8r_net_1\, S => 
        \I3.REGMAPl7r_net_1\, Y => \I3.VDBi_16l8r_net_1\);
    
    \I2.BNCID_VECTrff_4\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_4_261_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_4\);
    
    \I2.END_EVNT5_1144_1733\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT5_840\);
    
    TDCDA_padl21r : IB33
      port map(PAD => TDCDA(21), Y => TDCDA_cl21r);
    
    \I1.SSTATEL7R_3000\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.sstate_ns_0_iv_0_il3r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL7R_754\);
    
    \I2.REG_1_C1_I_1745\ : NOR2
      port map(A => REGl33r, B => \I2.N_121\, Y => 
        \I2.N_3830_adt_net_101622_\);
    
    \I2.PIPE10_DT_17_0L29R_1614\ : AND2
      port map(A => \I2.N_22_i_0_adt_net_855596__net_1\, B => 
        \I2.N_3822\, Y => \I2.PIPE10_DT_17l29r_adt_net_64809_\);
    
    \I2.TRGSERVl3r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l3r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVl3r_net_1\);
    
    DPR_padl9r : IB33
      port map(PAD => DPR(9), Y => DPR_cl9r);
    
    VAD_padl2r : IOB33PH
      port map(PAD => VAD(2), A => \I3.VADml2r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl2r);
    
    \I2.un1_STATE1_28_0\ : AOI21FTT
      port map(A => \I2.CHAINA_EN244_i_adt_net_855260__net_1\, B
         => \I2.N_148\, C => \I2.STATE1l13r_net_1\, Y => 
        \I2.un1_STATE1_28\);
    
    \I2.resyn_0_I2_BITCNT_n1_i_o3\ : AND2
      port map(A => \I2.BITCNT_c0\, B => \I2.BITCNTl1r_net_1\, Y
         => \I2.N_4327\);
    
    \I3.VDBi_40_0_i_m2l2r\ : MUX2L
      port map(A => REGl420r, B => REGl436r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_134\);
    
    \I2.ADOl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl9r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0_o2_1_725\ : OR2
      port map(A => \I2.N_128_0\, B => 
        \I2.N_74_ADT_NET_55281__325\, Y => \I2.N_74_103\);
    
    \I2.OFFSET_37_7l6r\ : MUX2L
      port map(A => \I2.N_681\, B => \I2.N_657\, S => 
        \I2.PIPE7_DTL25R_682\, Y => \I2.N_689\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I15_G0N_i_o4\ : NAND2
      port map(A => \I2.RAMDT4L12R_799\, B => 
        \I2.PIPE4_DTl15r_net_1\, Y => \I2.N_8_0\);
    
    \I2.SUB8_504\ : MUX2H
      port map(A => \I2.SUB8l1r_net_1\, B => \I2.SUB8_2l1r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855136__net_1\, Y => 
        \I2.SUB8_504_net_1\);
    
    \I3.REGMAPL9R_3030\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un41_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL9R_784\);
    
    REGl280r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_181_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl280r\);
    
    \I1.REG_1_113\ : MUX2H
      port map(A => \REGl212r\, B => \I1.N_1350\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_113_net_1\);
    
    CHAINA_EN244_pad : OB33PH
      port map(PAD => CHAINA_EN244, A => 
        \I2.CHAINA_EN244_i_adt_net_855264__net_1\);
    
    \I2.N_2828_ADT_NET_1062__ADT_NET_835312_RD1__2910\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2828_adt_net_1062__net_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.N_2828_ADT_NET_1062__ADT_NET_835312_RD1__379\);
    
    \I2.DTO_16_1_IV_0L27R_1078\ : AND2
      port map(A => \I2.DT_TEMPl27r_net_1\, B => 
        \I2.N_4671_adt_net_854600__net_1\, Y => 
        \I2.DTO_16_1l27r_adt_net_29240_\);
    
    \I2.RAMDT4L5R_3055\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_809\);
    
    \I1.REG_74_0_IVL167R_2067\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l167r_adt_net_133493_\);
    
    \I4.resyn_0_I4_LSRAM_FL_RADDR_0_sqmuxa_1\ : NOR2FT
      port map(A => \I4.STATE1l1r_net_1\, B => 
        \I4.LSRAM_FL_RADDR_0_sqmuxa\, Y => 
        \I4.LSRAM_FL_RADDR_0_sqmuxa_1\);
    
    \I3.VDBi_13l4r\ : AND3FFT
      port map(A => \I2.N_3877_adt_net_4723_\, B => 
        \I2.N_3877_adt_net_4725_\, C => \I3.REGMAPl2r_net_1\, Y
         => \I3.VDBi_13l4r_adt_net_284333_\);
    
    \I3.N_1413_i_i_o3\ : OR2
      port map(A => \I3.STATE1_ipl0r_net_1\, B => 
        \I3.STATE1_ipl3r_net_1\, Y => \I3.N_1764\);
    
    \I2.REG_1l37r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n5_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl37r);
    
    \I2.N_2864_0_adt_net_854264_\ : BFR
      port map(A => \I2.N_2864_0\, Y => 
        \I2.N_2864_0_adt_net_854264__net_1\);
    
    \I3.REG_1_292\ : MUX2L
      port map(A => VDB_inl10r, B => REGl111r, S => 
        \I3.N_318_adt_net_855888__net_1\, Y => \I3.REG_1_292_0\);
    
    \I2.N_152_i_adt_net_4109_\ : OR2
      port map(A => \I2.N_75\, B => 
        \I2.N_152_i_adt_net_54710__net_1\, Y => 
        \I2.N_152_i_adt_net_4109__net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I179_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl9r_net_1\, Y => \I2.ADD_21x21_fast_I179_Y_0\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I179_Y_2687\ : AO21FTT
      port map(A => \I2.N303_0\, B => \I2.N349\, C => 
        \I2.N481_adt_net_424213_\, Y => \I2.N481_adt_net_424221_\);
    
    \I3.RAMAD_VME_34\ : MUX2H
      port map(A => RAMAD_VMEl10r, B => \I3.REGl93r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_34_net_1\);
    
    \I3.PULSE_330_adt_net_854736_\ : BFR
      port map(A => \I3.PULSE_330_net_1\, Y => 
        \I3.PULSE_330_adt_net_854736__net_1\);
    
    \I1.REG_74_3L404R_1838\ : AO21
      port map(A => \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__363\, B
         => \I1.N_253\, C => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854396__net_1\, 
        Y => \I1.N_273_10_adt_net_114360_\);
    
    \I3.REGMAPl9r_adt_net_854316_\ : BFR
      port map(A => \I3.REGMAPl9r_adt_net_854320__net_1\, Y => 
        \I3.REGMAPl9r_adt_net_854316__net_1\);
    
    \I2.PIPE6_DT_456\ : MUX2H
      port map(A => \I2.PIPE5_DTl2r_net_1\, B => 
        \I2.PIPE6_DTl2r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_456_net_1\);
    
    \I3.VDBOFFB_30_IV_0L2R_2452\ : AO21
      port map(A => \REGl391r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l2r_adt_net_162738_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162745_\);
    
    \I3.PIPEA1_12l28r\ : NAND2FT
      port map(A => DPR_cl28r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, Y => 
        \I3.PIPEA1_12l28r_net_1\);
    
    \I2.BNCID_VECTrff_9_256_0_a2_0\ : NOR3FFT
      port map(A => TDCTRG_c, B => \I2.TRGARRl3r_net_1\, C => 
        \I2.TRGARRl2r_net_1\, Y => 
        \I2.BNCID_VECTrff_8_257_0_a2_0\);
    
    \I3.PIPEB_88\ : AO21
      port map(A => DPR_cl9r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_88_adt_net_160335_\, Y => 
        \I3.PIPEB_88_net_1\);
    
    \I2.NWRSRAMO\ : OR2
      port map(A => \I2.CLK_sram\, B => \I2.WROi_net_1\, Y => 
        NWRSRAMO_c);
    
    \I5.TEMPDATA_75\ : MUX2L
      port map(A => \I5.TEMPDATAl1r_net_1\, B => REGl126r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_75_net_1\);
    
    \I3.VAS_76\ : MUX2L
      port map(A => VAD_inl14r, B => \I3.VAS_i_0_il14r\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_76_net_1\);
    
    \I3.REG_44_i_a2_0l88r\ : NOR2
      port map(A => VDB_inl5r, B => \I3.N_98\, Y => \I3.N_1671\);
    
    \I2.FID_7_0_IVL6R_1721\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl54r, C => 
        \I2.FID_7l6r_adt_net_92927_\, Y => 
        \I2.FID_7l6r_adt_net_92935_\);
    
    \I2.ROFFSETl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_916_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl2r_net_1\);
    
    \I2.RAMAD1l16r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_670_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l16r_net_1\);
    
    \I2.OFFSETl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_564_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl4r_net_1\);
    
    \I1.REG_1_140\ : MUX2H
      port map(A => \REGl239r\, B => \I1.REG_74l239r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\, Y => 
        \I1.REG_1_140_net_1\);
    
    \I2.TDCDBSl21r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl21r, Q => 
        \I2.TDCDBSl21r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2610\ : AO21
      port map(A => \REGl174r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        C => \I3.VDBoffa_31l1r_adt_net_164416_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164451_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I184_Y\ : XOR2FT
      port map(A => \I2.N_40\, B => \I2.ADD_21x21_fast_I184_Y_0\, 
        Y => \I2.un27_pipe5_dt0l14r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_1_1\ : 
        NAND3FFT
      port map(A => \I2.N_107_adt_net_276024_\, B => 
        \I2.N_107_adt_net_256840_\, C => \I2.N_17\, Y => 
        \I2.N_108\);
    
    \I3.STATE2_NS_I_I_A5_0_A3L1R_2115\ : NOR3FTT
      port map(A => EVRDY_c, B => \I3.EFS_net_1\, C => \I3.N_258\, 
        Y => \I3.STATE2_ns_i_i_a5_0_a3l1r_adt_net_135757_\);
    
    \I3.TCNT3l3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT3_376_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT3l3r_net_1\);
    
    \I1.REG_74_0_IVL267R_1956\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, Y => 
        \I1.REG_74l267r_adt_net_124113_\);
    
    \I1.SBYTE_8_0_a2_il0r\ : AND2
      port map(A => \I1.N_371_i\, B => \I1.N_405\, Y => 
        \I1.N_186\);
    
    \I1.REG_1_300\ : MUX2H
      port map(A => \REGl399r\, B => \I1.REG_74l399r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\, Y => 
        \I1.REG_1_300_net_1\);
    
    \I3.VDBil7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_347_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil7r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I151_Y_i_1\ : NAND3
      port map(A => \I2.N_41\, B => \I2.N_63\, C => \I2.N_33\, Y
         => \I2.N_1_1\);
    
    \I2.PIPE7_DTL26R_2900\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_354\);
    
    \I2.PIPE1_DT_42_1_IVL11R_1457\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl43r_net_1\, C => 
        \I2.PIPE1_DT_42l11r_adt_net_49685_\, Y => 
        \I2.PIPE1_DT_42l11r_adt_net_49703_\);
    
    \I1.REG_1_116\ : MUX2H
      port map(A => \REGl215r\, B => \I1.REG_74l215r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_116_net_1\);
    
    \I5.TEMPDATAl1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_75_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl1r_net_1\);
    
    \I1.REG_74_8_0_o4_a0_0l324r_723\ : OR2
      port map(A => \I1.PAGECNTL5R_309\, B => \I1.PAGECNTL6R_249\, 
        Y => \I1.REG_74_1_A0_0L228R_101\);
    
    \I2.PIPE7_DTl25r_1575\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL25R_682\);
    
    \I1.REG_74_0_ivl388r\ : AO21
      port map(A => \REGl388r\, B => \I1.N_257\, C => 
        \I1.REG_74l388r_adt_net_111319_\, Y => 
        \I1.REG_74l388r_net_1\);
    
    \I1.REG_17_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_260\, B => \I1.N_242\, Y => 
        \I1.REG_17_sqmuxa\);
    
    \I2.DT_SRAM_i_m2l24r\ : MUX2L
      port map(A => \I2.N_4192\, B => \I2.PIPE2_DTl24r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668__net_1\, 
        Y => \I2.N_4194\);
    
    \I2.G_EVNT_NUM_926\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl8r_net_1\, B => \I2.N_4640\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_926_net_1\);
    
    \I2.TDCDBSl5r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl5r, Q => 
        \I2.TDCDBSl5r_net_1\);
    
    \I2.CHAINB_ERRS\ : DFFC
      port map(CLK => CLK_c, D => \I2.CHAINB_ERRS_525_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.CHAINB_ERRS_net_1\);
    
    \I3.VDBOFFB_30_IV_0L4R_2407\ : AND2
      port map(A => \REGl345r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        Y => \I3.VDBoffb_30l4r_adt_net_162334_\);
    
    \I2.OFFSET_37_14l1r\ : MUX2L
      port map(A => \I2.N_732\, B => \I2.N_684\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_740\);
    
    \I2.CRC32_12_0_0_x2l21r\ : XOR2FT
      port map(A => \I2.CRC32l21r_net_1\, B => \I2.N_4039_i_i\, Y
         => \I2.N_58_i_0_i_0\);
    
    \I3.VDBi_31l28r\ : MUX2L
      port map(A => \I3.REGl161r\, B => \I3.VDBi_20l28r\, S => 
        \I3.REGMAPl17r_adt_net_854284__net_1\, Y => 
        \I3.VDBi_31l28r_net_1\);
    
    \I2.ROFFSET_n5\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855700__net_1\, B => 
        \I2.ROFFSET_n5_tz_i\, Y => \I2.ROFFSET_n5_net_1\);
    
    \I3.VDBi_57_iv_0_0l2r\ : OR3
      port map(A => \I3.VDBi_57l2r_adt_net_145372_\, B => 
        \I3.VDBi_57l2r_adt_net_145380_\, C => 
        \I3.VDBi_57l2r_adt_net_145381_\, Y => \I3.VDBi_57l2r\);
    
    \I2.BNC_IDl2r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_9_1\, CLR => 
        \I2.N_4622_i_0\, SET => \I2.N_4610_i_0\, Q => 
        \I2.BNC_IDl2r_net_1\);
    
    \I2.RAMAD1_658\ : MUX2L
      port map(A => \I2.RAMAD1_12l4r_net_1\, B => 
        \I2.RAMAD1l4r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__173\, Y => 
        \I2.RAMAD1_658_net_1\);
    
    \I3.REGMAPl23r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un96_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl23r_net_1\);
    
    \I2.DTO_9_ivl11r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl11r_net_1\, 
        C => \I2.DTO_9l11r_adt_net_32812_\, Y => \I2.DTO_9l11r\);
    
    \I3.VDBml17r\ : MUX2L
      port map(A => \I3.VDBil17r_net_1\, B => \I3.N_159\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml17r_net_1\);
    
    \I3.VDBI_20_IVL12R_2203\ : AND2
      port map(A => REGl60r, B => 
        \I3.REGMAPl9r_adt_net_854308__net_1\, Y => 
        \I3.VDBi_20l12r_adt_net_140765_\);
    
    \I3.REGMAPl8r_1634\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un37_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL8R_741\);
    
    \I2.RAMAD_4_0l2r\ : MUX2H
      port map(A => \I2.RAMAD1l2r_net_1\, B => RAMAD_VMEl2r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_529\);
    
    \I1.sstatel3r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl7r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel3r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL2R_1510\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl34r_net_1\, C => 
        \I2.PIPE1_DT_42l2r_adt_net_51819_\, Y => 
        \I2.PIPE1_DT_42l2r_adt_net_51836_\);
    
    \I2.CRC32_814\ : MUX2L
      port map(A => \I2.CRC32l19r_net_1\, B => \I2.N_3936\, S => 
        \I2.N_2826_1_ADT_NET_794__330\, Y => \I2.CRC32_814_net_1\);
    
    \I2.PIPE1_DTl10r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_737_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl10r_net_1\);
    
    \I1.REG_74_0_IVL347R_1866\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l347r_adt_net_116412_\);
    
    \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834764_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_0_sqmuxa_i_0_N_3_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834764_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2553\ : AO21
      port map(A => \REGl201r\, B => \I3.REGMAPl22r_net_1\, C => 
        \I3.VDBoffa_31l4r_adt_net_163834_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163878_\);
    
    \I2.TDCDBSl2r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl2r, Q => 
        \I2.TDCDBSl2r_net_1\);
    
    \I1.REG_74_0_iv_i_a2l211r\ : AO21
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, C => 
        \I1.N_144_adt_net_129587_\, Y => \I1.N_144\);
    
    \I3.REGMAPl2r_1629\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un13_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL2R_736\);
    
    \I1.REG_5_sqmuxa_0_a2_0\ : OR3FTT
      port map(A => \I1.PAGECNTL7R_525\, B => \I1.PAGECNTL8R_457\, 
        C => \I1.N_1169_168\, Y => \I1.N_243\);
    
    \I2.RAMDT4L4R_3097\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl4r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L4R_883\);
    
    \I2.TDCDASl24r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl24r, Q => 
        \I2.TDCDASl24r_net_1\);
    
    \I1.REG_74_0_iv_0l367r\ : AO21
      port map(A => \REGl367r\, B => \I1.N_660\, C => 
        \I1.REG_74l367r_adt_net_113740_\, Y => \I1.REG_74l367r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I34_P0N_1282\ : OR2FT
      port map(A => \I2.LSRAM_OUTl13r_adt_net_854940__net_1\, B
         => \I2.PIPE7_DTl13r_net_1\, Y => \I2.N270_0_544\);
    
    \I2.DTO_16_1_IVL22R_1106\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855676__net_1\, B => 
        \I2.DTO_9l22r\, Y => \I2.DTO_16_1l22r_adt_net_30346_\);
    
    \I2.N_4547_1_adt_net_1209__adt_net_855616_\ : BFR
      port map(A => \I2.N_4547_1_adt_net_1209__net_1\, Y => 
        \I2.N_4547_1_adt_net_1209__adt_net_855616__net_1\);
    
    \I2.PIPE8_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_541_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl13r_net_1\);
    
    \I2.OFFSET_37_17l3r\ : MUX2L
      port map(A => \I2.N_758\, B => \I2.N_750\, S => 
        \I2.PIPE7_DTL26R_354\, Y => \I2.N_766\);
    
    \I2.N_2868_1_adt_net_836000_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2868_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\);
    
    \I3.TCNT_n0_0_0\ : OAI21
      port map(A => \I3.TCNTl0r_net_1\, B => 
        \I3.un1_STATE1_10_i_0\, C => \I3.N_1966_1\, Y => 
        \I3.TCNT_n0\);
    
    \I2.N_3883_adt_net_854632_\ : BFR
      port map(A => \I2.N_3883\, Y => 
        \I2.N_3883_adt_net_854632__net_1\);
    
    \I2.N_152_i_adt_net_54710_\ : OA21
      port map(A => \I2.PIPE4_DTL17R_636\, B => 
        \I2.PIPE4_DTL15R_637\, C => \I2.RAMDT4L5R_816\, Y => 
        \I2.N_152_i_adt_net_54710__net_1\);
    
    ADE_padl9r : OB33PH
      port map(PAD => ADE(9), A => ADE_cl9r);
    
    \I2.DTO_16_1_iv_1l1r\ : AO21FTT
      port map(A => \I2.DTO_1l1r_net_1\, B => \I2.N_196_53\, C
         => \I2.DTO_16_1_iv_1l1r_adt_net_35128_\, Y => 
        \I2.DTO_16_1_iv_1l1r_net_1\);
    
    \I2.PIPE4_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl10r_net_1\);
    
    \I3.N_1935_adt_net_855328_\ : BFR
      port map(A => \I3.N_1935\, Y => 
        \I3.N_1935_adt_net_855328__net_1\);
    
    \I2.EVRDYi\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVRDYi_496_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => EVRDY_c);
    
    \I2.DT_TEMPl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_792_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl31r_net_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I108_Y_1658\ : OAI21FTF
      port map(A => \I2.N460\, B => \I2.N329\, C => \I2.N328\, Y
         => \I2.N436_adt_net_70670_\);
    
    \I2.DTE_cl_0_sqmuxa_2_0_a2_0_a2_0_912\ : OR2FT
      port map(A => \I2.N_4241_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, Y => 
        \I2.DTE_CL_0_SQMUXA_2_0_290\);
    
    \I2.WOFFSET_827\ : MUX2L
      port map(A => 
        \I2.WOFFSETl0r_adt_net_854636__adt_net_855712__net_1\, B
         => \I2.WOFFSET_13l0r\, S => 
        \I2.N_2828_adt_net_1062__net_1\, Y => 
        \I2.WOFFSET_827_net_1\);
    
    \I2.CRC32_12_i_0l31r\ : NOR2
      port map(A => \I2.N_2867_1_adt_net_854964__net_1\, B => 
        \I2.N_244_i_i_0\, Y => \I2.N_3948\);
    
    \I3.RAMAD_VME_38\ : MUX2H
      port map(A => RAMAD_VMEl14r, B => \I3.REGl97r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_38_net_1\);
    
    \I2.DT_SRAM_0l26r\ : MUX2L
      port map(A => \I2.PIPE10_DTl26r_net_1\, B => 
        \I2.PIPE5_DTl26r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854220__net_1\, Y => 
        \I2.N_894\);
    
    \I3.REG_1l90r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_271_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl90r);
    
    \I3.STATE1_NS_0_IV_0_0L7R_2120\ : NOR2FT
      port map(A => 
        \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344__net_1\, 
        B => \I3.N_57_i_0_0_adt_net_854692__net_1\, Y => 
        \I3.STATE1_nsl7r_adt_net_136170_\);
    
    \I2.un2_evnt_word_I_5\ : XOR2
      port map(A => 
        \I2.WOFFSETl0r_adt_net_854636__adt_net_855712__net_1\, B
         => \I2.WOFFSETl1r_adt_net_854992__net_1\, Y => 
        \I2.I_5_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I185_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L5R_139\, B => 
        \I2.PIPE4_DTl15r_net_1\, Y => 
        \I2.ADD_21x21_fast_I185_Y_0\);
    
    \I3.REG_44_IL86R_2305\ : AOI21FTT
      port map(A => REGl86r, B => \I3.N_98_0\, C => \I3.N_1667\, 
        Y => \I3.N_1632_adt_net_150363_\);
    
    \I2.FIFO_END_EVNT_489\ : OAI21FTF
      port map(A => \I2.FIFO_END_EVNT_net_1\, B => 
        \I2.STATE3l5r_net_1\, C => 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\, Y => 
        \I2.FIFO_END_EVNT_489_net_1\);
    
    \I2.PIPE8_DT_534\ : MUX2L
      port map(A => \I2.PIPE8_DTl6r_net_1\, B => 
        \I2.PIPE8_DT_21l6r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_534_net_1\);
    
    \I2.STATE1l8r_1541\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3234_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1L8R_648\);
    
    \I2.G_EVNT_NUMl1r_928\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_933_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUML1R_306\);
    
    \I1.REG_1_165\ : MUX2H
      port map(A => \REGl264r\, B => \I1.REG_74l264r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y => 
        \I1.REG_1_165_net_1\);
    
    \I3.REG_0_sqmuxa_2_0_a2_0_a3\ : AND2
      port map(A => \I3.REGMAPl17r_adt_net_854296__net_1\, B => 
        \I3.N_1906_i_0_0_adt_net_855640__net_1\, Y => 
        \I3.REG_0_sqmuxa_2\);
    
    \I5.sstate1l4r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el9r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l4r_net_1\);
    
    \I5.REG_1_24\ : MUX2H
      port map(A => \I5.TEMPDATAl5r_net_1\, B => REGl441r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_24_net_1\);
    
    \I1.REG_16_sqmuxa_0_a2_0_720\ : OR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835132_RD1__884\, B
         => \I1.REG_74_1_A0_0L228R_102\, Y => \I1.N_253_98\);
    
    \I3.REG_1_180\ : MUX2L
      port map(A => VDB_inl31r, B => REGl79r, S => 
        \I3.N_1935_adt_net_855316__net_1\, Y => \I3.REG_1_180_0\);
    
    \I1.REG_74_12_300_N_15_adt_net_3731_\ : NAND2
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720__adt_net_835724_Rd1__net_1\, 
        B => \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__361\, Y => 
        \I1.REG_74_12_300_N_15_adt_net_3731__net_1\);
    
    \I2.REG_1l42r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n10_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REG_i_0_il42r);
    
    \I2.LEAD_FLAG6_637_1606\ : NOR2FT
      port map(A => LEAD_FLAGl0r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_637_adt_net_64628_\);
    
    \I2.un19_start_giro_i_0_o2\ : NOR2
      port map(A => \I2.FIFO_END_EVNT_net_1\, B => 
        \I2.EVNT_REJ_net_1\, Y => \I2.N_3850\);
    
    \I1.REG_74_0_iv_0l269r\ : AO21
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, C => 
        \I1.REG_74l269r_adt_net_123904_\, Y => \I1.REG_74l269r\);
    
    \I3.N_57_i_0_a3_0\ : NOR2
      port map(A => \I3.N_1919\, B => \I3.TCNTl4r_net_1\, Y => 
        \I3.N_57_i_0_0\);
    
    \I2.MIC_REG1L3R_ADT_NET_834596_RD1__2912\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_304_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1L3R_ADT_NET_834596_RD1__381\);
    
    \I3.REG_1_200\ : MUX2L
      port map(A => VDB_inl19r, B => \I3.REGl152r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\, Y => 
        \I3.REG_1_200_0\);
    
    \I2.EVNT_NUM_i_ml8r\ : NOR2
      port map(A => \I2.PIPE1_DT_42_3_0L28R_339\, B => 
        \I2.EVNT_NUMl8r_net_1\, Y => \I2.EVNT_NUM_i_m_il8r\);
    
    \I2.DTE_21_1_IV_0_0L7R_1315\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855120__net_1\, B => 
        \I2.EVNT_WORDl3r_net_1\, Y => 
        \I2.DTE_21_1l7r_adt_net_38855_\);
    
    \I2.un1_STATE3_10_1_adt_net_999_\ : OR3
      port map(A => \I2.STATE3L2R_413\, B => \I2.STATE3l9r_net_1\, 
        C => \I2.un1_STATE3_10_1_adt_net_17431__net_1\, Y => 
        \I2.un1_STATE3_10_1_adt_net_999__net_1\);
    
    \I3.VADm_0_a3l10r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl10r_net_1\, Y => \I3.VADml10r\);
    
    \I2.NWPIPE8_0\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, 
        SET => CLEAR_STAT_i_0, Q => \I2.NWPIPE8_I_0_I_0_0_6\);
    
    \I2.STATEe_illegalpipe2\ : DFFLC
      port map(CLK => CLK_c, D => \I2.STATEe_illegalpipe1_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.STATEe_illegalpipe2_net_1\);
    
    \I1.REG_1_167\ : MUX2H
      port map(A => \REGl266r\, B => \I1.REG_74l266r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y => 
        \I1.REG_1_167_net_1\);
    
    \I1.REG_1_148\ : MUX2H
      port map(A => \REGl247r\, B => \I1.REG_74l247r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_148_net_1\);
    
    \I3.VDBi_16_m_i_a2l11r\ : OR2
      port map(A => \I3.REGMAPL2R_736\, B => \I3.REGMAPL7R_459\, 
        Y => \I3.N_2018\);
    
    \I3.VDBi_371\ : MUX2L
      port map(A => \I3.VDBil31r_net_1\, B => \I3.VDBi_57l31r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_371_net_1\);
    
    \I2.LEAD_FLAG6_1_sqmuxa_i\ : OR2
      port map(A => END_FLUSH_560, B => 
        \I2.N_4527_adt_net_63801_\, Y => \I2.N_4527\);
    
    \I2.OFFSETl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_567_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl7r_net_1\);
    
    \I2.PIPE7_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl31r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl31r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I153_Y_i_o4\ : AND3
      port map(A => \I2.N_33_adt_net_55021_\, B => \I2.N_57\, C
         => \I2.N_33_adt_net_55020_\, Y => \I2.N_33\);
    
    \I2.PIPE5_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_701_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl25r_net_1\);
    
    NWEN_pad : OB33PH
      port map(PAD => NWEN, A => NWEN_c);
    
    \I5.SSTATE1SE_2_0_908\ : AND2
      port map(A => TICKL0R_558, B => \I5.N_74\, Y => 
        \I5.sstate1_ns_el3r_adt_net_9195_\);
    
    \I2.DT_SRAMl3r\ : MUX2L
      port map(A => \I2.N_871\, B => \I2.PIPE2_DTl3r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl3r_net_1\);
    
    REGl204r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_105_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl204r\);
    
    \I3.VDBi_353\ : MUX2L
      port map(A => \I3.VDBil13r_net_1\, B => \I3.VDBi_57l13r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_353_net_1\);
    
    \I2.PIPE7_DTL27R_2794\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_87\);
    
    \I2.STOP_RDSRAM_453_i\ : AND3FFT
      port map(A => \I2.STATE3l1r_net_1\, B => 
        \I2.ROFFSET_0_sqmuxa_1\, C => 
        \I2.STOP_RDSRAM_453_i_adt_net_1077__net_1\, Y => 
        \I2.STOP_RDSRAM_453_i_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_1\ : OA21
      port map(A => \I2.N_140_0_ADT_NET_947__328\, B => 
        \I2.N_139_0_adt_net_55124_\, C => \I2.RAMDT4L5R_136\, Y
         => \I2.N_107_adt_net_256840_\);
    
    \I2.SUB9l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_570_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l2r_net_1\);
    
    \I2.OFFSET_37_1l1r\ : MUX2L
      port map(A => \REGl350r\, B => \REGl286r\, S => 
        \I2.PIPE7_DTL27R_66\, Y => \I2.N_636\);
    
    \I2.G_EVNT_NUM_n10_0_o2\ : NAND2
      port map(A => \I2.N_207_549\, B => \I2.G_EVNT_NUMl9r_net_1\, 
        Y => \I2.N_218\);
    
    \I2.DT_SRAM_0l4r\ : MUX2L
      port map(A => \I2.PIPE10_DTl4r_net_1\, B => 
        \I2.PIPE5_DTl4r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854220__net_1\, Y => 
        \I2.N_872\);
    
    \I1.un1_sbyte13_1_i_1_adt_net_854520_\ : BFR
      port map(A => \I1.un1_sbyte13_1_i_1\, Y => 
        \I1.un1_sbyte13_1_i_1_adt_net_854520__net_1\);
    
    \I2.OFFSET_37_10l0r\ : MUX2L
      port map(A => \I2.N_699\, B => \I2.N_691\, S => 
        \I2.PIPE7_DTL26R_351\, Y => \I2.N_707\);
    
    \I2.RAMAD1_12l1r\ : MUX2L
      port map(A => \I2.TDCDASl20r_net_1\, B => 
        \I2.TDCDBSl20r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855176__net_1\, Y => 
        \I2.RAMAD1_12l1r_net_1\);
    
    \I1.REG_74_12_300_m8_i_0\ : XOR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__761\, B
         => \I1.REG_74_12_300_N_13_Rd1__net_1\, Y => 
        \I1.REG_74_12_300_m8_i_0_adt_net_120083_\);
    
    \I3.REG1_139\ : MUX2L
      port map(A => VDB_inl6r, B => \I3.REG1l6r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG1_139_net_1\);
    
    \I3.VADm_0_a3l27r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl27r_net_1\, Y => \I3.VADml27r\);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_500\ : MUX2H
      port map(A => \I2.PIPE4_DTl22r_net_1\, B => 
        \I2.LSRAM_RADDRil1r_net_1\, S => \I2.N_4642\, Y => 
        \I2.LSRAM_RADDRi_500\);
    
    \I2.FCNT_105\ : NOR2
      port map(A => \I2.FCNT_c0\, B => \I2.un1_STATE1_22\, Y => 
        \I2.N_1236\);
    
    \I2.PIPE4_DTL6R_2963\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL6R_480\);
    
    REGl210r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_111_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl210r\);
    
    \I3.TCNT2_i_0_il2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT2_394_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT2_i_0_il2r_net_1\);
    
    \I2.PIPE2_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl7r_net_1\);
    
    \I1.REG_74_0_IVL388R_1805\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.REG_28_sqmuxa\, 
        Y => \I1.REG_74l388r_adt_net_111319_\);
    
    \I3.PIPEA1_325\ : MUX2L
      port map(A => \I3.PIPEA1l27r_net_1\, B => 
        \I3.PIPEA1_12l27r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, Y => 
        \I3.PIPEA1_325_net_1\);
    
    \I1.REG_74_0_ivl241r\ : AO21
      port map(A => \REGl241r\, B => \I1.N_113\, C => 
        \I1.REG_74l241r_adt_net_126641_\, Y => \I1.REG_74l241r\);
    
    \I2.STATEe_ns_il1r\ : AOI21FTF
      port map(A => \I2.CHAIN_ERRS_net_1\, B => 
        \I2.N_3496_adt_net_926__net_1\, C => 
        \I2.STATEe_ns_i_0_il1r\, Y => \I2.STATEe_ns_il1r_net_1\);
    
    \I2.PIPE4_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl9r_net_1\);
    
    \I2.DTE_1_866\ : MUX2L
      port map(A => \I2.DTE_1l28r_Rd1__net_1\, B => 
        \I2.DTE_21_1l28r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835988_Rd1__net_1\, Y => 
        \I2.DTE_1l28r\);
    
    \I2.LEAD_FLAG6l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_642_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl5r);
    
    \I3.VDBi_40_1l1r\ : MUX2L
      port map(A => REGl118r, B => \I3.VDBi_31l1r_net_1\, S => 
        \I3.REGMAPl16r_net_1\, Y => \I3.N_339\);
    
    \I3.REG_1l101r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_282_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl101r);
    
    \I3.VDBml23r\ : MUX2L
      port map(A => \I3.VDBil23r_net_1\, B => \I3.N_165\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml23r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I52_Y\ : AO21
      port map(A => \I2.N273\, B => \I2.N304_0_adt_net_86999_\, C
         => \I2.N300_0_adt_net_87051_\, Y => \I2.N302_0\);
    
    \I2.PIPE4_DTL9R_2955\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL9R_472\);
    
    \I1.N_347_adt_net_854788_\ : BFR
      port map(A => \I1.N_347\, Y => 
        \I1.N_347_adt_net_854788__net_1\);
    
    RAMAD_padl12r : OB33PH
      port map(PAD => RAMAD(12), A => RAMAD_cl12r);
    
    \I1.REG_74_0_iv_i_a2l208r\ : AO21
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, C => 
        \I1.N_1347_adt_net_129845_\, Y => \I1.N_1347\);
    
    \I3.REG_1l56r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_157_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl56r);
    
    \I2.DT_TEMPl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_769_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl8r_net_1\);
    
    \I2.DT_TEMPl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_763_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl2r_net_1\);
    
    \I2.DTO_1l17r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l17r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l17r_Rd1__net_1\);
    
    \I3.TCNT3_i_0_il4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT3_375_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT3_i_0_il4r_net_1\);
    
    \I2.N_2826_1_adt_net_40744_\ : OR3FTT
      port map(A => \I2.N_4641\, B => 
        \I2.STATE2l1r_adt_net_855132__net_1\, C => 
        \I2.N_2826_1_adt_net_40738__net_1\, Y => 
        \I2.N_2826_1_adt_net_40744__net_1\);
    
    REGl192r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_93_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl192r\);
    
    \I1.REG_5_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_243\, B => \I1.N_255\, Y => 
        \I1.REG_5_sqmuxa\);
    
    \I3.un3_noe32wi_0_a2_i\ : OR2
      port map(A => NOE16W_c, B => \I3.LWORDS_net_1\, Y => 
        NOE32W_c);
    
    \I2.PIPE10_DT_17_i_0l18r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855592__net_1\, B => 
        \I2.PIPE9_DTl18r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l18r_net_1\);
    
    \I5.sstate1l6r\ : DFFC
      port map(CLK => CLK_c, D => \I5.N_98\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l6r_net_1\);
    
    \I2.DTO_9_iv_ml28r_adt_net_857_\ : OAI21TTF
      port map(A => \I2.N_4283_i_0_adt_net_854968__net_1\, B => 
        \I2.DT_TEMPl28r_net_1\, C => 
        \I2.DTO_9_iv_ml28r_adt_net_28906__net_1\, Y => 
        \I2.DTO_9_iv_ml28r_adt_net_857__net_1\);
    
    \I2.MIC_ERR_REGSl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_355_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl26r_net_1\);
    
    \I5.SSTATE1SE_7_0_0_905\ : AO21FTF
      port map(A => TICKL0R_558, B => \I5.sstate1l5r_net_1\, C
         => \I5.N_130\, Y => \I5.sstate1_ns_el8r_adt_net_8891_\);
    
    FID_padl29r : OB33PH
      port map(PAD => FID(29), A => FID_cl29r);
    
    \I3.un5_noe16ri_0_i_a3\ : AOI21TTF
      port map(A => \I3.N_268\, B => \I3.N_290_adt_net_4891_\, C
         => NOEAD_c, Y => NOE16R_c);
    
    \I3.PULSE_330_adt_net_854732_\ : BFR
      port map(A => \I3.PULSE_330_net_1\, Y => 
        \I3.PULSE_330_adt_net_854732__net_1\);
    
    \I2.EVNT_NUMl10r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_953_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl10r_net_1\);
    
    \I2.BNCID_VECT_tile_0_I_5_i\ : INV
      port map(A => TDCTRG_c, Y => \I2.TDCTRG_c_i_0\);
    
    \I1.REG_74_0_ivl381r\ : AO21
      port map(A => \REGl381r\, B => \I1.N_257\, C => 
        \I1.REG_74l381r_adt_net_111921_\, Y => \I1.REG_74l381r\);
    
    \I2.DTO_16_1l6r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l6r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l6r_Rd1__net_1\);
    
    \I2.PIPE10_DT_17_il16r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l3r_net_1\, C => \I2.PIPE10_DT_17_i_0l16r_net_1\, 
        Y => \I2.N_3802\);
    
    \I1.REG_74_2_0l404r\ : NOR2
      port map(A => \I1.PAGECNT_320_adt_net_854872__net_1\, B => 
        \I1.PAGECNT_319_net_1\, Y => \I1.REG_74_2_0l404r_Ra1_\);
    
    \I2.LEAD_FLAG6_644_1599\ : NOR2FT
      port map(A => LEAD_FLAGl7r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_644_adt_net_63844_\);
    
    \I3.VDBi_342\ : MUX2L
      port map(A => \I3.VDBil2r_net_1\, B => \I3.VDBi_57l2r\, S
         => \I3.un1_STATE1_13_1_adt_net_1351__net_1\, Y => 
        \I3.VDBi_342_net_1\);
    
    \I3.VDBI_16_M_I_2L3R_2254\ : AO21FTT
      port map(A => REGl35r, B => \I3.REGMAPL7R_460\, C => 
        \I3.N_1907_265\, Y => 
        \I3.VDBi_16_m_i_2_il3r_adt_net_144610_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I113_Y\ : NOR3
      port map(A => \I2.N330\, B => \I2.I92_un1_Y\, C => 
        \I2.I113_un1_Y\, Y => \I2.N451_i\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I65_Y\ : AND2
      port map(A => \I2.N255_0\, B => \I2.N252_0\, Y => \I2.N315\);
    
    \I3.VDBOFFA_31_IV_0L1R_2608\ : AO21
      port map(A => \REGl190r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.VDBoffa_31l1r_adt_net_164408_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164449_\);
    
    \I2.OFFSET_37_24l1r\ : MUX2L
      port map(A => \I2.N_812\, B => \I2.N_804\, S => 
        \I2.PIPE7_DTL26R_360\, Y => \I2.N_820\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I18_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L5R_820\, B => 
        \I2.PIPE4_DTl18r_net_1\, Y => \I2.N_63\);
    
    \I5.SBYTEl6r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_71_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl6r_net_1\);
    
    \I3.N_1645_i_i_o3_1\ : OR2FT
      port map(A => \I3.STATE1_IPL9R_419\, B => 
        \I3.REGMAPL0R_421\, Y => \I3.N_1905_1\);
    
    \I2.DT_SRAMl29r\ : MUX2L
      port map(A => \I2.N_897\, B => \I2.PIPE2_DTl29r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl29r_net_1\);
    
    \I3.VDBi_57l7r_adt_net_142952_\ : NOR2FT
      port map(A => REGl39r, B => \I3.N_2033\, Y => 
        \I3.VDBi_57l7r_adt_net_142952__net_1\);
    
    \I1.REG_1_163\ : MUX2H
      port map(A => \REGl262r\, B => \I1.REG_74l262r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y => 
        \I1.REG_1_163_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I25_Y\ : OAI21FTT
      port map(A => \I2.N_3558_i_net_1\, B => \I2.SUB8l15r_net_1\, 
        C => \I2.N288_adt_net_68878_\, Y => \I2.N290\);
    
    \I2.PIPE8_DT_21l5r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl5r\, B => \I2.N_571\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l5r_net_1\);
    
    \I2.PIPE2_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl30r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl30r_net_1\);
    
    \I1.REG_74_0_IV_0L369R_1832\ : AND2
      port map(A => \FBOUTl4r\, B => \I1.N_593\, Y => 
        \I1.REG_74l369r_adt_net_113568_\);
    
    \I3.VDBi_40_0_a3_0l5r\ : NOR3
      port map(A => \I3.N_1948\, B => 
        \I3.VDBi_31_i_a3_0_1l5r_adt_net_143649_\, C => 
        \I3.VDBi_31_i_a3_0_1l5r_adt_net_143654_\, Y => 
        \I3.N_1772_adt_net_143698_\);
    
    \I3.PIPEA_8_0l14r\ : MUX2L
      port map(A => DPR_cl14r, B => \I3.PIPEA1l14r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855348__net_1\, Y => \I3.N_223\);
    
    \I3.DS_i_a3\ : OR2
      port map(A => DS0B_c, B => DS1B_c, Y => \I3.N_95\);
    
    \I2.N346_adt_net_4075_\ : AO21
      port map(A => \I2.N232\, B => 
        \I2.N346_adt_net_69448__net_1\, C => \I2.N311\, Y => 
        \I2.N346_adt_net_4075__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I3_P0N_i_o3\ : NOR2
      port map(A => \I2.RAMDT4L10R_766\, B => 
        \I2.PIPE4_DTl3r_adt_net_854548__net_1\, Y => \I2.N_28_0\);
    
    \I3.VDBi_57l8r_adt_net_142596_\ : AO21
      port map(A => \I3.N_2271\, B => \I3.N_2037\, C => 
        \I3.VDBi_57l8r_adt_net_142588__net_1\, Y => 
        \I3.VDBi_57l8r_adt_net_142596__net_1\);
    
    \I2.STATE3l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3l3r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL2R_1512\ : AO21FTT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        B => \I2.PIPE1_DT_12l2r_net_1\, C => 
        \I2.PIPE1_DT_42l2r_adt_net_51829_\, Y => 
        \I2.PIPE1_DT_42l2r_adt_net_51838_\);
    
    \I3.REGMAPL57R_2992\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un231_reg_ads_0_a2_4_a3_net_1\, Q => 
        \I3.REGMAPL57R_539\);
    
    \I2.CRC32_808\ : MUX2L
      port map(A => \I2.CRC32l13r_net_1\, B => \I2.N_3930\, S => 
        \I2.N_2826_1_ADT_NET_794__331\, Y => \I2.CRC32_808_net_1\);
    
    \I3.REG_1l57r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_158_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl57r);
    
    REGl352r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_253_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl352r\);
    
    \I1.REG_74_0_IVL243R_1983\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_10_sqmuxa_adt_net_854716__net_1\, Y => 
        \I1.REG_74l243r_adt_net_126469_\);
    
    \I3.VDBi_55l3r\ : MUX2H
      port map(A => \I3.VDBil3r_net_1\, B => \I3.RAMDTSl3r_net_1\, 
        S => \I3.N_57_i_0_0_adt_net_854688__net_1\, Y => 
        \I3.VDBi_55l3r_net_1\);
    
    VAD_padl29r : IOB33PH
      port map(PAD => VAD(29), A => \I3.VADml29r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl29r);
    
    \I3.TCNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_383_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTl1r_net_1\);
    
    \I2.PIPE8_DT_21l1r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl1r\, B => \I2.N_567\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l1r_net_1\);
    
    REGl299r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_200_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl299r\);
    
    \I3.un1_REGMAP_30_0_a2_0\ : NOR3FTT
      port map(A => \I3.un1_REGMAP_30_0_a2_0_adt_net_134424_\, B
         => \I3.REGMAP_I_0_IL30R_772\, C => \I3.REGMAPL29R_771\, 
        Y => \I3.un1_REGMAP_30_0_a2_0_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I172_Y\ : XOR2
      port map(A => \I2.N357_0\, B => 
        \I2.ADD_21x21_fast_I172_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l2r\);
    
    \I2.OFFSET_37_27l3r\ : MUX2L
      port map(A => \I2.N_838\, B => \I2.N_822\, S => 
        \I2.PIPE7_DTL25R_687\, Y => \I2.N_846\);
    
    \I2.RAMAD_4_0l3r\ : MUX2H
      port map(A => \I2.RAMAD1l3r_net_1\, B => RAMAD_VMEl3r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_530\);
    
    \I2.SUB9_1_ADD_18x18_fast_I5_P0N\ : OR2
      port map(A => \I2.N_3543_i_i\, B => \I2.G_1_0\, Y => 
        \I2.N241\);
    
    \I2.SUB9l12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_580_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l12r_net_1\);
    
    \I2.PIPE5_DT_682\ : MUX2L
      port map(A => \I2.PIPE5_DTl6r_net_1\, B => 
        \I2.PIPE5_DT_6l6r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_682_net_1\);
    
    \I3.un224_reg_ads_0_a2_3_a3\ : NOR3
      port map(A => \I3.N_546\, B => \I3.N_558\, C => \I3.N_578\, 
        Y => \I3.un224_reg_ads_0_a2_3_a3_net_1\);
    
    \I3.PIPEA1_12l22r\ : AND2
      port map(A => DPR_cl22r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854496__net_1\, Y => 
        \I3.PIPEA1_12l22r_net_1\);
    
    \I3.VDBoffb_52\ : OR3
      port map(A => \I3.VDBoffb_52_adt_net_163170_\, B => 
        \I3.VDBoffb_30l0r_adt_net_163129_\, C => 
        \I3.VDBoffb_30l0r_adt_net_163130_\, Y => 
        \I3.VDBoffb_52_net_1\);
    
    \I2.PIPE6_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_480_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl26r_net_1\);
    
    \I2.PIPE8_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_559_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl31r_net_1\);
    
    \I2.L2SERV_922\ : XOR2
      port map(A => \I2.RPAGEl12r\, B => \I2.L2SERVe\, Y => 
        \I2.L2SERV_922_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I99_Y\ : AO21
      port map(A => \I2.N346_adt_net_4075__net_1\, B => 
        \I2.N463_adt_net_70886_\, C => \I2.N338\, Y => \I2.N463\);
    
    \I2.MIC_ERR_REGS_365\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl37r_net_1\, B => 
        \I2.MIC_ERR_REGSl36r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_365_net_1\);
    
    \I5.AIR_WDATAl8r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_58_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl8r_net_1\);
    
    \I1.REG_1_166\ : MUX2H
      port map(A => \REGl265r\, B => \I1.REG_74l265r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y => 
        \I1.REG_1_166_net_1\);
    
    \I2.TRGCNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGCNT_n1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGCNT_i_0_il1r\);
    
    \I2.PIPE1_DT_42_1_IVL23R_1375\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855032__net_1\, 
        B => \I2.TDCDASl23r_net_1\, Y => 
        \I2.PIPE1_DT_42l23r_adt_net_46639_\);
    
    \I1.BYTECNT_312\ : MUX2H
      port map(A => \I1.BYTECNTl2r_adt_net_855020__net_1\, B => 
        \I1.N_174\, S => \I1.N_1383\, Y => \I1.BYTECNT_312_net_1\);
    
    \I2.FID_7_0_iv_0l5r\ : OAI21FTF
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl5r_net_1\, 
        C => \I2.FID_7_0_iv_0l5r_adt_net_93017_\, Y => 
        \I2.FID_7_0_iv_0l5r_net_1\);
    
    \I2.CRC32l29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_824_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l29r_net_1\);
    
    \I3.REG_0_sqmuxa_3_0_a2_0_a3\ : AND2
      port map(A => \I3.REGMAPl55r_net_1\, B => 
        \I3.N_1906_i_0_0_adt_net_855636__net_1\, Y => 
        \I3.REG_0_sqmuxa_3\);
    
    \I2.FID_7_0_ivl15r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl15r_net_1\, 
        C => \I2.FID_7l15r_adt_net_17901_\, Y => \I2.FID_7l15r\);
    
    \I2.DTO_16_1_IV_0L7R_1186\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.DTE_2_1l7r_net_1\, Y => 
        \I2.DTO_16_1l7r_adt_net_33728_\);
    
    \I2.DTE_21_1_iv_0_0l22r\ : AO21
      port map(A => \I2.DTE_1l22r_Rd1__net_1\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835168_Rd1__net_1\, 
        C => \I2.DTE_21_1l22r_adt_net_37395_Rd1__net_1\, Y => 
        \I2.DTE_21_1l22r_Rd1_\);
    
    \I1.REG_74_0_iv_i_a2l200r\ : AO21
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_1339_adt_net_130533_\, Y => \I1.N_1339\);
    
    \I5.REG_1l431r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_44_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl431r);
    
    \I1.REG_74_0_ivl310r\ : AO21
      port map(A => \REGl310r\, B => \I1.N_185\, C => 
        \I1.REG_74l310r_adt_net_119905_\, Y => \I1.REG_74l310r\);
    
    \I2.WOFFSETl0r_adt_net_854644_\ : BFR
      port map(A => \I2.WOFFSETl0r_net_1\, Y => 
        \I2.WOFFSETl0r_adt_net_854644__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I178_Y_2730\ : AND2
      port map(A => \I2.N297_0\, B => \I2.N300_0\, Y => 
        \I2.N479_adt_net_642266_\);
    
    \I1.REG_1_81\ : MUX2H
      port map(A => \REGl180r\, B => \I1.REG_74l180r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\, Y
         => \I1.REG_1_81_net_1\);
    
    \I3.VDBOFFA_31_IV_0L0R_2634\ : OR3
      port map(A => \I3.VDBoffa_31l0r_adt_net_164645_\, B => 
        \I3.VDBoffa_31l0r_adt_net_164639_\, C => 
        \I3.VDBoffa_31l0r_adt_net_164640_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164649_\);
    
    \I3.un1_STATE1_5_i_a2_0_a3\ : NOR2
      port map(A => \I3.N_311\, B => \I3.STATE1_ipl7r\, Y => 
        \I3.N_1409\);
    
    \I2.EVNT_REJ_2_SQMUXA_1060\ : AND3FTT
      port map(A => \I2.un21_sram_empty_NE_net_1\, B => 
        \I2.N_118_i_1_adt_net_1122__net_1\, C => 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26950_\, Y => 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26951_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I177_Y_2688\ : AO21
      port map(A => \I2.N285\, B => \I2.N296_0_adt_net_86398_\, C
         => \I2.N475_adt_net_87328__net_1\, Y => 
        \I2.N477_adt_net_438351_\);
    
    \I2.N_2826_1_ADT_NET_794__2889\ : OAI21FTF
      port map(A => \I2.N_4261_304\, B => \I2.N_4282\, C => 
        \I2.N_2826_1_adt_net_40744__net_1\, Y => 
        \I2.N_2826_1_ADT_NET_794__330\);
    
    \I2.FID_7_0_ivl17r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl17r_net_1\, 
        C => \I2.FID_7l17r_adt_net_17713_\, Y => \I2.FID_7l17r\);
    
    \I2.LSRAM_WADDRl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_WADDR_382_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_WADDRl1r_net_1\);
    
    REGl391r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_292_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl391r\);
    
    \I2.MIC_ERR_REGSl45r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_374_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl45r_net_1\);
    
    \I3.VDBI_57_0_IV_0L20R_2170\ : AO21
      port map(A => \I3.VDBil20r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l20r_adt_net_139281_\, Y => 
        \I3.VDBi_57l20r_adt_net_139291_\);
    
    \I2.PIPE1_DT_42_1_ivl17r\ : OR3
      port map(A => \I2.PIPE1_DT_42l17r_adt_net_47637_\, B => 
        \I2.PIPE1_DT_42l17r_adt_net_47649_\, C => 
        \I2.PIPE1_DT_42l17r_adt_net_47650_\, Y => 
        \I2.PIPE1_DT_42l17r\);
    
    \I2.PIPE6_DT_473\ : MUX2H
      port map(A => \I2.PIPE5_DTl19r_net_1\, B => 
        \I2.PIPE6_DTl19r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_473_net_1\);
    
    \I2.DTE_21_1_IV_0L6R_1320\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855124__net_1\, B => 
        \I2.EVNT_WORDl2r_net_1\, Y => 
        \I2.DTE_21_1l6r_adt_net_38967_\);
    
    \I2.PIPE1_DT_42_1_IVL11R_1458\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855228__net_1\, B => 
        \I2.MIC_ERR_REGSl11r_net_1\, C => 
        \I2.PIPE1_DT_42l11r_adt_net_49703_\, Y => 
        \I2.PIPE1_DT_42l11r_adt_net_49704_\);
    
    \I3.TCNT3l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT3_374_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT3l5r_net_1\);
    
    \I3.un136_reg_ads_0_a2_2_a2\ : OR2
      port map(A => \I3.N_555\, B => \I3.N_549\, Y => \I3.N_584\);
    
    \I2.PIPE10_DT_616\ : MUX2L
      port map(A => \I2.PIPE10_DTl11r_net_1\, B => 
        \I2.PIPE9_DTl11r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_616_net_1\);
    
    \I1.N_1169_adt_net_854824_\ : BFR
      port map(A => \I1.N_1169\, Y => 
        \I1.N_1169_adt_net_854824__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I119_Y_i_o4\ : OR2
      port map(A => 
        \I2.N_3_0_adt_net_1070__adt_net_855604__net_1\, B => 
        \I2.N_3_0_adt_net_59703_\, Y => \I2.N_3_0\);
    
    \I2.SUB9_574\ : MUX2H
      port map(A => \I2.SUB9l6r_net_1\, B => \I2.SUB9_1l6r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_574_net_1\);
    
    \I3.un47_reg_ads_0_a2_0_a2_994\ : OR2FT
      port map(A => \I3.WRITES_8\, B => \I3.N_546_374\, Y => 
        \I3.N_547_372\);
    
    \I2.L2TYPE_4_il11r\ : OAI21FTF
      port map(A => \I2.L2TYPEl11r_net_1\, B => \I2.N_4467\, C
         => \I2.N_4441_adt_net_67338_\, Y => \I2.N_4441\);
    
    DTO_padl5r : IOB33PH
      port map(PAD => DTO(5), A => \I2.DTO_1l5r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl5r);
    
    \I1.ISCK_0_sqmuxa_0_0_a2\ : NAND3FFT
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__863\, B => 
        \I1.N_359\, C => \I1.sstatel4r_net_1\, Y => \I1.N_656\);
    
    \I3.VDBI_57_0_IV_0_0L8R_2222\ : AND2
      port map(A => \I3.PIPEAl8r_net_1\, B => \I3.N_90_i_0\, Y
         => \I3.VDBi_57l8r_adt_net_142780_\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__3103\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__889\);
    
    \I2.PIPE6_DT_481\ : MUX2H
      port map(A => \I2.PIPE5_DTl27r_net_1\, B => 
        \I2.PIPE6_DTl27r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_481_net_1\);
    
    \I2.FID_7_ivl2r\ : OR2
      port map(A => \I2.FID_7l2r_adt_net_93358_\, B => 
        \I2.FID_7l2r_adt_net_93359_\, Y => \I2.FID_7l2r\);
    
    \I1.REG_74_0_ivl216r\ : AO21
      port map(A => \REGl216r\, B => \I1.N_89\, C => 
        \I1.REG_74l216r_adt_net_129120_\, Y => \I1.REG_74l216r\);
    
    \I3.REGMAPL7R_2943\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un33_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL7R_460\);
    
    \I2.OFFSET_37_20l0r\ : MUX2L
      port map(A => \I2.N_779\, B => \I2.N_771\, S => 
        \I2.PIPE7_DTL26R_356\, Y => \I2.N_787\);
    
    TDCDRYA_pad : IB33
      port map(PAD => TDCDRYA, Y => TDCDRYA_c);
    
    \I3.VDBOFFB_30_IV_0L7R_2360\ : AO21
      port map(A => \REGl316r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        C => \I3.VDBoffb_30l7r_adt_net_161764_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161793_\);
    
    \I3.REGMAPl1r_1618\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un10_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL1R_725\);
    
    ADO_padl4r : OB33PH
      port map(PAD => ADO(4), A => ADO_cl4r);
    
    \I2.DTO_16_1_ivl23r\ : OR2
      port map(A => \I2.DTO_16_1l23r_adt_net_30115_\, B => 
        \I2.DTO_16_1l23r_adt_net_30116_\, Y => \I2.DTO_16_1l23r\);
    
    \I3.un224_reg_ads_0_a2_3_a2_995\ : NAND2
      port map(A => \I3.LWORDS_787\, B => \I3.N_545\, Y => 
        \I3.N_546_373\);
    
    \I1.BITCNTL0R_3051\ : DFFC
      port map(CLK => CLK_c, D => \I1.BITCNT_317_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BITCNTL0R_805\);
    
    \I3.STATE2_0_sqmuxa_2_i_o3_877\ : NAND2FT
      port map(A => \I3.DSS_718\, B => \I3.N_258\, Y => 
        \I3.N_281_255\);
    
    \I5.COMMANDl12r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_49_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl12r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L0R_2477\ : AND2
      port map(A => \REGl285r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163086_\);
    
    \I2.un1_STATE1_9_i_a3\ : NOR3
      port map(A => \I2.STATE1l18r_net_1\, B => 
        \I2.STATE1l10r_net_1\, C => \I2.STATE1l13r_net_1\, Y => 
        \I2.N_3306\);
    
    \I2.DT_TEMPl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_772_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl11r_net_1\);
    
    \I2.RAMAD_4l5r\ : MUX2L
      port map(A => \I2.N_532\, B => \I1.BYTECNTl5r_net_1\, S => 
        LOAD_RES, Y => \I2.RAMAD_4l5r_net_1\);
    
    \I3.PULSE_331\ : AO21
      port map(A => \I3.N_311_adt_net_854748__net_1\, B => 
        \I3.N_118_adt_net_147476_\, C => 
        \I3.PULSE_331_adt_net_147557_\, Y => \I3.PULSE_331_net_1\);
    
    \I3.VDBI_57_0_IVL10R_2215\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => 
        \I3.VDBi_55l10r_net_1\, C => 
        \I3.VDBi_57l10r_adt_net_141883_\, Y => 
        \I3.VDBi_57l10r_adt_net_141884_\);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854260_\ : BFR
      port map(A => \I2.WR_SRAM_2_adt_net_748__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854260__net_1\);
    
    \I2.PIPE8_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_538_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl10r_net_1\);
    
    \I1.N_161_adt_net_121649_\ : OAI21FTF
      port map(A => \I1.REG_74_12_300_N_11_adt_net_120111_\, B
         => \I1.REG_74_12_284_m10_i_0_i\, C => \I1.N_1370\, Y => 
        \I1.N_161_adt_net_121649__net_1\);
    
    \I3.PIPEAl29r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEA_260_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl29r_net_1\);
    
    \I2.ADOl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl7r);
    
    \I5.DATAl15r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l15r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl132r);
    
    \I2.PIPE1_DT_42_1_IVL19R_1397\ : NOR2FT
      port map(A => REGl423r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, Y => 
        \I2.PIPE1_DT_42l19r_adt_net_47255_\);
    
    \I1.REG_74_12_0l188r_894\ : NAND3
      port map(A => \I1.N_347_adt_net_854788__net_1\, B => 
        \I1.REG_74_i_o2_i_0l364r_net_1\, C => \I1.N_57_9_i\, Y
         => \I1.N_65_12_272\);
    
    \I1.REG_74_0_IVL274R_1949\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, Y => 
        \I1.REG_74l274r_adt_net_123474_\);
    
    \I5.TEMPDATAl2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_76_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl2r_net_1\);
    
    \I3.PULSEl8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_338_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl8r);
    
    \I2.LSRAM_IN_412\ : MUX2L
      port map(A => \I2.PIPE5_DTl28r_net_1\, B => 
        \I2.LSRAM_INl28r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_412_net_1\);
    
    \I1.PAGECNTL9R_2850\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854856__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL9R_244\);
    
    \I2.STATE1_ns_il9r\ : OA21TTF
      port map(A => \I2.CHAINA_EN244_i_adt_net_855260__net_1\, B
         => \I2.END_CHAINA1_net_1\, C => \I2.N_3288\, Y => 
        \I2.N_3208_i_0\);
    
    \I2.un1_DTO_cl_0_sqmuxa_0_0_o2_1\ : OR2FT
      port map(A => \I2.N_2870\, B => 
        \I2.un1_DTO_cl_0_sqmuxa_adt_net_22686_\, Y => 
        \I2.un1_DTO_cl_0_sqmuxa\);
    
    \I2.FIDl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_416_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl0r);
    
    \I2.DTO_16_1_iv_0_0l12r\ : OR2
      port map(A => \I2.DTO_16_1l12r_adt_net_32633_\, B => 
        \I2.DTO_16_1l12r_adt_net_32634_\, Y => \I2.DTO_16_1l12r\);
    
    \I2.un1_TOKOUT_FL_0_sqmuxa_0_o3_0\ : OR2
      port map(A => \I2.STATE1L8R_648\, B => \I2.STATE1L13R_601\, 
        Y => \I2.N_3890\);
    
    \I3.TCNT_N1_0_0_2136\ : XOR2FT
      port map(A => \I3.TCNTl0r_net_1\, B => \I3.TCNTl1r_net_1\, 
        Y => \I3.TCNT_n1_adt_net_137059_\);
    
    REGl390r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_291_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl390r\);
    
    \I5.SDAin_m_1\ : NOR3FFT
      port map(A => \I5.sstate1l1r_net_1\, B => \I5.N_101\, C => 
        \I5.COMMANDl0r_net_1\, Y => \I5.SDAin_m_1_net_1\);
    
    \I5.COMMAND_4l1r\ : MUX2L
      port map(A => \I5.AIR_WDATAl1r_net_1\, B => REGl102r, S => 
        REGl7r, Y => \I5.COMMAND_4l1r_net_1\);
    
    \I3.REG_1_215\ : MUX2L
      port map(A => VDB_inl2r, B => REGl408r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_215_0\);
    
    \I2.PIPE9_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_277_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl8r_net_1\);
    
    \I3.UN1_STATE2_15_1_ADT_NET_1342__2859\ : OR2
      port map(A => \I3.STATE2_nsl0r_adt_net_136048_\, B => 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\, Y => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__253\);
    
    \I1.REG_1_290\ : MUX2H
      port map(A => \REGl389r\, B => \I1.REG_74l389r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y => 
        \I1.REG_1_290_net_1\);
    
    \I2.L2TYPEl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_591_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl2r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L4R_2409\ : AO21
      port map(A => \REGl401r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l4r_adt_net_162314_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162358_\);
    
    \I3.VDBOFFB_56_2420\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl4r_net_1\, Y => 
        \I3.VDBoffb_56_adt_net_162410_\);
    
    \I2.DTE_21_1_IV_0L19R_1266\ : AO21
      port map(A => \I2.DT_TEMPl19r_net_1\, B => \I2.N_4038\, C
         => \I2.DTE_21_1l19r_adt_net_37709_\, Y => 
        \I2.DTE_21_1l19r_adt_net_37723_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I153_Y\ : XOR2FT
      port map(A => \I2.N445_i\, B => 
        \I2.ADD_18x18_fast_I153_Y_0\, Y => \I2.SUB9_1l16r\);
    
    \I3.REG_44_IL85R_2306\ : AOI21FTT
      port map(A => REGl85r, B => \I3.N_98_0\, C => \I3.N_1665\, 
        Y => \I3.N_1631_adt_net_150433_\);
    
    \I1.REG_74L388R_1802\ : AND2FT
      port map(A => \I1.N_330_i_0_i\, B => \I1.N_584\, Y => 
        \I1.N_257_adt_net_111267_\);
    
    \I3.VASl15r_968\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_77_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VAS_I_0_IL15R_346\);
    
    \I2.SUB9_1_ADD_18x18_fast_I63_Y\ : AND2
      port map(A => \I2.N300\, B => \I2.N296\, Y => \I2.N331\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I58_Y\ : AO21
      port map(A => \I2.N264_0\, B => \I2.N308_0_adt_net_86497_\, 
        C => \I2.N308_0_adt_net_86492_\, Y => \I2.N308_0\);
    
    \I3.VDBil18r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_358_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil18r_net_1\);
    
    \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146197_\ : AND2
      port map(A => \I3.N_2034\, B => \I3.RAMDTSl0r_net_1\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146197__net_1\);
    
    REGl284r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_185_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl284r\);
    
    \I2.PIPE7_DTL27R_2795\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_88\);
    
    \I3.UN224_REG_ADS_0_A2_3_A2_2_2647\ : AND3FFT
      port map(A => \I3.VAS_I_0_IL7R_747\, B => \I3.VASL6R_748\, 
        C => \I3.N_545_adt_net_165680_\, Y => 
        \I3.N_545_adt_net_165682_\);
    
    \I3.VDBI_57_0_IVL22R_2162\ : AO21
      port map(A => \I3.VDBil22r_net_1\, B => 
        \I3.N_1910_0_adt_net_854344__net_1\, C => 
        \I3.VDBi_57l22r_adt_net_139083_\, Y => 
        \I3.VDBi_57l22r_adt_net_139087_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I5_P0N_i_a4\ : OR2
      port map(A => \I2.RAMDT4L5R_809\, B => 
        \I2.PIPE4_DTl5r_adt_net_854420__net_1\, Y => \I2.N_89\);
    
    \I3.VADm_0_a3l25r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl25r_net_1\, Y => \I3.VADml25r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I190_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_799\, B => 
        \I2.PIPE4_DTl20r_net_1\, Y => 
        \I2.ADD_21x21_fast_I190_Y_0_0\);
    
    \I2.PIPE8_DT_556\ : MUX2L
      port map(A => \I2.PIPE8_DTl28r_net_1\, B => \I2.N_4399\, S
         => \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_556_net_1\);
    
    \I2.PIPE8_DT_21l9r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl9r\, B => \I2.N_575\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l9r_net_1\);
    
    \I2.PIPE10_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_625_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl20r_net_1\);
    
    \I3.VDBi_31l17r\ : MUX2L
      port map(A => \I3.REGl150r\, B => \I3.VDBi_20l17r\, S => 
        \I3.REGMAPl17r_adt_net_854280__net_1\, Y => 
        \I3.VDBi_31l17r_net_1\);
    
    \I3.un5_noe16ri_0_i_o2\ : AND2
      port map(A => \I3.N_268\, B => \I3.N_290_adt_net_4891_\, Y
         => \I3.N_290\);
    
    \I3.VAS_73\ : MUX2L
      port map(A => VAD_inl11r, B => \I3.VASl11r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_73_net_1\);
    
    \I2.N_4667_1_ADT_NET_1046__2755\ : OAI21FTF
      port map(A => \I2.N_4261\, B => \I2.N_4283_I_0_41\, C => 
        \I2.STATE2L2R_589\, Y => \I2.N_4667_1_ADT_NET_1046__31\);
    
    \I3.REGMAPl0r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un2_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl0r_net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854568_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854568__net_1\);
    
    \I2.CRC32_818\ : MUX2L
      port map(A => \I2.CRC32l23r_net_1\, B => \I2.N_3940\, S => 
        \I2.N_2826_1_ADT_NET_794__330\, Y => \I2.CRC32_818_net_1\);
    
    \I3.un54_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.un231_reg_ads_1\, B => \I3.N_573\, Y => 
        \I3.un54_reg_ads_0_a2_1_a3_net_1\);
    
    \I1.REG_74l244r\ : OR3
      port map(A => \I1.N_201_9\, B => 
        \I1.N_113_adt_net_3714__net_1\, C => \I1.REG_9_sqmuxa\, Y
         => \I1.N_113\);
    
    \I3.REG3l405r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_226_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l405r_net_1\);
    
    \I2.DTE_21_1_IV_0_IL25R_1243\ : AND2
      port map(A => \I2.DT_TEMPl25r_net_1\, B => \I2.N_4038_233\, 
        Y => \I2.N_4644_adt_net_37053_\);
    
    \I1.REG_74_0_IVL361R_1846\ : AND2
      port map(A => \FBOUTl4r\, B => \I1.REG_25_sqmuxa\, Y => 
        \I1.REG_74l361r_adt_net_114783_\);
    
    \I2.BNCID_VECTROR_9_TZ_1420\ : AO21
      port map(A => \I2.BNCID_VECTra14_1_net_1\, B => 
        \I2.BNCID_VECTro_14\, C => 
        \I2.BNCID_VECTror_9_tz_adt_net_48091_\, Y => 
        \I2.BNCID_VECTror_9_tz_adt_net_48099_\);
    
    \I5.SDAOUT_12_IV_0_A2_917\ : OR3FFT
      port map(A => \I5.SDAout_net_1\, B => 
        \I5.N_64_adt_net_855868__net_1\, C => 
        \I5.sstate1l11r_net_1\, Y => \I5.N_150_adt_net_9846_\);
    
    \I1.REG_1_293\ : MUX2H
      port map(A => \REGl392r\, B => \I1.REG_74l392r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y => 
        \I1.REG_1_293_net_1\);
    
    \I3.REG_1l408r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_215_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl408r);
    
    \I2.PIPE6_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_457_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl3r_net_1\);
    
    \I2.MIC_REG3l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_321_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l4r_net_1\);
    
    \I2.PIPE4_DTl19r_1527\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl19r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL19R_634\);
    
    \I2.NWPIPE8\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, 
        SET => CLEAR_STAT_i_0, Q => \I2.NWPIPE8_I_0_I_0_0_5\);
    
    \I2.L2TYPE_600\ : MUX2L
      port map(A => \I2.L2TYPEl11r_net_1\, B => \I2.N_4441\, S
         => \I2.N_4482_0\, Y => \I2.L2TYPE_600_net_1\);
    
    VAD_padl18r : OTB33PH
      port map(PAD => VAD(18), A => \I3.VADml18r\, EN => 
        NOEAD_c_i_0);
    
    \I2.PIPE7_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl23r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl23r_net_1\);
    
    \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_28030_\ : NAND2
      port map(A => NOESRAME_C_833, B => \I2.STATE2L5R_508\, Y
         => 
        \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_28030__net_1\);
    
    \I2.PIPE9_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_274_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl5r_net_1\);
    
    TDCDA_padl4r : IB33
      port map(PAD => TDCDA(4), Y => TDCDA_cl4r);
    
    \I3.UN1_STATE1_13_1_ADT_NET_1351__2802\ : OR3
      port map(A => \I3.un1_STATE1_13_1_adt_net_137890__net_1\, B
         => \I3.un1_STATE1_13_1_adt_net_137896__net_1\, C => 
        \I3.un1_STATE1_13_1_adt_net_137902__net_1\, Y => 
        \I3.UN1_STATE1_13_1_ADT_NET_1351__114\);
    
    \I3.REG_1l417r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_224_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl417r);
    
    \I2.DTO_1l6r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l6r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l6r_Rd1__net_1\);
    
    \I3.VDBI_57_IVL4R_2252\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => 
        \I3.VDBi_55l4r_net_1\, C => 
        \I3.VDBi_57l4r_adt_net_144439_\, Y => 
        \I3.VDBi_57l4r_adt_net_144440_\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855032_\ : BFR
      port map(A => \I2.PIPE1_DT_2_SQMUXA_ADT_NET_803__299\, Y
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855032__net_1\);
    
    \I1.ISI_54\ : MUX2H
      port map(A => F_SI_c, B => \I1.N_1193\, S => \I1.N_1375\, Y
         => \I1.ISI_54_net_1\);
    
    \I3.VDBOFFA_45_2618\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal1r_net_1\, Y => 
        \I3.VDBoffa_45_adt_net_164498_\);
    
    VAD_padl23r : OTB33PH
      port map(PAD => VAD(23), A => \I3.VADml23r\, EN => 
        NOEAD_c_i_0);
    
    \I2.TRGSERV_2_I_17\ : XOR2
      port map(A => \I2.DWACT_ADD_CI_0_g_array_12_0l0r\, B => 
        \I2.TRGSERVl3r_net_1\, Y => \I2.TRGSERV_2l3r\);
    
    \I2.RAMAD1_12l2r\ : MUX2L
      port map(A => \I2.TDCDASl0r_net_1\, B => 
        \I2.TDCDBSl0r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855176__net_1\, Y => 
        \I2.RAMAD1_12l2r_net_1\);
    
    \I2.PIPE7_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl3r_net_1\);
    
    \I2.END_TDC5\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_TDC4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_TDC5_net_1\);
    
    \I1.N_237_adt_net_854804_\ : BFR
      port map(A => \I1.N_237\, Y => 
        \I1.N_237_adt_net_854804__net_1\);
    
    \I3.un1_singcyc8_i_0_o2\ : NAND2
      port map(A => \I3.CYCS_net_1\, B => \I3.CYCS1_i_0\, Y => 
        \I3.N_1918\);
    
    \I2.PIPE8_DT_21_il28r\ : OA21TTF
      port map(A => \I2.N_4418\, B => \I2.PIPE7_DTl28r_net_1\, C
         => \I2.PIPE8_DT_21_i_1l28r_net_1\, Y => \I2.N_4399\);
    
    \I2.PIPE1_DT_42_1_IVL22R_1383\ : OAI21FTF
      port map(A => REGl442r, B => 
        \I2.N_3234_adt_net_855648__net_1\, C => 
        \I2.PIPE1_DT_42l22r_adt_net_46757_\, Y => 
        \I2.PIPE1_DT_42l22r_adt_net_46763_\);
    
    \I3.REGMAPl18r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un71_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl18r_net_1\);
    
    \I3.un227_reg_ads_0_a2_3_a3_2\ : OR3
      port map(A => \I3.WRITES_8\, B => \I3.VASl12r_net_1\, C => 
        \I3.N_562\, Y => \I3.un227_reg_ads_2\);
    
    \I3.VDBil14r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_354_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil14r_net_1\);
    
    \I2.un1_tdc_res_45_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl413r, Y => 
        \I2.N_4626_i_0\);
    
    \I2.RAMDT4L11R_2924\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl11r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L11R_441\);
    
    \I2.PIPE5_DT_6_0l28r\ : MUX2L
      port map(A => \I2.PIPE4_DTl28r_net_1\, B => 
        \I2.PIPE5_DT_6l28r_adt_net_53820_\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\, Y => 
        \I2.PIPE5_DT_6l28r\);
    
    \I1.N_145_adt_net_854772_\ : BFR
      port map(A => \I1.N_145\, Y => 
        \I1.N_145_adt_net_854772__net_1\);
    
    \I2.DTO_16_1_IV_0L31R_1064\ : AND2
      port map(A => \I2.DT_SRAMl31r_net_1\, B => 
        \I2.N_182_ADT_NET_1007__385\, Y => 
        \I2.DTO_16_1l31r_adt_net_28246_\);
    
    RAMAD_padl15r : OB33PH
      port map(PAD => RAMAD(15), A => RAMAD_cl15r);
    
    \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_995\ : NOR3
      port map(A => \I2.N_4646_1_ADT_NET_19635__185\, B => 
        \I2.N_4646_1_ADT_NET_19637_RD1__523\, C => 
        \I2.END_EVNT2_403\, Y => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_adt_net_19813_\);
    
    \I2.DTE_21_1_0_IVL31R_1226\ : AND2FT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855192__net_1\, 
        B => \I2.DT_TEMPl31r_net_1\, Y => 
        \I2.DTE_21_1l31r_adt_net_36411_\);
    
    FID_padl11r : OB33PH
      port map(PAD => FID(11), A => FID_cl11r);
    
    \I3.VDBOFFB_59_2366\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl7r_net_1\, Y => 
        \I3.VDBoffb_59_adt_net_161840_\);
    
    \I1.BYTECNT_N2_I_O2_1777\ : AND2
      port map(A => \I1.BYTECNT_I_0_IL1R_435\, B => 
        \I1.BYTECNTL0R_436\, Y => \I1.N_323_adt_net_108906_\);
    
    F_SCK_pad : OB33PH
      port map(PAD => F_SCK, A => \F_SCK_c\);
    
    \I2.PIPE6_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_472_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl18r_net_1\);
    
    \I3.REGMAPl13r_1619\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un54_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL13R_726\);
    
    \I2.STATE5_ns_i_0l0r\ : AOI21FTF
      port map(A => \I2.STATE5l0r_net_1\, B => \I2.N_4338_1\, C
         => \I2.STATE5_ns_i_0_1_il0r\, Y => 
        \I2.STATE5_ns_i_0l0r_net_1\);
    
    \I2.FID_424\ : MUX2H
      port map(A => FID_cl8r, B => \I2.FID_7l8r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        Y => \I2.FID_424_net_1\);
    
    \I1.SBYTE_8_0_a2_i_o2l0r\ : OR2
      port map(A => \I1.sstatel9r_net_1\, B => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854912__net_1\, Y
         => \I1.N_362\);
    
    DTE_padl14r : IOB33PH
      port map(PAD => DTE(14), A => \I2.DTE_1l14r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl14r);
    
    \I2.resyn_0_I2_BITCNT_938\ : MUX2H
      port map(A => \I2.BITCNTl2r_net_1\, B => \I2.N_4323\, S => 
        \I2.BITCNTe\, Y => \I2.BITCNT_938\);
    
    \I2.DTO_16_1_iv_0_a2_4tt_18_m2_0_a2\ : NAND3FTT
      port map(A => \I2.ENDF_net_1\, B => 
        \I2.STATE2l4r_adt_net_855684__net_1\, C => 
        \I2.TEMPF_adt_net_855740__adt_net_855896__net_1\, Y => 
        \I2.DTO_16_1_iv_0_a2_4tt_18_m2_0_a2_net_1\);
    
    \I1.REG_74_2_2L340R_1873\ : NOR2
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720__adt_net_835724_Rd1__net_1\, 
        B => \I1.PAGECNTL6R_836\, Y => 
        \I1.REG_74_2_2_il340r_adt_net_117061_\);
    
    NOE16W_pad : OB33PH
      port map(PAD => NOE16W, A => NOE16W_c);
    
    \I2.OFFSET_37_9l0r\ : MUX2L
      port map(A => \REGl389r\, B => \REGl325r\, S => 
        \I2.PIPE7_DTL27R_85\, Y => \I2.N_699\);
    
    \I3.WRITES\ : DFFC
      port map(CLK => CLK_c, D => \I3.WRITES_23_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.WRITES_8\);
    
    \I1.REG_74_0_ivl308r\ : AO21
      port map(A => \REGl308r\, B => \I1.N_177\, C => 
        \I1.REG_74l308r_adt_net_120180_\, Y => 
        \I1.REG_74l308r_net_1\);
    
    \I1.SBYTE_8_0_il5r\ : OA21
      port map(A => \I1.N_602_i\, B => REGl88r, C => 
        \I1.N_204_adt_net_105924_\, Y => \I1.N_204\);
    
    \I3.UN1_STATE1_13_1_ADT_NET_1351__2803\ : OR3
      port map(A => \I3.un1_STATE1_13_1_adt_net_137890__net_1\, B
         => \I3.un1_STATE1_13_1_adt_net_137896__net_1\, C => 
        \I3.un1_STATE1_13_1_adt_net_137902__net_1\, Y => 
        \I3.UN1_STATE1_13_1_ADT_NET_1351__115\);
    
    \I2.PIPE10_DT_17_I_A3_2L13R_1607\ : OR2
      port map(A => \I2.SUB9_i_0_il13r\, B => \I2.SUB9l12r_net_1\, 
        Y => \I2.N_3822_adt_net_64757_\);
    
    \I3.VDBOFFB_30_IV_0L7R_2363\ : OR2
      port map(A => \I3.VDBoffb_30l7r_adt_net_161791_\, B => 
        \I3.VDBoffb_30l7r_adt_net_161792_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161797_\);
    
    \I2.OFFSET_37_15l7r\ : MUX2L
      port map(A => \REGl236r\, B => \REGl172r\, S => 
        \I2.PIPE7_DTL27R_67\, Y => \I2.N_754\);
    
    \I3.PULSEl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_331_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl1r);
    
    \I3.un1_REGMAP_34_0_a2_0_a2_746\ : NOR2FT
      port map(A => \I3.UN1_REGMAP_30_375\, B => 
        \I3.N_178_ADT_NET_1360__127\, Y => \I3.UN1_REGMAP_34_124\);
    
    \I2.DTE_21_1_IVL11R_1296\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, 
        B => \I2.DT_TEMPl11r_net_1\, C => 
        \I2.DTE_21_1l11r_adt_net_38399_\, Y => 
        \I2.DTE_21_1l11r_adt_net_38414_\);
    
    \I1.COMMAND_52\ : MUX2L
      port map(A => 
        \PULSEl0r_adt_net_854532__adt_net_855544__net_1\, B => 
        \I1.COMMAND_net_1\, S => \I1.N_1384\, Y => 
        \I1.COMMAND_52_0\);
    
    \I0.COM_SERSi_1454\ : DFFC
      port map(CLK => CLK_c, D => \I0.COM_SERF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => COM_SERS_561);
    
    \I1.REG_74_1_i_a2_a0l404r\ : OR2FT
      port map(A => \I1.REG_74_1_i_a2_a0_2l404r\, B => 
        \I1.N_1367_i_adt_net_112072_\, Y => \I1.N_1367_i\);
    
    \I2.DTO_16_1_IV_0_0L18R_1129\ : AO21
      port map(A => \I2.N_197_152\, B => 
        \I2.DTO_16_1l18r_adt_net_756__net_1\, C => 
        \I2.DTO_16_1l18r_adt_net_31333_\, Y => 
        \I2.DTO_16_1l18r_adt_net_31346_\);
    
    \I2.DTE_21_1_IV_0L20R_1259\ : AND2FT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_288\, B => 
        \I2.DT_SRAMl20r_net_1\, Y => 
        \I2.DTE_21_1l20r_adt_net_37605_\);
    
    \I3.TCNT2_394\ : MUX2H
      port map(A => \I3.TCNT2_i_0_il2r_net_1\, B => 
        \I3.TCNT2_n2_net_1\, S => TICKL0R_558, Y => 
        \I3.TCNT2_394_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I46_Y_1676\ : AND2FT
      port map(A => \I2.LSRAM_OUTl16r\, B => 
        \I2.PIPE7_DTl16r_net_1\, Y => \I2.N296_0_adt_net_86403_\);
    
    \I2.REG_1_n15_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => REGl47r, Y => \I2.REG_1_n15_0_net_1\);
    
    \I2.EVNT_WORD_716\ : MUX2H
      port map(A => \I2.EVNT_WORDl3r_net_1\, B => \I2.I_13_1\, S
         => \I2.N_2864_0_adt_net_854276__net_1\, Y => 
        \I2.EVNT_WORD_716_net_1\);
    
    \I2.ROFFSET_224\ : NAND2FT
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855704__net_1\, B => 
        \I2.ROFFSETl0r_net_1\, Y => \I2.N_1355\);
    
    \I2.TRGSERVl0r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.DWACT_ADD_CI_0_partial_sum_1l0r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGSERVl0r_net_1\);
    
    \I2.PIPE4_DTL7R_2965\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL7R_482\);
    
    \I3.VDBi_40_0l5r\ : OAI21TTF
      port map(A => \I3.N_1772_adt_net_143698_\, B => 
        \I3.N_1772_adt_net_143704_\, C => 
        \I3.VDBi_40l5r_adt_net_143744_\, Y => \I3.VDBi_40l5r\);
    
    \I1.REG_74_0_ivl283r\ : AO21
      port map(A => \REGl283r\, B => \I1.N_153\, C => 
        \I1.REG_74l283r_adt_net_122463_\, Y => \I1.REG_74l283r\);
    
    \I3.VDBi_57_iv_0_0_a2_13l7r\ : NOR3FTT
      port map(A => \I3.REGMAPl17r_adt_net_854296__net_1\, B => 
        \I3.N_2014\, C => \I3.REGMAPL55R_782\, Y => \I3.N_2046\);
    
    \I1.REG_1_67\ : MUX2H
      port map(A => \REGl166r\, B => \I1.REG_74l166r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, Y => 
        \I1.REG_1_67_net_1\);
    
    \I2.PIPE7_DTl12r_1586\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL12R_693\);
    
    \I3.VDBi_57_iv_0_0l6r\ : OR3
      port map(A => \I3.VDBi_57l6r_adt_net_143394_\, B => 
        \I3.VDBi_57l6r_adt_net_143402_\, C => 
        \I3.VDBi_57l6r_adt_net_143403_\, Y => \I3.VDBi_57l6r\);
    
    \I1.REG_2_sqmuxa_adt_net_855392_\ : BFR
      port map(A => \I1.REG_2_sqmuxa\, Y => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\);
    
    \I3.un235_reg_ads_0_a2_2_a3\ : NOR3
      port map(A => \I3.N_547\, B => \I3.N_558\, C => \I3.N_634\, 
        Y => \I3.un235_reg_ads_0_a2_2_a3_net_1\);
    
    \I3.VDBil31r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_371_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil31r_net_1\);
    
    \I2.OFFSET_37_12l3r\ : MUX2L
      port map(A => \REGl344r\, B => \I2.N_718\, S => 
        \I2.PIPE7_DTL26R_358\, Y => \I2.N_726\);
    
    \I1.N_50_0_ADT_NET_1409__2749\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__200\, B => 
        \I1.N_50_0_ADT_NET_109751__258\, Y => 
        \I1.N_50_0_ADT_NET_1409__22\);
    
    \I3.TCNT2_396\ : XOR2
      port map(A => \I3.TCNT2_i_0_il0r_net_1\, B => TICKL0R_558, 
        Y => \I3.TCNT2_396_net_1\);
    
    \I1.REG_74_0_ivl190r\ : AO21
      port map(A => \REGl190r\, B => \I1.N_65\, C => 
        \I1.REG_74l190r_adt_net_131441_\, Y => \I1.REG_74l190r\);
    
    \I3.TCNT2_n5\ : XOR2
      port map(A => \I3.TCNT2l5r_net_1\, B => \I3.TCNT2_c4\, Y
         => \I3.TCNT2_n5_net_1\);
    
    \I2.SUB9_581\ : MUX2H
      port map(A => \I2.SUB9_i_0_il13r\, B => \I2.SUB9_1l13r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_581_net_1\);
    
    \I1.REG_9_sqmuxa_adt_net_854728_\ : BFR
      port map(A => \I1.REG_9_sqmuxa\, Y => 
        \I1.REG_9_sqmuxa_adt_net_854728__net_1\);
    
    DTO_padl4r : IOB33PH
      port map(PAD => DTO(4), A => \I2.DTO_1l4r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl4r);
    
    \I2.SUB9l14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_582_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l14r_net_1\);
    
    \I2.CRC32_12_0_0_x2l26r\ : XOR2FT
      port map(A => \I2.CRC32l26r_net_1\, B => \I2.N_4271_i_i\, Y
         => \I2.N_127_i_0_i_0\);
    
    \I2.DTE_1_860\ : MUX2L
      port map(A => \I2.DTE_1l22r_Rd1__net_1\, B => 
        \I2.DTE_21_1l22r_Rd1_\, S => 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\, Y => 
        \I2.DTE_1l22r\);
    
    \I1.REG_74_0_IVL375R_1824\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l375r_adt_net_112915_\);
    
    \I2.ROFFSET_c1\ : NAND2
      port map(A => \I2.ROFFSETl0r_net_1\, B => 
        \I2.ROFFSETl1r_net_1\, Y => \I2.ROFFSET_c1_net_1\);
    
    \I2.END_EVNT2_1141\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT1_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT2_403\);
    
    \I2.DTO_16_1_ivl10r\ : OR2
      port map(A => \I2.DTO_16_1l10r_adt_net_33065_\, B => 
        \I2.DTO_16_1l10r_adt_net_33066_\, Y => \I2.DTO_16_1l10r\);
    
    \I1.N_341_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_341_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_341_Rd1__net_1\);
    
    \I1.REG_1_86\ : MUX2H
      port map(A => \REGl185r\, B => \I1.REG_74l185r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, Y => 
        \I1.REG_1_86_net_1\);
    
    \I1.N_113_adt_net_126306_\ : OAI21TTF
      port map(A => \I1.REG_74_1_396_m7_i_3\, B => 
        \I1.REG_74_8_308_N_6_i\, C => 
        \I1.N_113_adt_net_126301__net_1\, Y => 
        \I1.N_113_adt_net_126306__net_1\);
    
    \I1.REG_74_12_348_M9_I_1855\ : NOR2FT
      port map(A => \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, 
        B => \I1.PAGECNTl5r_net_1\, Y => 
        \I1.REG_74_12_348_m9_i_adt_net_115429_\);
    
    \I3.TCNT3_i_0_il2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT3_377_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT3_i_0_il2r_net_1\);
    
    \I2.STATEel3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATEe_ns_il1r_net_1\, CLR
         => \I2.STATEe_i_0l0r_net_1\, Q => \I2.STATEe_ipl3r\);
    
    \I2.DTE_21_1l16r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l16r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l16r_Rd1__net_1\);
    
    \I2.N507_adt_net_56251_\ : AO21
      port map(A => \I2.PIPE4_DTL12R_511\, B => 
        \I2.PIPE4_DTL14R_639\, C => \I2.RAMDT4L5R_814\, Y => 
        \I2.N507_adt_net_56251__net_1\);
    
    \I3.REGMAPl9r_adt_net_854324_\ : BFR
      port map(A => \I3.REGMAPl9r_adt_net_854328__net_1\, Y => 
        \I3.REGMAPl9r_adt_net_854324__net_1\);
    
    REGl353r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_254_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl353r\);
    
    \I2.ADO_3l12r\ : MUX2H
      port map(A => \I2.RPAGEl12r\, B => \I2.WPAGEl12r_net_1\, S
         => NOESRAME_c, Y => \I2.ADO_3l12r_net_1\);
    
    DTE_padl27r : IOB33PH
      port map(PAD => DTE(27), A => \I2.DTE_1l27r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl27r);
    
    \I2.MIC_ERR_REGSl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_358_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl29r_net_1\);
    
    \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832_\ : BFR
      port map(A => \I2.un1_STATE3_10_1_adt_net_999__net_1\, Y
         => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\);
    
    \I2.N_4547_1_adt_net_1209_\ : NAND2
      port map(A => \I2.PIPE4_DTl31r_net_1\, B => REGl0r, Y => 
        \I2.N_4547_1_adt_net_1209__net_1\);
    
    SP5_pad : OB33PH
      port map(PAD => SP5, A => \GND\);
    
    \I2.un1_tdc_res_25_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl417r, Y => 
        \I2.N_4606_i_0\);
    
    \I2.PIPE8_DT_16_0l17r\ : MUX2H
      port map(A => \I2.PIPE8_DTl17r_net_1\, B => 
        \I2.PIPE7_DTl17r_net_1\, S => 
        \I2.N_565_0_adt_net_855736__net_1\, Y => \I2.N_583\);
    
    \I2.OFFSET_37_10l3r\ : MUX2L
      port map(A => \I2.N_702\, B => \I2.N_694\, S => 
        \I2.PIPE7_DTL26R_353\, Y => \I2.N_710\);
    
    \I2.BNCID_VECTror_10_tz\ : AOI21
      port map(A => \I2.BNCID_VECTra14_1_net_1\, B => 
        \I2.BNCID_VECTro_6\, C => \I2.BNCID_VECTria_7_0_net_1\, Y
         => \I2.BNCID_VECTror_10_tz_adt_net_48171_\);
    
    \I2.LSRAM_INl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_388_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl4r_net_1\);
    
    \I2.EVNT_WORD_725\ : MUX2H
      port map(A => \I2.EVNT_WORDl12r_net_1\, B => \I2.I_73\, S
         => \I2.N_2864_0_adt_net_854268__net_1\, Y => 
        \I2.EVNT_WORD_725_net_1\);
    
    \I5.REG_1l418r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_31_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl418r);
    
    \I2.BNCID_VECT_tile_I_6_0\ : XOR2
      port map(A => \I2.TRGSERVl0r_net_1\, B => 
        \I2.WADDR_REG1l0r\, Y => \I2.I_6_0_i_0_i\);
    
    \I2.DTE_21_1_IV_0L12R_1290\ : AND2
      port map(A => \I2.DTE_1l12r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1l12r_adt_net_38283_\);
    
    \I3.VDBm_0l24r\ : MUX2L
      port map(A => \I3.PIPEAl24r_net_1\, B => 
        \I3.PIPEBl24r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_166\);
    
    \I3.N_1917_adt_net_855336_\ : BFR
      port map(A => \I3.N_1917\, Y => 
        \I3.N_1917_adt_net_855336__net_1\);
    
    \I2.REG_1_c8_i_a2_0\ : AND3FFT
      port map(A => REGl39r, B => REGl40r, C => \I2.N_126\, Y => 
        \I2.N_129\);
    
    \I2.PIPE8_DT_21l3r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl3r\, B => \I2.N_569\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l3r_net_1\);
    
    \I2.DTE_21_1_IVL11R_1298\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l11r\, C
         => \I2.DTE_21_1l11r_adt_net_38416_\, Y => 
        \I2.DTE_21_1l11r_adt_net_38417_\);
    
    \I5.SDAout_12_iv_0_o4\ : AO21FTT
      port map(A => \I5.N_64\, B => \I5.COMMANDl0r_net_1\, C => 
        \I5.N_71_adt_net_9287_\, Y => \I5.N_71\);
    
    \I2.L2TYPEl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_595_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl6r_net_1\);
    
    \I2.EVNT_NUM_c5\ : AND2
      port map(A => \I2.EVNT_NUMl5r_net_1\, B => 
        \I2.EVNT_NUM_c4_net_1\, Y => \I2.EVNT_NUM_c5_net_1\);
    
    \I2.LSRAM_IN_405\ : MUX2L
      port map(A => \I2.PIPE5_DTl21r_net_1\, B => 
        \I2.LSRAM_INl21r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_405_net_1\);
    
    REGl214r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_115_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl214r\);
    
    AMB_padl5r : IB33
      port map(PAD => AMB(5), Y => AMB_c_i_0_il5r);
    
    \I3.PIPEA1_12l8r\ : AND2
      port map(A => DPR_cl8r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854508__net_1\, Y => 
        \I3.PIPEA1_12l8r_net_1\);
    
    \I1.REG_74_0_ivl171r\ : AO21
      port map(A => \REGl171r\, B => \I1.N_41\, C => 
        \I1.REG_74l171r_adt_net_133149_\, Y => \I1.REG_74l171r\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854628_\ : BFR
      port map(A => \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\, Y
         => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854628__net_1\);
    
    \I2.DTO_16_1_iv_0_o2_0_i_o2l21r\ : OAI21FTF
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.N_182_ADT_NET_1007__155\, Y => \I2.N_197\);
    
    \I2.STOP_RDSRAM_453_i_adt_net_1077_\ : AO21
      port map(A => \I2.STATE3l3r_net_1\, B => \I2.N_145\, C => 
        \I2.STOP_RDSRAM_net_1\, Y => 
        \I2.STOP_RDSRAM_453_i_adt_net_1077__net_1\);
    
    \I2.N_182_ADT_NET_1007__2915\ : OR2
      port map(A => \I2.STATE2l0r_net_1\, B => 
        \I2.STATE2_nsl2r_adt_net_24911_\, Y => 
        \I2.N_182_ADT_NET_1007__386\);
    
    \I1.ISI_0_sqmuxa_1_0_i_o2_0\ : OR2
      port map(A => \I1.sstatel3r_net_1\, B => 
        \I1.sstatel6r_net_1\, Y => \I1.N_366\);
    
    \I2.PIPE4_DTl15r_1530\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl15r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL15R_637\);
    
    \I2.MAJORITY_REG_IL5R_1019\ : AOI21
      port map(A => \I2.MIC_REG2_i_0_il5r_net_1\, B => 
        \I2.MIC_REG1l5r_net_1\, C => \I2.MIC_REG3l5r_net_1\, Y
         => \I2.N_4431_adt_net_22416_\);
    
    \I3.VDBm_il7r\ : MUX2L
      port map(A => \I3.VDBil7r_net_1\, B => \I3.N_129\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.N_11\);
    
    \I2.PIPE5_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_699_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl23r_net_1\);
    
    \I5.SBYTEl0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_65_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl0r_net_1\);
    
    \I5.REG_1l427r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_40_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl427r);
    
    \I2.DT_SRAM_0_i_m2l2r\ : MUX2L
      port map(A => \I2.PIPE10_DTl2r_net_1\, B => 
        \I2.PIPE5_DTl2r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854204__net_1\, Y => 
        \I2.N_4191\);
    
    \I3.PIPEAl18r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_249_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl18r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I144_Y_2656\ : OR2
      port map(A => \I2.N516_adt_net_87903__net_1\, B => 
        \I2.N326_0\, Y => \I2.N510_adt_net_220925_\);
    
    \I2.PIPE1_DT_42_1_IVL6R_1486\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl2r\, Y => 
        \I2.PIPE1_DT_42l6r_adt_net_50930_\);
    
    \I5.DATAl13r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l13r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl130r);
    
    \I2.FID_7_0_IVL0R_1734\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl48r, C => 
        \I2.FID_7l0r_adt_net_93569_\, Y => 
        \I2.FID_7l0r_adt_net_93577_\);
    
    \I3.REG_1_155\ : MUX2L
      port map(A => VDB_inl6r, B => REGl54r, S => 
        \I3.N_1935_adt_net_855332__net_1\, Y => \I3.REG_1_155_0\);
    
    \I3.VDBOFFA_31_IV_0L7R_2504\ : AO21
      port map(A => \REGl268r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        C => \I3.VDBoffa_31l7r_adt_net_163284_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163313_\);
    
    \I2.PIPE8_DT_538\ : MUX2L
      port map(A => \I2.PIPE8_DTl10r_net_1\, B => 
        \I2.PIPE8_DT_21l10r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_538_net_1\);
    
    \I3.REG_1_265\ : MUX2H
      port map(A => REGl84r, B => \I3.N_1630\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_265_0\);
    
    \I2.L2SERVl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_922_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEl12r\);
    
    \I1.REG_74_0_ivl319r\ : AO21
      port map(A => \REGl319r\, B => \I1.N_193\, C => 
        \I1.REG_74l319r_adt_net_119131_\, Y => \I1.REG_74l319r\);
    
    \I3.VDBi_55l12r\ : MUX2H
      port map(A => \I3.VDBil12r_net_1\, B => 
        \I3.RAMDTSl12r_net_1\, S => 
        \I3.N_57_i_0_0_adt_net_854692__net_1\, Y => 
        \I3.VDBi_55l12r_net_1\);
    
    \I4.STATE1l0r\ : DFFC
      port map(CLK => CLK_c, D => \I4.STATE1_nsl2r\, CLR => 
        CLEAR_STAT_i_0, Q => \I4.STATE1l0r_net_1\);
    
    \I2.un6_tdcgdb1_1\ : XOR2
      port map(A => \I2.TDCl1r_net_1\, B => \I2.TDCDBSl25r_net_1\, 
        Y => \I2.un6_tdcgdb1_1_net_1\);
    
    \I2.G_EVNT_NUM_n5_i_0_a2\ : NOR2FT
      port map(A => \I2.N_4669_adt_net_855052__net_1\, B => 
        \I2.G_EVNT_NUMl5r_net_1\, Y => \I2.N_319\);
    
    \I2.DT_SRAM_0_i_m2l13r\ : MUX2L
      port map(A => \I2.PIPE10_DTl13r_net_1\, B => 
        \I2.PIPE5_DTl13r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854224__net_1\, Y => 
        \I2.N_4046\);
    
    MTDCRESB_pad : OB33PH
      port map(PAD => MTDCRESB, A => MTDCRESB_c);
    
    \I2.FID_7_0_ivl31r\ : AO21
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOS_i_il31r\, C
         => \I2.FID_7l31r_adt_net_18465_\, Y => \I2.FID_7l31r\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I138_Y_0_1579\ : NOR3FTT
      port map(A => \I2.N_112_2\, B => 
        \I2.ADD_21x21_fast_I138_Y_0_0\, C => 
        \I2.N_114_adt_net_275800_\, Y => 
        \I2.N513_i_adt_net_58503_\);
    
    \I3.UN131_REG_ADS_0_A2_1_A2_2649\ : OR2FT
      port map(A => \I3.VASl4r_net_1\, B => \I3.VASl1r_net_1\, Y
         => \I3.N_586_adt_net_165970_\);
    
    \I3.REG_1_283\ : MUX2L
      port map(A => VDB_inl1r, B => REGl102r, S => 
        \I3.N_318_adt_net_855888__net_1\, Y => \I3.REG_1_283_0\);
    
    \I3.VDBi_40_0_i_m2l11r\ : MUX2L
      port map(A => REGl429r, B => REGl445r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_1856\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I180_UN1_Y_2669\ : AND2
      port map(A => \I2.N305_0\, B => 
        \I2.N258_0_adt_net_854936__net_1\, Y => 
        \I2.I180_un1_Y_adt_net_309337_\);
    
    \I2.OFFSET_561\ : MUX2L
      port map(A => \I2.OFFSETl1r_net_1\, B => \I2.OFFSET_37l1r\, 
        S => \I2.un1_NWPIPE7_2_net_1\, Y => \I2.OFFSET_561_net_1\);
    
    \I1.REG_74_0_IV_0_0_O2L253R_1964\ : OR3
      port map(A => \I1.N_374\, B => \I1.N_395\, C => \I1.N_592\, 
        Y => \I1.N_658_adt_net_124758_\);
    
    \I1.REG_1_304\ : MUX2H
      port map(A => \REGl403r\, B => \I1.REG_74l403r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\, Y => 
        \I1.REG_1_304_net_1\);
    
    \I2.L2TYPE_4_i_o2l3r\ : AND2FT
      port map(A => \I2.N_4454\, B => \I2.N_4461\, Y => 
        \I2.N_4465\);
    
    \I3.VDBm_0l3r\ : MUX2L
      port map(A => \I3.PIPEAl3r_net_1\, B => \I3.PIPEBl3r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_145\);
    
    \I2.REG_1_n9\ : XOR2FT
      port map(A => \I2.N_3837_i_0\, B => \I2.REG_1_n9_0_net_1\, 
        Y => \I2.REG_1_n9_net_1\);
    
    \I1.BYTECNT_313\ : MUX2H
      port map(A => \I1.BYTECNT_i_0_il1r_net_1\, B => \I1.N_1161\, 
        S => \I1.N_1383\, Y => \I1.BYTECNT_313_net_1\);
    
    \I3.VADm_0_a3l28r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl28r_net_1\, Y => \I3.VADml28r\);
    
    \I2.STATE4_ns_i_0_o2l1r\ : NAND2
      port map(A => \I2.L1AF2_net_1\, B => \I2.L1AF3_i_0\, Y => 
        \I2.N_4464\);
    
    \I2.PIPE8_DT_16_0l7r\ : MUX2H
      port map(A => \I2.PIPE8_DTl7r_net_1\, B => 
        \I2.PIPE7_DTl7r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_573\);
    
    \I2.DTO_9_IVL7R_1183\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        B => \I2.DTE_2_1l7r_net_1\, Y => 
        \I2.DTO_9l7r_adt_net_33660_\);
    
    \I2.un7_bnc_id_1_I_20\ : XOR2
      port map(A => \I2.N_37\, B => \I2.BNC_IDl4r_net_1\, Y => 
        \I2.I_20_0\);
    
    \I2.SUB9_1_ADD_18x18_fast_I109_Y\ : AND2FT
      port map(A => \I2.I109_un1_Y\, B => 
        \I2.N439_i_adt_net_71055_\, Y => \I2.N439_i\);
    
    TDCDA_padl27r : IB33
      port map(PAD => TDCDA(27), Y => TDCDA_cl27r);
    
    \I2.PIPE1_DT_42_1_IVL17R_1409\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\, B => 
        \I2.PIPE1_DT_30l17r_net_1\, C => 
        \I2.PIPE1_DT_42l17r_adt_net_47635_\, Y => 
        \I2.PIPE1_DT_42l17r_adt_net_47650_\);
    
    \I2.LEAD_FLAG6l6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_643_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl6r);
    
    \I2.un1_NWPIPE7_2\ : OR2FT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855156__net_1\, B
         => \I2.un1_NWPIPE7_2_adt_net_73606_\, Y => 
        \I2.un1_NWPIPE7_2_net_1\);
    
    \I2.DTO_9_iv_0l31r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl31r_net_1\, 
        C => \I2.DTO_9l31r_adt_net_27894_\, Y => \I2.DTO_9l31r\);
    
    \I2.PIPE1_DT_42_1_IVL13R_1444\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl9r\, Y => 
        \I2.PIPE1_DT_42l13r_adt_net_49201_\);
    
    \I3.NOEDTKi\ : DFFS
      port map(CLK => CLK_c, D => \I3.NOEDTKi_111_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => NOEDTK_c);
    
    \I3.un1_STATE2_15_1_adt_net_147708_\ : OR3
      port map(A => \I3.N_1879\, B => 
        \I3.un1_STATE2_15_1_adt_net_147701__net_1\, C => 
        \I3.STATE2l3r_net_1\, Y => 
        \I3.un1_STATE2_15_1_adt_net_147708__net_1\);
    
    \I1.REG_74_1_380_m8_i_0_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.REG_74_1_380_m8_i_0_Ra1_\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.REG_74_1_380_m8_i_0_Rd1__net_1\);
    
    \I2.DTE_21_1_iv_0_18_N_8_i_0_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1_iv_0_18_N_8_i_0\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_Rd1__net_1\);
    
    \I1.REG_74_0_ivl301r\ : AO21
      port map(A => \REGl301r\, B => \I1.N_177\, C => 
        \I1.REG_74l301r_adt_net_120782_\, Y => \I1.REG_74l301r\);
    
    \I2.PIPE4_DTL10R_2959\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL10R_476\);
    
    \I2.DTO_16_1_IVL22R_1107\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.G_EVNT_NUMl6r_net_1\, Y
         => \I2.DTO_16_1l22r_adt_net_30352_\);
    
    \I1.SBYTE_61\ : MUX2L
      port map(A => \FBOUTl3r\, B => \I1.N_202\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_61_net_1\);
    
    \I1.REG_1_230\ : MUX2H
      port map(A => \REGl329r\, B => \I1.REG_74l329r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y => 
        \I1.REG_1_230_net_1\);
    
    \I3.REG_1l68r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_169_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl68r);
    
    RAMDT_padl10r : IOB33PH
      port map(PAD => RAMDT(10), A => \I1.RAMDT_SPI_1l3r_net_1\, 
        EN => \I1.RAMDT_SPI_E_0\, Y => RAMDT_inl10r);
    
    \I2.L2ARRl1r_1496\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_943_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRL1R_603\);
    
    \I2.END_EVNT7\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT6_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT7_net_1\);
    
    \I2.DTO_16_1_IV_0_0L6R_1193\ : AO21
      port map(A => \I2.N_197\, B => \I2.DT_SRAMl6r_net_1\, C => 
        \I2.DTO_16_1l6r_adt_net_33912_\, Y => 
        \I2.DTO_16_1l6r_adt_net_33922_\);
    
    \I1.REG_74_0_iv_i_a2l199r\ : AO21
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_1338_adt_net_130619_\, Y => \I1.N_1338\);
    
    \I1.REG_74_0_IVL341R_1872\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l341r_adt_net_116928_\);
    
    \I1.REG_74L220R_2010\ : AND3FFT
      port map(A => \I1.REG_74_1_a0_0l228r_adt_net_854832__net_1\, 
        B => \I1.REG_74_12_220_m9_i_a6_0\, C => 
        \I1.N_89_adt_net_128729_\, Y => \I1.N_89_adt_net_128731_\);
    
    \I2.PIPE1_DT_746\ : MUX2L
      port map(A => \I2.PIPE1_DTl19r_net_1\, B => 
        \I2.PIPE1_DT_42l19r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854572__net_1\, 
        Y => \I2.PIPE1_DT_746_net_1\);
    
    \I2.OFFSET_37_25l7r\ : MUX2L
      port map(A => \REGl260r\, B => \REGl196r\, S => 
        \I2.PIPE7_DTL27R_87\, Y => \I2.N_834\);
    
    \I2.DTE_21_1_0_IV_0_0L29R_1233\ : AO21
      port map(A => \I2.STATE2L3R_440\, B => \I2.N_4159\, C => 
        \I2.DTE_21_1l29r_adt_net_36650_\, Y => 
        \I2.DTE_21_1l29r_adt_net_36651_\);
    
    \I2.EVNT_NUM_n5\ : NOR2
      port map(A => EV_RES_c, B => \I2.EVNT_NUM_n5_tz_i\, Y => 
        \I2.EVNT_NUM_n5_net_1\);
    
    \I1.REG_1_105\ : MUX2H
      port map(A => \REGl204r\, B => \I1.N_1343\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_105_net_1\);
    
    VAD_padl27r : OTB33PH
      port map(PAD => VAD(27), A => \I3.VADml27r\, EN => 
        NOEAD_c_i_0);
    
    \I3.RAMAD_VMEl16r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_40_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl16r);
    
    \I5.AIR_START_16\ : OR2
      port map(A => \I5.N_463\, B => \TICKl3r\, Y => 
        \I5.AIR_START_16_net_1\);
    
    \I3.REGMAPL55R_3027\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un224_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL55R_781\);
    
    \I2.CRC32_12_0_0_m2l24r\ : MUX2H
      port map(A => \I2.N_4194\, B => \I2.DT_TEMPl24r_net_1\, S
         => \I2.N_4667_1_adt_net_1046__adt_net_854428__net_1\, Y
         => \I2.N_4270_i_i\);
    
    \I2.CRC32_1_sqmuxa_1_i_o2_925\ : OR2
      port map(A => \I2.STATE2L4R_291\, B => \I2.STATE2L3R_437\, 
        Y => \I2.N_4261_303\);
    
    \I2.OFFSET_37_12l5r\ : MUX2L
      port map(A => \REGl346r\, B => \I2.N_720\, S => 
        \I2.PIPE7_DTL26R_357\, Y => \I2.N_728\);
    
    \I3.un15_tcnt4\ : AND2
      port map(A => \I3.un12_tcnt3_net_1\, B => 
        \I3.un15_tcnt4_adt_net_165652_\, Y => 
        \I3.un15_tcnt4_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I136_Y_0_o2_m4_1\ : 
        AO21TTF
      port map(A => \I2.N_2358_tz_tz\, B => 
        \I2.N_152_i_0_adt_net_502546_\, C => 
        \I2.N_163_0_adt_net_55087_\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_1_i\);
    
    \I1.REG_15_sqmuxa_adt_net_109461_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => 
        \I1.REG_15_sqmuxa_adt_net_109461_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.REG_15_sqmuxa_adt_net_109461_Rd1__net_1\);
    
    \I1.REG_1_107\ : MUX2H
      port map(A => \REGl206r\, B => \I1.N_282\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_107_net_1\);
    
    \I5.COMMANDl8r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_45_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl8r_net_1\);
    
    \I3.VDBml11r\ : MUX2L
      port map(A => \I3.VDBil11r_net_1\, B => \I3.N_153\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml11r_net_1\);
    
    \I3.VDBoff_122\ : MUX2L
      port map(A => \I3.VDBoffl6r_net_1\, B => \I3.N_79\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_122_net_1\);
    
    \I3.UN1_REGMAP_34_5_0_A2_I_O2_I_A2_2_O2_2087\ : NOR2
      port map(A => \I3.REGMAP_I_0_IL45R_452\, B => 
        \I3.REGMAPL44R_451\, Y => \I3.N_2086_adt_net_134541_\);
    
    \I2.LSRAM_WADDRl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_WADDR_381_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_WADDRl0r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I10_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L5R_815\, B => 
        \I2.PIPE4_DTL10R_791\, Y => \I2.N_59\);
    
    \I2.OFFSET_37_22l3r\ : MUX2L
      port map(A => \REGl240r\, B => \REGl176r\, S => 
        \I2.PIPE7_DTL27R_82\, Y => \I2.N_806\);
    
    \I2.PIPE10_DT_17_I_A3_2L13R_1608\ : OR2
      port map(A => \I2.SUB9_i_0_il11r\, B => \I2.SUB9l10r_net_1\, 
        Y => \I2.N_3822_adt_net_64759_\);
    
    \I1.REG_1_233\ : MUX2H
      port map(A => \REGl332r\, B => \I1.REG_74l332r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y
         => \I1.REG_1_233_net_1\);
    
    \I3.REG_1l71r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_172_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl71r);
    
    \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__2826\ : OAI21TTF
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096__net_1\, B
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        C => \I2.FIRST_TDC_1_sqmuxa_net_1\, Y => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__170\);
    
    \I2.TDCDASl19r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl19r, Q => 
        \I2.TDCDASl19r_net_1\);
    
    \I3.VDBi_29l8r\ : MUX2L
      port map(A => \I3.REGl99r\, B => \I3.VDBi_20l8r\, S => 
        \I3.REGMAPl14r_net_1\, Y => \I3.VDBi_29l8r_net_1\);
    
    \I2.PIPE1_DT_744\ : MUX2L
      port map(A => \I2.PIPE1_DTl17r_net_1\, B => 
        \I2.PIPE1_DT_42l17r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854572__net_1\, 
        Y => \I2.PIPE1_DT_744_net_1\);
    
    \I3.un1_STATE2_13_adt_net_1333_\ : OR3
      port map(A => \I3.N_12180_i\, B => 
        \I3.un1_STATE2_13_adt_net_150841__net_1\, C => 
        \I3.un1_STATE2_13_adt_net_150833__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__net_1\);
    
    \I2.DTO_16_1_iv_0_o2_0_i_o2l21r_774\ : OAI21FTF
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.N_182_ADT_NET_1007__155\, Y => \I2.N_197_152\);
    
    \I2.REG_1_n14\ : XOR2FT
      port map(A => \I2.N_3842_i_0\, B => \I2.REG_1_n14_0_net_1\, 
        Y => \I2.REG_1_n14_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL4R_1501\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, B => 
        \I2.PIPE1_DT_30l4r_net_1\, C => 
        \I2.PIPE1_DT_42l4r_adt_net_51418_\, Y => 
        \I2.PIPE1_DT_42l4r_adt_net_51434_\);
    
    \I2.LSRAM_WADDRl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_WADDR_383_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_WADDRl2r_net_1\);
    
    \I3.TCNTl1r_1167\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_383_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTL1R_429\);
    
    \I3.REG_1_168\ : MUX2L
      port map(A => VDB_inl19r, B => REGl67r, S => 
        \I3.N_1935_adt_net_855324__net_1\, Y => \I3.REG_1_168_0\);
    
    \I3.REGMAPL26R_2985\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un111_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL26R_532\);
    
    \I3.VDBOFFA_31_IV_0L0R_2625\ : AO21
      port map(A => \REGl197r\, B => \I3.REGMAPl22r_net_1\, C => 
        \I3.VDBoffa_31l0r_adt_net_164594_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164638_\);
    
    \I2.NWPIPE10\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE9_0_7\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE10_net_1\);
    
    \I2.FIDl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_436\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl20r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I152_Y_0\ : AO21
      port map(A => \I2.N498_0_adt_net_598283_\, B => 
        \I2.N498_0_adt_net_598321_\, C => 
        \I2.N498_0_adt_net_56940_\, Y => \I2.N498_0\);
    
    \I5.un1_SENS_ADDR_1_I_15\ : AND2
      port map(A => \I5.DWACT_ADD_CI_0_TMPl0r\, B => 
        \I5.SENS_ADDRl1r_net_1\, Y => 
        \I5.DWACT_ADD_CI_0_g_array_1l0r\);
    
    \I5.CHAIN_SELECT\ : DFFC
      port map(CLK => CLK_c, D => \I5.CHAIN_SELECT_11_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.CHAIN_SELECT_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I9_G0N_0_o3\ : AND2
      port map(A => \I2.RAMDT4L5R_817\, B => 
        \I2.PIPE4_DTl9r_net_1\, Y => \I2.N_16\);
    
    \I3.VDBI_57_IV_0_0L7R_2229\ : OA21TTF
      port map(A => \I3.VDBi_57l7r_adt_net_143036__net_1\, B => 
        \I3.VDBi_57l7r_adt_net_143037__net_1\, C => 
        \I3.N_1905_1_adt_net_855384__net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_143103_\);
    
    \I1.REG_74_0_iv_0_0l246r\ : AO21
      port map(A => \REGl246r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l246r_adt_net_126121_\, Y => \I1.REG_74l246r\);
    
    \I2.OFFSET_37_2l3r\ : MUX2L
      port map(A => \REGl384r\, B => \REGl320r\, S => 
        \I2.PIPE7_DTL27R_71\, Y => \I2.N_646\);
    
    \I3.PIPEAl0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_231_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl0r_net_1\);
    
    \I2.PIPE6_DT_484\ : MUX2H
      port map(A => \I2.PIPE5_DTl30r_net_1\, B => 
        \I2.PIPE6_DTl30r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_484_net_1\);
    
    \I2.ROFFSET_c8\ : NOR2FT
      port map(A => \I2.ROFFSETl8r_net_1\, B => 
        \I2.ROFFSET_c7_net_1\, Y => \I2.ROFFSET_c8_net_1\);
    
    \I2.un1_tdc_res_31_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl414r, Y => 
        \I2.N_4612_i_0\);
    
    \I3.PIPEA1_327\ : MUX2L
      port map(A => \I3.PIPEA1l29r_net_1\, B => 
        \I3.PIPEA1_12l29r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, Y => 
        \I3.PIPEA1_327_net_1\);
    
    \I2.OFFSET_37_20l3r\ : MUX2L
      port map(A => \I2.N_782\, B => \I2.N_774\, S => 
        \I2.PIPE7_DTL26R_358\, Y => \I2.N_790\);
    
    \I2.un21_pipe5_dt_0\ : XOR2
      port map(A => \I2.RAMDT4l0r_net_1\, B => 
        \I2.RAMDT4l6r_net_1\, Y => \I2.un21_pipe5_dt_0_net_1\);
    
    \I1.REG_74_0_IVL291R_1928\ : NOR2FT
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l291r_adt_net_121775_\);
    
    \I3.VDBil16r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_356_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil16r_net_1\);
    
    \I2.PIPE10_DT_625\ : MUX2L
      port map(A => \I2.PIPE10_DTl20r_net_1\, B => \I2.N_3806\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_625_net_1\);
    
    \I5.REG_1l429r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_42_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl429r);
    
    \I2.L2TYPEl0r_1542\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_589_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL0R_649\);
    
    \I1.REG_1_303\ : MUX2H
      port map(A => \REGl402r\, B => \I1.REG_74l402r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\, Y => 
        \I1.REG_1_303_net_1\);
    
    \I3.REGMAP_i_0_il45r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un206_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il45r_net_1\);
    
    \I1.REG_74_13_388_M8_I_1783\ : OAI21FTT
      port map(A => \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, 
        B => \I1.REG_74_13_388_N_16_adt_net_109531_\, C => 
        \I1.REG_74_12_300_N_15\, Y => 
        \I1.REG_74_13_388_N_11_adt_net_109571_\);
    
    \I2.un1_STATE1_38_0\ : AO21FTT
      port map(A => \I2.N_3292\, B => 
        \I2.un1_STATE1_38_adt_net_52564_\, C => 
        \I2.un1_STATE1_38_adt_net_52557_\, Y => 
        \I2.un1_STATE1_38\);
    
    \I5.SBYTE_68\ : MUX2H
      port map(A => \I5.SBYTEl3r_net_1\, B => \I5.N_20\, S => 
        \I5.N_406\, Y => \I5.SBYTE_68_net_1\);
    
    \I2.RAMAD_4_0l13r\ : MUX2H
      port map(A => \I2.RAMAD1l13r_net_1\, B => RAMAD_VMEl13r, S
         => \REG_i_il5r_adt_net_855552__net_1\, Y => \I2.N_540\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I179_Y\ : OR3
      port map(A => \I2.N302_0\, B => \I2.N481_adt_net_424217_\, 
        C => \I2.N481_adt_net_424221_\, Y => 
        \I2.N481_adt_net_88982_\);
    
    \I2.RAMDT4L12R_3071\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_825\);
    
    \I2.MIC_ERR_REGS_375\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl47r_net_1\, B => 
        \I2.MIC_ERR_REGSl46r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_375_net_1\);
    
    VAD_padl15r : IOB33PH
      port map(PAD => VAD(15), A => \I3.VADml15r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl15r);
    
    \I1.REG_9_sqmuxa_0_a2_0_0_a2\ : NAND3FFT
      port map(A => \I1.PAGECNTL7R_525\, B => \I1.N_1169\, C => 
        \I1.PAGECNTL8R_457\, Y => \I1.N_240\);
    
    \I3.VDBi_57l7r_adt_net_3750_\ : AO21
      port map(A => REGl7r, B => 
        \I3.VDBi_57l7r_adt_net_142960__net_1\, C => 
        \I3.VDBi_57l7r_adt_net_142961__net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_3750__net_1\);
    
    \I1.SBYTE_8_0_il3r\ : OA21
      port map(A => \I1.N_602_i\, B => REGl86r, C => 
        \I1.N_202_adt_net_105770_\, Y => \I1.N_202\);
    
    \I3.REG_1l109r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_290_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl109r);
    
    \I2.PIPE4_DTl11r_1147\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL11R_409\);
    
    \I2.UN1_REG80_I_1703\ : NOR3FTT
      port map(A => \I2.N_3824_adt_net_90289_\, B => REGl41r, C
         => REGl40r, Y => \I2.N_3824_adt_net_90295_\);
    
    REGl181r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_82_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl181r\);
    
    \I2.DTO_16_1_IV_0L27R_1079\ : AND2
      port map(A => \I2.DTO_1l27r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l27r_adt_net_29242_\);
    
    \I3.REGMAPl11r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un47_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl11r_net_1\);
    
    \I3.PIPEAl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_233_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl2r_net_1\);
    
    \I1.un1_sbyte13_1_i_0_s_830\ : AO21
      port map(A => \I1.N_370_adt_net_854904__net_1\, B => 
        \I1.un1_sbyte13_1_i_1_adt_net_106369__adt_net_854528__net_1\, 
        C => \PULSE_0L0R_ADT_NET_834380_RD1__199\, Y => 
        \I1.UN1_SBYTE13_1_I_1_208\);
    
    \I4.un4_bcnt_I_8\ : AND2
      port map(A => \I4.bcntl1r_net_1\, B => \I4.bcntl0r_net_1\, 
        Y => \I4.N_7\);
    
    \I2.un7_bnc_id_1_I_51\ : AND2
      port map(A => \I2.BNC_IDl8r_net_1\, B => 
        \I2.DWACT_FINC_El4r\, Y => \I2.N_14\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I167_Y\ : AO21TTF
      port map(A => \I2.N516\, B => \I2.N504_adt_net_88887_\, C
         => \I2.N357_1\, Y => \I2.N504\);
    
    \I1.REG_74_0_IV_0_O2L253R_1827\ : AOI21TTF
      port map(A => \I1.N_238_Rd1__adt_net_854884__net_1\, B => 
        \I1.REG_74_5_404_m1_e_0_net_1\, C => 
        \I1.REG_74_12_300_N_15\, Y => \I1.N_395_adt_net_113231_\);
    
    \I3.VDBOFFA_31_IV_0L7R_2509\ : OR3
      port map(A => \I3.VDBoffa_31l7r_adt_net_163317_\, B => 
        \I3.VDBoffa_31l7r_adt_net_163313_\, C => 
        \I3.VDBoffa_31l7r_adt_net_163314_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163320_\);
    
    \I3.UN1_STATE2_9_2310\ : NOR2
      port map(A => \I3.STATE2l0r_net_1\, B => 
        \I3.STATE2l1r_net_1\, Y => 
        \I3.un1_STATE2_9_adt_net_154004_\);
    
    \I3.VDBm_0l23r\ : MUX2L
      port map(A => \I3.PIPEAl23r_net_1\, B => 
        \I3.PIPEBl23r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_165\);
    
    \I2.N_199_0_ADT_NET_1054__2761\ : OAI21FTT
      port map(A => \I2.STATE2L3R_440\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.DTE_CL_0_SQMUXA_2_0_287\, Y => 
        \I2.N_199_0_ADT_NET_1054__37\);
    
    \I3.un1_NOEDTKi_0_sqmuxa_adt_net_135826_\ : AND2
      port map(A => \I3.ASBS_net_1\, B => \I3.STATE1_ipl5r\, Y
         => \I3.un1_NOEDTKi_0_sqmuxa_adt_net_135826__net_1\);
    
    \I1.REG_1_103\ : MUX2H
      port map(A => \REGl202r\, B => \I1.N_1341\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\, Y => 
        \I1.REG_1_103_net_1\);
    
    \I3.NRDMEBi_2_sqmuxa_2_1_a3\ : NOR2
      port map(A => \I3.N_1622_1\, B => 
        \I3.STATE2_ns_i_i_a5_0_a3l1r_adt_net_135757_\, Y => 
        \I3.N_12180_i\);
    
    \I2.PIPE8_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_547_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl19r_net_1\);
    
    \I2.DTE_21_1_iv_2l1r\ : AO21
      port map(A => \I2.STATE2L3R_440\, B => 
        \I2.DTO_9_ivl1r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39593_\, Y => 
        \I2.DTE_21_1_iv_2_il1r\);
    
    \I3.UN21_REG_ADS_0_A2_0_A3_1_2651\ : OR3
      port map(A => \I3.VASl12r_net_1\, B => \I3.VASl4r_net_1\, C
         => \I3.VASl2r_net_1\, Y => 
        \I3.un60_reg_ads_3_adt_net_166295_\);
    
    REGl195r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_96_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl195r\);
    
    \I2.RAMADl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l7r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl7r);
    
    \I1.REG_3_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_254_196\, B => \I1.N_242\, Y => 
        \I1.REG_3_sqmuxa\);
    
    \I3.RAMAD_VMEl6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_30_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl6r);
    
    \I2.TRGARR_3_I_21\ : AND2
      port map(A => \I2.DWACT_ADD_CI_0_g_array_1l0r\, B => 
        \I2.TRGARRl2r_net_1\, Y => 
        \I2.DWACT_ADD_CI_0_g_array_12l0r\);
    
    \I2.N_1170_adt_net_1217__adt_net_855700_\ : BFR
      port map(A => \I2.N_1170_adt_net_1217__net_1\, Y => 
        \I2.N_1170_adt_net_1217__adt_net_855700__net_1\);
    
    \I3.STATE1l7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl3r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl7r\);
    
    \I3.un2_reg_ads_0_a2_0_a3\ : NOR3FTT
      port map(A => \I3.WRITES_8\, B => \I3.N_581\, C => 
        \I3.un41_reg_ads_2\, Y => 
        \I3.un2_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.PIPE5_DT_6l2r\ : MUX2L
      port map(A => \I2.PIPE4_DTl2r_net_1\, B => \I2.N_1071\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, Y
         => \I2.PIPE5_DT_6l2r_net_1\);
    
    \I2.DTO_16_1_IV_0_0L19R_1123\ : AND2
      port map(A => \I2.DTO_1l19r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l19r_adt_net_30970_\);
    
    \I3.VDBi_40_1l3r\ : AND2FT
      port map(A => \I3.REGMAPl16r_net_1\, B => 
        \I3.VDBi_31l3r_net_1\, Y => \I3.N_341\);
    
    \I2.BNCID_VECT_tile_I_7\ : AND3FFT
      port map(A => \I2.I_6_2_i_0_i\, B => \I2.I_6_1_i_0_i\, C
         => \I2.N_13_adt_net_47925_\, Y => \I2.N_13\);
    
    \I1.REG_1_292\ : MUX2H
      port map(A => \REGl391r\, B => \I1.REG_74l391r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y => 
        \I1.REG_1_292_net_1\);
    
    \I1.REG_74_1_404_m7_i_a5_0\ : OR2FT
      port map(A => \I1.REG_74_2_0l404r_Rd1__net_1\, B => 
        \I1.REG_74_1_a0_0l228r_adt_net_854832__net_1\, Y => 
        \I1.REG_74_1_396_N_12\);
    
    \I2.DTE_1_851\ : MUX2L
      port map(A => \I2.DTE_1l11r_Rd1__net_1\, B => 
        \I2.DTE_21_1l11r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, Y => 
        \I2.DTE_1l11r\);
    
    \I1.REG_74_0_ivl297r\ : AO21
      port map(A => \REGl297r\, B => \I1.N_169\, C => 
        \I1.REG_74l297r_adt_net_121126_\, Y => \I1.REG_74l297r\);
    
    NMRSFIF_pad : OB33PH
      port map(PAD => NMRSFIF, A => NMRSFIF_c_c);
    
    \I1.REG_74_4_i_a2_404_N_4_i_adt_net_1465_\ : AND2
      port map(A => \I1.N_268_Rd1__net_1\, B => \I1.N_254_194\, Y
         => \I1.REG_74_4_i_a2_404_N_4_i_adt_net_1465__net_1\);
    
    \I3.REGMAPl17r_adt_net_854292_\ : BFR
      port map(A => \I3.REGMAPl17r_adt_net_854300__net_1\, Y => 
        \I3.REGMAPl17r_adt_net_854292__net_1\);
    
    \I3.EVREAD_DS_1_sqmuxa_i_s\ : AND2
      port map(A => \I3.N_1465\, B => \I3.un15_anycyc_net_1\, Y
         => \I3.N_1861\);
    
    \I2.PIPE1_DT_12l4r\ : MUX2L
      port map(A => \I2.TDCDASl4r_net_1\, B => 
        \I2.TDCDASl2r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855104__net_1\, Y
         => \I2.PIPE1_DT_12l4r_net_1\);
    
    \I2.TOKENB_TIMOUT_2_0_a3\ : AND3
      port map(A => \I2.N_177\, B => \I2.TOKENB_CNTl1r_net_1\, C
         => \I2.TOKENB_CNTl0r_net_1\, Y => \I2.TOKENB_TIMOUT_2\);
    
    \I3.VDBi_55l10r\ : MUX2H
      port map(A => \I3.VDBil10r_net_1\, B => 
        \I3.RAMDTSl10r_net_1\, S => 
        \I3.N_57_i_0_0_adt_net_854696__net_1\, Y => 
        \I3.VDBi_55l10r_net_1\);
    
    \I1.REG_1_294\ : MUX2H
      port map(A => \REGl393r\, B => \I1.REG_74l393r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y => 
        \I1.REG_1_294_net_1\);
    
    \I3.REG_44_i_o2_0l83r\ : NAND2
      port map(A => \I3.STATE1_ipl8r\, B => \I3.REGMAPl13r_net_1\, 
        Y => \I3.N_98_0\);
    
    \I1.un1_sbyte13_1_i_0_s_832\ : AO21
      port map(A => \I1.N_370_adt_net_854904__net_1\, B => 
        \I1.un1_sbyte13_1_i_1_adt_net_106369__adt_net_854528__net_1\, 
        C => \PULSE_0L0R_ADT_NET_834380_RD1__199\, Y => 
        \I1.UN1_SBYTE13_1_I_1_210\);
    
    \I2.WOFFSET_836\ : MUX2L
      port map(A => \I2.WOFFSETl9r_Rd1__net_1\, B => 
        \I2.N_4252_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835304_Rd1__net_1\, Y
         => \I2.WOFFSETl9r\);
    
    \I3.RAMAD_VMEl13r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_37_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl13r);
    
    \I2.TDCDBSl22r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl22r, Q => 
        \I2.TDCDBSl22r_net_1\);
    
    \I2.DTO_9_IVL14R_1146\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl14r_net_1\, C => 
        \I2.DTO_9l14r_adt_net_32134_\, Y => 
        \I2.DTO_9l14r_adt_net_32142_\);
    
    \I3.un37_reg_ads_0_a2_1_a2_0\ : OR2
      port map(A => \I3.N_547\, B => \I3.N_553\, Y => \I3.N_637\);
    
    \I2.BNCID_VECT_tile_0_DOUTl1r\ : MUX2L
      port map(A => \I2.DIN_REG1l1r\, B => \I2.DOUT_TMPl1r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl9r\);
    
    \I1.REG_1_106\ : MUX2H
      port map(A => \REGl205r\, B => \I1.N_280\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_106_net_1\);
    
    \I2.LSRAM_IN_407\ : MUX2L
      port map(A => \I2.PIPE5_DTl23r_net_1\, B => 
        \I2.LSRAM_INl23r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_407_net_1\);
    
    \I2.REG_1l34r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl34r);
    
    REGl167r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_68_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl167r\);
    
    \I2.TDCGDB1_1473\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => TDCGDB_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.TDCGDB1_580\);
    
    \I1.REG_74_1_380_m8_i_x3\ : XOR2
      port map(A => \I1.PAGECNTl9r_net_1\, B => 
        \I1.REG_74_1_380_N_14\, Y => \I1.REG_74_1_380_N_15_i_i_i\);
    
    \I1.REG_74_0_IVL381R_1812\ : AND2
      port map(A => \FBOUTl0r\, B => \I1.REG_28_sqmuxa\, Y => 
        \I1.REG_74l381r_adt_net_111921_\);
    
    \I3.STATE1_ns_0_iv_0_0_a3_0_1_0l7r\ : NOR3FTT
      port map(A => \I3.N_58_i_0_adt_net_134395_\, B => 
        \I3.REGMAPL25R_776\, C => \I3.REGMAPL22R_775\, Y => 
        \I3.N_58_i_0\);
    
    \I2.RAMAD1_12l12r\ : MUX2L
      port map(A => \I2.TDCDASl23r_net_1\, B => 
        \I2.TDCDBSl23r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855176__net_1\, Y => 
        \I2.RAMAD1_12l12r_net_1\);
    
    \I3.VDBi_57l7r_adt_net_143034_\ : AO21
      port map(A => \I3.N_2037\, B => \I3.N_2270\, C => 
        \I3.VDBi_57l7r_adt_net_143017__net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_143034__net_1\);
    
    \I3.un1_NRDMEBi_2_sqmuxa_3\ : AOI21TTF
      port map(A => \I3.STATE2l1r_net_1\, B => \I3.N_297\, C => 
        \I3.un1_NRDMEBi_2_sqmuxa_3_adt_net_153598_\, Y => 
        \I3.un1_NRDMEBi_2_sqmuxa_3_net_1\);
    
    \I2.FID_7_0_IVL25R_985\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl25r_net_1\, 
        Y => \I2.FID_7l25r_adt_net_19021_\);
    
    \I1.BYTECNTL3R_2917\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_311_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTL3R_434\);
    
    \I2.PIPE9_DT_276\ : MUX2L
      port map(A => \I2.PIPE9_DTl7r_net_1\, B => 
        \I2.PIPE8_DTl7r_net_1\, S => \I2.NWPIPE8_i_0_i_0_0\, Y
         => \I2.PIPE9_DT_276_net_1\);
    
    \I3.VDBoff_119\ : MUX2L
      port map(A => \I3.VDBoffl3r_net_1\, B => \I3.N_2067\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_119_net_1\);
    
    \I3.PIPEA1_12l13r\ : AND2
      port map(A => DPR_cl13r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854504__net_1\, Y => 
        \I3.PIPEA1_12l13r_net_1\);
    
    \I3.STATE2_NS_0L0R_2118\ : AOI21TTF
      port map(A => \I3.N_203_adt_net_854976__net_1\, B => 
        \I3.STATE2_ns_i_i_a5_0_a3l1r_adt_net_135757_\, C => 
        \I3.STATE2l4r_net_1\, Y => 
        \I3.STATE2_nsl0r_adt_net_136048_\);
    
    \I2.CRC32_12_0_0_x2l29r\ : XOR2FT
      port map(A => \I2.CRC32l29r_net_1\, B => \I2.N_4157_i_i\, Y
         => \I2.N_18_i_0_i_0\);
    
    \I1.REG_74L220R_2009\ : AND2FT
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__831\, B => 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__net_1\, Y => 
        \I1.N_89_adt_net_128729_\);
    
    SP3_pad : OB33PH
      port map(PAD => SP3, A => \GND\);
    
    \I2.PIPE6_DT_485\ : MUX2H
      port map(A => \I2.PIPE5_DTl31r_net_1\, B => 
        \I2.PIPE6_DTl31r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_485_net_1\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855532_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__281\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\);
    
    \I2.PIPE1_DT_42_1_ivl1r\ : OR3
      port map(A => \I2.PIPE1_DT_42l1r_adt_net_52046_\, B => 
        \I2.PIPE1_DT_42l1r_adt_net_52044_\, C => 
        \I2.PIPE1_DT_42l1r_adt_net_52045_\, Y => 
        \I2.PIPE1_DT_42l1r\);
    
    \I2.OFFSET_37_22l5r\ : MUX2L
      port map(A => \REGl242r\, B => \REGl178r\, S => 
        \I2.PIPE7_DTL27R_79\, Y => \I2.N_808\);
    
    REGl342r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_243_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl342r\);
    
    \I2.PIPE5_DT_676\ : MUX2L
      port map(A => \I2.PIPE5_DTl0r_net_1\, B => 
        \I2.PIPE5_DT_6l0r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_676_net_1\);
    
    \I2.OFFSET_37_6l5r\ : MUX2L
      port map(A => \I2.N_672\, B => \I2.N_664\, S => 
        \I2.PIPE7_DTL26R_352\, Y => \I2.N_680\);
    
    \I3.un51_reg_ads_0_a2_0_a3_0\ : NAND3
      port map(A => \I3.VASl4r_net_1\, B => \I3.VASl2r_net_1\, C
         => \I3.N_552\, Y => \I3.un41_reg_ads_0_a2_3_a3_0\);
    
    \I3.PIPEB_99\ : AO21
      port map(A => DPR_cl20r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\, 
        C => \I3.PIPEB_99_adt_net_159873_\, Y => 
        \I3.PIPEB_99_net_1\);
    
    \I3.STATE1_NS_1_IV_0L5R_2122\ : OA21
      port map(A => \I3.N_1920\, B => \I3.STATE1_ipl6r\, C => 
        \I3.DSS_9\, Y => \I3.STATE1_nsl5r_adt_net_136318_\);
    
    \I1.REG_74_0_ivl196r\ : AO21
      port map(A => \REGl196r\, B => \I1.N_65_92\, C => 
        \I1.REG_74l196r_adt_net_130925_\, Y => 
        \I1.REG_74l196r_net_1\);
    
    \I3.STATE1l1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_tr24_i_0_net_1\, CLR
         => \I3.N_1311_0\, Q => \I3.STATE1_ipl1r\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2520\ : AO21
      port map(A => \REGl211r\, B => 
        \I3.REGMAPl23r_adt_net_855012__net_1\, C => 
        \I3.N_2070_adt_net_163466_\, Y => 
        \I3.N_2070_adt_net_163501_\);
    
    \I2.LSRAM_INl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_414_0_0_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl31r_net_1\);
    
    \I2.PIPE1_DT_12l11r\ : MUX2L
      port map(A => \I2.TDCDASl11r_net_1\, B => 
        \I2.TDCDASl9r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, Y
         => \I2.PIPE1_DT_12l11r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2423\ : AND2
      port map(A => \REGl288r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162516_\);
    
    \I3.REG_1l137r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_185_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl137r\);
    
    \I2.un1_tdc_res_28_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl413r, Y => 
        \I2.N_4609_i_0\);
    
    \I1.REG_2_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_242\, B => \I1.N_259\, Y => 
        \I1.REG_2_sqmuxa\);
    
    \I1.PAGECNT_n8_i_i\ : OAI21
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_854520__net_1\, 
        B => \I1.N_409_i_i_0_i\, C => \I1.N_473_206\, Y => 
        \I1.N_1379\);
    
    \I3.STATE2l0r_1613\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE2_nsl4r\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.STATE2L0R_720\);
    
    \I5.COMMAND_50\ : MUX2H
      port map(A => \I5.COMMANDl13r_net_1\, B => 
        \I5.COMMAND_4l13r_net_1\, S => \I5.sstate1l13r_net_1\, Y
         => \I5.COMMAND_50_net_1\);
    
    \I5.AIR_WDATA_9l10r\ : AND2
      port map(A => \I5.SENS_ADDRl1r_net_1\, B => 
        \I5.sstate2l3r_net_1\, Y => \I5.AIR_WDATA_9l10r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L7R_2501\ : AO21
      port map(A => \REGl228r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.VDBoffa_31l7r_adt_net_163272_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163310_\);
    
    \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r\ : AO21FTT
      port map(A => \I3.N_2031\, B => \I3.N_1923\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_adt_net_146111_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_net_1\);
    
    \I2.RAMDT4L5R_2809\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_137\);
    
    \I1.REG_74_0_IVL230R_1996\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_9_sqmuxa_adt_net_854728__net_1\, Y => 
        \I1.REG_74l230r_adt_net_127624_\);
    
    \I2.PIPE4_DTl13r_1534\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl13r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL13R_641\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I187_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl17r_net_1\, Y => 
        \I2.ADD_21x21_fast_I187_Y_0\);
    
    \I2.FID_7_0_ivl30r\ : AO21
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl30r_net_1\, 
        C => \I2.FID_7l30r_adt_net_18559_\, Y => \I2.FID_7l30r\);
    
    \I2.DTO_9_IVL24R_1091\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => \I2.N_4194\, C
         => \I2.DTO_9l24r_adt_net_29794_\, Y => 
        \I2.DTO_9l24r_adt_net_29802_\);
    
    \I3.REG_1_219\ : MUX2L
      port map(A => VDB_inl6r, B => REGl412r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_219_0\);
    
    \I1.REG_1_155\ : MUX2H
      port map(A => \REGl254r\, B => \I1.REG_74l254r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_155_net_1\);
    
    \I1.REG_74_i_o2_0_0_m9_i_0_0\ : MUX2L
      port map(A => \I1.PAGECNTl5r_net_1\, B => 
        \I1.REG_74_1_396_m7_i_a5_0\, S => 
        \I1.REG_74_i_o2_0_0_364_N_14\, Y => 
        \I1.REG_74_i_o2_0_0_m9_i_0_0_net_1\);
    
    \I2.DTE_21_1_iv_2l3r\ : AO21
      port map(A => \I2.STATE2L3R_440\, B => 
        \I2.DTO_9_ivl3r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39313_\, Y => 
        \I2.DTE_21_1_iv_2_il3r\);
    
    \I1.N_50_0_ADT_NET_1409__2747\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__541\, B => 
        \I1.N_50_0_ADT_NET_109751__256\, Y => 
        \I1.N_50_0_ADT_NET_1409__20\);
    
    DTE_padl9r : IOB33PH
      port map(PAD => DTE(9), A => \I2.DTE_1l9r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl9r);
    
    \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836_\ : BFR
      port map(A => \I2.un1_STATE3_10_1_adt_net_999__net_1\, Y
         => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\);
    
    \I2.DTESl2r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl2r, Q => 
        \I2.DTESl2r_net_1\);
    
    \I1.REG_1_157\ : MUX2H
      port map(A => \REGl256r\, B => \I1.REG_74l256r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_157_net_1\);
    
    REGl357r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_258_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl357r\);
    
    \I3.DSSF1_2_I_I_O3_I_A3_2348\ : AND2
      port map(A => DS0B_c, B => DS1B_c, Y => 
        \I3.N_306_adt_net_161608_\);
    
    \I2.PIPE1_DT_30l10r\ : MUX2L
      port map(A => \I2.TDCDBSl10r_net_1\, B => 
        \I2.TDCDBSl8r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, Y
         => \I2.PIPE1_DT_30l10r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I121_Y_I_O2_1584\ : NOR2FT
      port map(A => \I2.N_64_0_adt_net_855028__net_1\, B => 
        \I2.N_28_0\, Y => \I2.N_29_i_0_adt_net_59529_\);
    
    \I2.PIPE1_DT_30l19r\ : MUX2L
      port map(A => \I2.TDCDBSl19r_net_1\, B => 
        \I2.TDCDBSl17r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, Y
         => \I2.PIPE1_DT_30l19r_net_1\);
    
    \I2.PIPE7_DTl25r_1578\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL25R_685\);
    
    \I3.un6_cycs_i_a3_0_a3\ : NOR2
      port map(A => \I3.CYCS_net_1\, B => \I3.ASBS_net_1\, Y => 
        \I3.N_1512\);
    
    \I2.REG_1_n14_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => REGl46r, Y => \I2.REG_1_n14_0_net_1\);
    
    \I2.REG_1_n3\ : XOR2
      port map(A => \I2.N_3831\, B => \I2.REG_1_n3_0_net_1\, Y
         => \I2.REG_1_n3_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I145_Y\ : AO21
      port map(A => \I2.N400_adt_net_88380_\, B => 
        \I2.N411_adt_net_4092__net_1\, C => \I2.N363\, Y => 
        \I2.N513\);
    
    \I2.BNCID_VECT_tile_0_DIN_REG1l3r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl11r_net_1\, Q => 
        \I2.DIN_REG1l3r\);
    
    \I3.un3_noe32wi_0_a2_i_o2\ : OR2
      port map(A => \I3.MBLTCYC_423\, B => 
        \I3.N_264_0_ADT_NET_1653_RD1__147\, Y => \I3.N_268\);
    
    \I3.VDBOFFA_31_IV_0L3R_2567\ : AND2
      port map(A => \REGl216r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.VDBoffa_31l3r_adt_net_164036_\);
    
    \I3.VDBI_57_IV_0_0L0R_2286\ : OA21TTF
      port map(A => \I3.VDBi_57l0r_adt_net_146601_\, B => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r\, C => 
        \I3.N_1905_1_adt_net_855384__net_1\, Y => 
        \I3.VDBi_57l0r_adt_net_146655_\);
    
    \I2.ROFFSET_906\ : MUX2H
      port map(A => \I2.ROFFSETl12r_net_1\, B => 
        \I2.ROFFSET_n12_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_906_net_1\);
    
    \I2.DT_SRAM_0_il17r\ : MUX2H
      port map(A => \I2.PIPE5_DTl17r_net_1\, B => 
        \I2.PIPE10_DTl17r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854216__net_1\, Y => 
        \I2.N_4645\);
    
    \I2.DTE_21_1l7r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l7r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l7r_Rd1__net_1\);
    
    \I5.DATAl9r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l9r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl126r);
    
    \I2.STATE1_ns_i_o3_i_a3l14r\ : AND2FT
      port map(A => \I2.N_3272_345\, B => \I2.STATE1l5r_net_1\, Y
         => \I2.N_158\);
    
    \I2.ADO_3l3r\ : MUX2L
      port map(A => \I2.WOFFSETl4r_adt_net_854980__net_1\, B => 
        \I2.ROFFSETl4r_net_1\, S => NOESRAME_C_243, Y => 
        \I2.ADO_3l3r_net_1\);
    
    \I3.REGMAPl2r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un13_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl2r_net_1\);
    
    \I2.WOFFSET_13_il6r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_31\, Y => \I2.N_4249\);
    
    \I2.FID_7_0_IVL25R_986\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl73r, C => 
        \I2.FID_7l25r_adt_net_19021_\, Y => 
        \I2.FID_7l25r_adt_net_19029_\);
    
    \I3.VDBOFFA_31_IV_0L3R_2569\ : AND2
      port map(A => \REGl272r\, B => \I3.REGMAPl31r_net_1\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164044_\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854580_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854580__net_1\);
    
    \I1.REG_1_245\ : MUX2H
      port map(A => \REGl344r\, B => \I1.REG_74l344r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_245_net_1\);
    
    \I5.COMMANDl11r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_48_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl11r_net_1\);
    
    \I1.REG_1_78\ : MUX2H
      port map(A => \REGl177r\, B => \I1.REG_74l177r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\, Y => 
        \I1.REG_1_78_net_1\);
    
    \I2.NPRSFIF\ : DFFC
      port map(CLK => CLK_c, D => \I2.NPRSFIF_328_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => NMRSFIF_c_c);
    
    ADE_padl2r : OB33PH
      port map(PAD => ADE(2), A => ADE_cl2r);
    
    \I3.VDBI_57_IV_0_0L0R_2285\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854356__net_1\, B
         => \I3.VDBoffl0r_net_1\, Y => 
        \I3.VDBi_57l0r_adt_net_146651_\);
    
    \I2.MIC_ERR_REGSl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_330_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl1r_net_1\);
    
    VDB_padl14r : IOB33PH
      port map(PAD => VDB(14), A => \I3.VDBml14r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl14r);
    
    \I2.N_152_i_0_adt_net_4117_\ : OR2
      port map(A => \I2.N_112_1\, B => 
        \I2.N_152_i_0_adt_net_55693__net_1\, Y => 
        \I2.N_152_i_0_adt_net_4117__net_1\);
    
    \I2.DTE_21_1_IV_2L3R_1336\ : OAI21TTF
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855208__net_1\, 
        B => \I2.DT_TEMPl3r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39303_\, Y => 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39312_\);
    
    \I1.REG_9_sqmuxa_adt_net_854724_\ : BFR
      port map(A => \I1.REG_9_sqmuxa\, Y => 
        \I1.REG_9_sqmuxa_adt_net_854724__net_1\);
    
    \I2.BNCID_VECT_tile_I_6_3\ : XOR2
      port map(A => \I2.WADDR_REG1l3r\, B => 
        \I2.TRGSERVl3r_net_1\, Y => \I2.I_6_3_i_0_i\);
    
    \I2.DT_SRAMl25r\ : MUX2L
      port map(A => \I2.N_893\, B => \I2.PIPE2_DTl25r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl25r_net_1\);
    
    \I2.DTE_1l4r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l4r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l4r_Rd1__net_1\);
    
    \I1.REG_15_sqmuxa_0_a2_897\ : OR2
      port map(A => \I1.REG_15_sqmuxa_adt_net_1457__net_1\, B => 
        \I1.N_254_277\, Y => \I1.REG_15_SQMUXA_275\);
    
    PWR_i : PWR
      port map(Y => \VCC\);
    
    \I2.resyn_0_I2_TRGCNT_c3_i\ : OAI21TTF
      port map(A => \I2.TRGCNT_i_0_il3r\, B => 
        \I2.un9_tdctrgi_i_0\, C => \I2.N_3764_adt_net_16233_\, Y
         => \I2.N_3764\);
    
    \I2.PIPE8_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_534_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl6r_net_1\);
    
    \I3.DSSF1_42\ : MUX2L
      port map(A => \I3.DSSF1_net_1\, B => \I3.N_306\, S => 
        \I3.N_1512\, Y => \I3.DSSF1_42_net_1\);
    
    \I2.DTE_21_1_iv_0_x2l13r\ : XOR2
      port map(A => \I2.CRC32l9r_net_1\, B => 
        \I2.CRC32l21r_net_1\, Y => \I2.N_44_i_0\);
    
    \I2.WOFFSETl0r_adt_net_854636__adt_net_855712_\ : BFR
      port map(A => \I2.WOFFSETl0r_adt_net_854636__net_1\, Y => 
        \I2.WOFFSETl0r_adt_net_854636__adt_net_855712__net_1\);
    
    \I3.PIPEA_8l6r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854480__net_1\, B => 
        \I3.N_215\, Y => \I3.PIPEA_8l6r_net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854576_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854576__net_1\);
    
    \I2.DTO_16_1_IV_0L27R_1080\ : AO21
      port map(A => \I2.G_EVNT_NUMl11r_net_1\, B => \I2.N_457\, C
         => \I2.DTO_16_1l27r_adt_net_29240_\, Y => 
        \I2.DTO_16_1l27r_adt_net_29251_\);
    
    \I2.PIPE1_DT_30l14r\ : MUX2L
      port map(A => \I2.TDCDBSl14r_net_1\, B => 
        \I2.TDCDBSl12r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, Y
         => \I2.PIPE1_DT_30l14r_net_1\);
    
    \I2.MIC_ERR_REGS_355\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl27r_net_1\, B => 
        \I2.MIC_ERR_REGSl26r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_355_net_1\);
    
    \I3.REG_1_181\ : MUX2L
      port map(A => VDB_inl0r, B => \I3.REGl133r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, Y => 
        \I3.REG_1_181_0\);
    
    \I2.un2_evnt_word_I_52\ : XOR2
      port map(A => \I2.N_19\, B => \I2.WOFFSETl9r\, Y => 
        \I2.I_52\);
    
    REGl362r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_263_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl362r\);
    
    \I2.BNCID_VECTror_9_tz\ : AND2
      port map(A => \I2.BNCID_VECTra12_1_net_1\, B => 
        \I2.BNCID_VECTro_12\, Y => 
        \I2.BNCID_VECTror_9_tz_adt_net_48087_\);
    
    \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1570_\ : NAND3FFT
      port map(A => \I3.REGMAPl34r_net_1\, B => 
        \I3.REGMAPl43r_net_1\, C => \I3.N_560_adt_net_134484_\, Y
         => \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1570__net_1\);
    
    \I2.TDCDASl16r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl16r, Q => 
        \I2.TDCDASl16r_net_1\);
    
    \I2.REG_1l34r_1456\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL34R_563);
    
    \I2.PIPE8_DT_531\ : MUX2L
      port map(A => \I2.PIPE8_DTl3r_net_1\, B => 
        \I2.PIPE8_DT_21l3r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_531_net_1\);
    
    \I2.DTO_16_1l26r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l26r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l26r_Rd1__net_1\);
    
    \I2.STATE2L3R_2920\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl2r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L3R_437\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855412_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__321\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\);
    
    \I3.un136_reg_ads_0_a2_2_a2_0_987\ : NAND2FT
      port map(A => \I3.VASl2r_net_1\, B => \I3.N_548_368\, Y => 
        \I3.N_549_365\);
    
    \I2.PIPE5_DT_6l14r\ : MUX2L
      port map(A => \I2.PIPE4_DTl14r_net_1\, B => \I2.N_1083\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\, Y
         => \I2.PIPE5_DT_6l14r_net_1\);
    
    \I2.N_118_i_1_adt_net_1122_\ : OR3
      port map(A => \I2.sram_empty_1_i_0_i\, B => 
        \I2.sram_empty_3_i_0_i\, C => 
        \I2.N_118_i_1_adt_net_24217__net_1\, Y => 
        \I2.N_118_i_1_adt_net_1122__net_1\);
    
    \I4.bcnt_3l3r\ : AND2
      port map(A => \I4.N_48_3\, B => \I4.I_13_0\, Y => 
        \I4.bcnt_3l3r_net_1\);
    
    \I3.VDBi_57_0_ivl26r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l26r_net_1\, C
         => \I3.VDBi_57l26r_adt_net_138577_\, Y => 
        \I3.VDBi_57l26r\);
    
    \I1.REG_1_153\ : MUX2H
      port map(A => \REGl252r\, B => \I1.REG_74l252r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_153_net_1\);
    
    \I2.PIPE9_DT_272\ : MUX2L
      port map(A => \I2.PIPE9_DTl3r_net_1\, B => 
        \I2.PIPE8_DTl3r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_272_net_1\);
    
    \I1.N_273_6_i_0_adt_net_854796_\ : BFR
      port map(A => \I1.N_273_6_i_0\, Y => 
        \I1.N_273_6_i_0_adt_net_854796__net_1\);
    
    \I2.STATE1l6r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3875_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1l6r_net_1\);
    
    \I2.RAMAD1_666\ : MUX2L
      port map(A => \I2.RAMAD1_12l12r_net_1\, B => 
        \I2.RAMAD1l12r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__171\, Y => 
        \I2.RAMAD1_666_net_1\);
    
    \I3.VDBOFFB_30_IV_0L7R_2361\ : AO21
      port map(A => \REGl340r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l7r_adt_net_161768_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161794_\);
    
    \I1.NWRLUT\ : DFFS
      port map(CLK => CLK_c, D => \I1.NWRLUTi_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => NWRLUT_c);
    
    REGl198r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_99_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl198r\);
    
    \I3.un1_STATE2_11_adt_net_153679_\ : NAND2FT
      port map(A => DPR_cl31r, B => DPR_cl30r, Y => 
        \I3.un1_STATE2_11_adt_net_153679__net_1\);
    
    \I3.PIPEA_8_0l24r\ : MUX2L
      port map(A => DPR_cl24r, B => \I3.PIPEA1l24r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855360__net_1\, Y => \I3.N_233\);
    
    \I2.DTO_9_IVL11R_1162\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        B => \I2.DTE_2_1l11r_net_1\, Y => 
        \I2.DTO_9l11r_adt_net_32804_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I201_Y\ : XOR2FT
      port map(A => \I2.N516\, B => \I2.SUB_21x21_fast_I201_Y_0\, 
        Y => \I2.SUB8_2l5r\);
    
    \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834772_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_0_sqmuxa_i_0_N_3_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834772_Rd1__net_1\);
    
    \I1.N_268_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_268_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_268_Rd1__net_1\);
    
    \I2.STATE4_ns_i_0_m2l1r\ : MUX2L
      port map(A => \I2.N_4464\, B => \I2.N_4462\, S => REGl1r, Y
         => \I2.N_4481\);
    
    \I2.LSRAM_RDi_486\ : MUX2H
      port map(A => \I2.N_4524\, B => \I2.LSRAM_RDi_net_1\, S => 
        END_FLUSH_560, Y => \I2.LSRAM_RDi_486_net_1\);
    
    \I2.DT_SRAM_0l3r\ : MUX2L
      port map(A => \I2.PIPE10_DTl3r_net_1\, B => 
        \I2.PIPE5_DTl3r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, Y => 
        \I2.N_871\);
    
    \I3.REG_1_i_il1r\ : AO21
      port map(A => \I3.REG3l1r_net_1\, B => \I3.REG2l1r_net_1\, 
        C => \REGl1r_adt_net_21137_\, Y => REGl1r);
    
    \I2.SUB9_1_ADD_18x18_fast_I112_Y\ : OA21
      port map(A => \I2.N336\, B => \I2.N329\, C => 
        \I2.N448_i_adt_net_71546_\, Y => \I2.N448_i\);
    
    DTO_padl8r : IOB33PH
      port map(PAD => DTO(8), A => \I2.DTO_1l8r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl8r);
    
    \I2.WROi_793\ : MUX2L
      port map(A => \I2.WROi_net_1\, B => \I2.WROi_10\, S => 
        \I2.un1_DTO_cl_0_sqmuxa\, Y => \I2.WROi_793_net_1\);
    
    \I3.VDBi_345\ : MUX2L
      port map(A => \I3.VDBil5r_net_1\, B => \I3.VDBi_57l5r\, S
         => \I3.un1_STATE1_13_1_adt_net_1351__net_1\, Y => 
        \I3.VDBi_345_net_1\);
    
    \I3.VDBI_57_IV_0_0L2R_2265\ : AO21
      port map(A => \I3.VDBil2r_net_1\, B => \I3.N_2048\, C => 
        \I3.VDBi_57l2r_adt_net_145368_\, Y => 
        \I3.VDBi_57l2r_adt_net_145381_\);
    
    \I1.REG_74_1_380_m8_i_o3\ : NAND3
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        B => \I1.PAGECNTl7r_net_1\, C => 
        \I1.PAGECNTl6r_adt_net_854924__net_1\, Y => 
        \I1.REG_74_1_380_N_14\);
    
    \I2.PIPE1_DT_42_1_IV_2L27R_1363\ : NOR2
      port map(A => \I2.TDCDASl27r_net_1\, B => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855036__net_1\, 
        Y => \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46027_\);
    
    \I1.REG_74_0_IV_0L215R_2019\ : AND2
      port map(A => \REGl215r\, B => \I1.N_89_164\, Y => 
        \I1.REG_74l215r_adt_net_129206_\);
    
    \I2.EVNT_WORDl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_720_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl7r_net_1\);
    
    \I2.L2TYPEl1r_1550\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_590_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_I_0_IL1R_657\);
    
    \I2.WPAGE_0_sqmuxa_0_a6_0_a2\ : AND2FT
      port map(A => NOESRAME_C_242, B => \I2.STATE2l1r\, Y => 
        \I2.WPAGEe\);
    
    \I3.un1_NOEDTKi_0_sqmuxa_1_0\ : OR3
      port map(A => \I3.N_1516\, B => 
        \I3.un1_NOEDTKi_0_sqmuxa_1_adt_net_159328_\, C => 
        \I3.un1_NOEDTKi_0_sqmuxa\, Y => 
        \I3.un1_NOEDTKi_0_sqmuxa_1\);
    
    \I2.PIPE6_DT_0_sqmuxa_i_m2_1\ : MUX2L
      port map(A => LEAD_FLAGl6r, B => LEAD_FLAGl4r, S => 
        \I2.PIPE5_DTL22R_666\, Y => \I2.N_4544\);
    
    \I2.PIPE1_DT_42_1_IVL5R_1494\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855224__net_1\, B => 
        \I2.MIC_ERR_REGSl5r_net_1\, C => 
        \I2.PIPE1_DT_42l5r_adt_net_51185_\, Y => 
        \I2.PIPE1_DT_42l5r_adt_net_51186_\);
    
    \I1.REG_74l348r\ : OR3FFT
      port map(A => \I1.REG_24_sqmuxa\, B => \I1.REG_74_0l348r\, 
        C => \I1.N_41_9_adt_net_854784__net_1\, Y => \I1.N_217\);
    
    \I2.DTESl18r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl18r, Q => 
        \I2.DTESl18r_net_1\);
    
    \I2.OFFSET_37_16l7r\ : MUX2L
      port map(A => \REGl268r\, B => \REGl204r\, S => 
        \I2.PIPE7_DTL27R_75\, Y => \I2.N_762\);
    
    \I2.DTO_1_883\ : MUX2L
      port map(A => \I2.DTO_1l9r_Rd1__net_1\, B => 
        \I2.DTO_16_1l9r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834772_Rd1__net_1\, Y
         => \I2.DTO_1l9r\);
    
    VDB_padl27r : IOB33PH
      port map(PAD => VDB(27), A => \I3.VDBml27r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl27r);
    
    \I2.STATEe_nsl0r\ : AO21
      port map(A => \I2.N_3510\, B => \I2.STATEel4r_net_1\, C => 
        \I2.STATEe_nsl0r_adt_net_23014_\, Y => 
        \I2.STATEe_nsl0r_net_1\);
    
    \I1.SSTATE_TR18_0_A2_0_A4_1763\ : AND2FT
      port map(A => \I1.COMMAND_716\, B => \I1.LUT_760\, Y => 
        \I1.sstate_ns_il5r_adt_net_107266_\);
    
    \I3.PIPEA1_306\ : MUX2L
      port map(A => \I3.PIPEA1l8r_net_1\, B => 
        \I3.PIPEA1_12l8r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__254\, Y => 
        \I3.PIPEA1_306_net_1\);
    
    \I1.REG_1_156\ : MUX2H
      port map(A => \REGl255r\, B => \I1.REG_74l255r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_156_net_1\);
    
    \I1.sstate_ns_0_iv_0_0_o2_0l2r\ : OR3FFT
      port map(A => \I1.BYTECNT_314_net_1\, B => 
        \I1.N_304_RA1__216\, C => \I1.BYTECNT_306_net_1\, Y => 
        \I1.N_317_Ra1_\);
    
    \I1.REG_1_114\ : MUX2H
      port map(A => \REGl213r\, B => \I1.REG_74l213r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_114_net_1\);
    
    \I3.REG_1_194\ : MUX2L
      port map(A => VDB_inl13r, B => \I3.REGl146r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, Y => 
        \I3.REG_1_194_0\);
    
    \I2.DT_TEMP_7l25r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854236__net_1\, B => 
        \I2.DT_SRAMl25r_net_1\, Y => \I2.DT_TEMP_7l25r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL1R_1519\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, B => 
        \I2.PIPE1_DT_30l1r_net_1\, C => 
        \I2.PIPE1_DT_42l1r_adt_net_52031_\, Y => 
        \I2.PIPE1_DT_42l1r_adt_net_52046_\);
    
    \I2.un28_sram_empty_10_0\ : MUX2L
      port map(A => \I2.N_628\, B => \I2.N_627\, S => 
        \I2.RPAGEL14R_613\, Y => \I2.N_629\);
    
    \I2.DTESl14r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl14r, Q => 
        \I2.DTESl14r_net_1\);
    
    \I3.REGMAP_i_0_a2_8l52r\ : NOR2
      port map(A => \I3.REGMAPL11R_743\, B => \I3.REGMAPL12R_746\, 
        Y => \I3.N_590\);
    
    \I3.REGMAP_I_0_A2L52R_2092\ : NOR3FTT
      port map(A => \I3.N_638_adt_net_134637_\, B => 
        \I3.REGMAPl6r_net_1\, C => \I3.REGMAPl50r_net_1\, Y => 
        \I3.N_638_adt_net_134643_\);
    
    \I2.un2_evnt_word_I_16\ : AND3
      port map(A => \I2.WOFFSETl0r_adt_net_854636__net_1\, B => 
        \I2.WOFFSETl1r_adt_net_854992__net_1\, C => 
        \I2.WOFFSETl2r_adt_net_854984__net_1\, Y => 
        \I2.DWACT_FINC_E_0l0r\);
    
    \I2.DTE_21_1_iv_0_o2_1_0l21r\ : OAI21FTT
      port map(A => \I2.STATE2L3R_440\, B => \I2.N_4283_I_0_234\, 
        C => \I2.DTO_cl_0_sqmuxa_0_adt_net_855200__net_1\, Y => 
        \I2.N_4038\);
    
    \I1.PAGECNT_325_1231\ : MUX2H
      port map(A => \I1.PAGECNTl2r_adt_net_834908_Rd1__net_1\, B
         => \I1.PAGECNT_n2\, S => 
        \I1.PAGECNTe_adt_net_854892__net_1\, Y => 
        \I1.PAGECNT_325_493\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I140_Y_0_o2_1\ : OR3FFT
      port map(A => \I2.N_107\, B => \I2.N_128_133\, C => 
        \I2.N_74_i_0_i_adt_net_54331_\, Y => \I2.N_74_i_0_i\);
    
    \I3.un166_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_580\, Y => 
        \I3.un166_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.PIPE10_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_615_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl10r_net_1\);
    
    \I2.PIPE8_DT_549\ : MUX2L
      port map(A => \I2.PIPE8_DTl21r_net_1\, B => 
        \I2.PIPE8_DT_21l21r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_549_net_1\);
    
    \I1.REG_74_0_IV_0L217R_2017\ : AND2
      port map(A => \FBOUTl4r\, B => \I1.REG_7_sqmuxa\, Y => 
        \I1.REG_74l217r_adt_net_129034_\);
    
    \I2.RAMADl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l17r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl17r);
    
    \I1.REG_74_0_IVL302R_1916\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l302r_adt_net_120696_\);
    
    \I2.PIPE1_DT_42_1_IVL28R_1361\ : NOR3FFT
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096__net_1\, B
         => \I2.TDCDASl28r_net_1\, C => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        Y => \I2.PIPE1_DT_42l28r_adt_net_45929_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I200_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl4r\, B => 
        \I2.PIPE7_DTl4r_net_1\, Y => \I2.SUB_21x21_fast_I200_Y_0\);
    
    \I5.sstate1l1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.N_95\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l1r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL13R_1445\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl45r_net_1\, C => 
        \I2.PIPE1_DT_42l13r_adt_net_49191_\, Y => 
        \I2.PIPE1_DT_42l13r_adt_net_49209_\);
    
    \I2.DTE_21_1_ivl15r\ : AO21
      port map(A => \I2.DTE_1l15r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.DTE_21_1l15r_adt_net_37953_\, Y => \I2.DTE_21_1l15r\);
    
    \I2.I_1335_s\ : XOR2
      port map(A => \I2.SUB8l3r_net_1\, B => \I2.OFFSETl0r_net_1\, 
        Y => \I2.SUB9_1l2r\);
    
    \I3.VDBI_20_IVL11R_2208\ : AND2
      port map(A => REGl59r, B => 
        \I3.REGMAPl9r_adt_net_854320__net_1\, Y => 
        \I3.VDBi_20l11r_adt_net_141166_\);
    
    \I2.EVNT_NUMl2r_1489\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_961_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUML2R_596\);
    
    \I1.REG_74_0_IVL398R_1791\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_30_sqmuxa_adt_net_854372__net_1\, Y => 
        \I1.REG_74l398r_adt_net_110272_\);
    
    \I2.un2_evnt_word_I_66\ : XOR2
      port map(A => \I2.WOFFSETl11r\, B => \I2.N_9_1\, Y => 
        \I2.I_66\);
    
    \I2.SUB9_1_ADD_18x18_fast_I70_Y\ : AO21
      port map(A => \I2.N307_1\, B => \I2.N304\, C => \I2.N303\, 
        Y => \I2.N338\);
    
    \I3.VDBi_20_ivl4r\ : NOR3
      port map(A => \I3.REGMAPL7R_460\, B => \I3.N_1907_264\, C
         => \I3.REGMAPl3r_net_1\, Y => 
        \I3.VDBi_20l4r_adt_net_414785_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I206_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl10r\, B => 
        \I2.PIPE7_DTl10r_net_1\, Y => 
        \I2.SUB_21x21_fast_I206_Y_0\);
    
    \I3.REG_1l54r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_155_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl54r);
    
    \I1.PAGECNT_320_adt_net_854876_\ : BFR
      port map(A => \I1.PAGECNT_320_net_1\, Y => 
        \I1.PAGECNT_320_adt_net_854876__net_1\);
    
    \I1.REG_1_232\ : MUX2H
      port map(A => \REGl331r\, B => \I1.REG_74l331r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y => 
        \I1.REG_1_232_net_1\);
    
    \I3.VDBI_57_IV_0_0L6R_2238\ : AO21
      port map(A => \I3.VDBil6r_net_1\, B => \I3.N_2048\, C => 
        \I3.VDBi_57l6r_adt_net_143390_\, Y => 
        \I3.VDBi_57l6r_adt_net_143403_\);
    
    \I2.LSRAM_INl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_400_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl16r_net_1\);
    
    \I2.PIPE9_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_273_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl4r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I2_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L9R_768\, B => \I2.PIPE4_DTL2R_513\, 
        Y => \I2.N_52_0\);
    
    \I2.WR_SRAM_2_ADT_NET_748__2762\ : OAI21FTF
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__889\, B => 
        \I2.N_4030\, C => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20049__net_1\, Y => 
        \I2.WR_SRAM_2_ADT_NET_748__39\);
    
    \I1.BYTECNT_306\ : MUX2H
      port map(A => \I1.BYTECNTl8r_net_1\, B => \I1.N_1162\, S
         => \I1.N_1383_225\, Y => \I1.BYTECNT_306_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I50_Y_1685\ : AND2FT
      port map(A => \I2.LSRAM_OUTl15r\, B => 
        \I2.PIPE7_DTl15r_net_1\, Y => \I2.N300_0_adt_net_87046_\);
    
    \I1.REG_1_80\ : MUX2H
      port map(A => \REGl179r\, B => \I1.REG_74l179r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\, Y => 
        \I1.REG_1_80_net_1\);
    
    \I2.CRC32l30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_825_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l30r_net_1\);
    
    \I2.DT_SRAM_i_m2l17r\ : MUX2L
      port map(A => \I2.N_4645\, B => \I2.PIPE2_DTl17r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.N_188\);
    
    LSRAM_FL_RADDRl1r : DFFC
      port map(CLK => CLK_c, D => \I4.LSRAM_FL_RADDR_10\, CLR => 
        CLEAR_STAT_i_0, Q => \LSRAM_FL_RADDRl1r\);
    
    \I3.REGMAPl55r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un224_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPl55r_net_1\);
    
    \I2.DTE_1l17r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l17r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l17r_Rd1__net_1\);
    
    \I1.REG_74_3l188r\ : OR2
      port map(A => \I1.N_1370_adt_net_112317_\, B => 
        \I1.N_41_9_ADT_NET_3739__93\, Y => \I1.N_97_2\);
    
    \I3.VDBI_20_IVL12R_2204\ : NOR2FT
      port map(A => \I3.N_2018\, B => \I3.N_1907\, Y => 
        \I3.VDBi_20l12r_adt_net_140770_\);
    
    \I2.N_565_0_adt_net_855732_\ : BFR
      port map(A => \I2.N_565_0\, Y => 
        \I2.N_565_0_adt_net_855732__net_1\);
    
    \I2.un28_sram_empty_9_0\ : MUX2L
      port map(A => \I2.L2TYPE_I_0_IL13R_660\, B => 
        \I2.L2TYPE_I_0_IL5R_659\, S => \I2.RPAGEL15R_519\, Y => 
        \I2.N_628\);
    
    \I1.BITCNT_n0_i_o3_0\ : AO21FTF
      port map(A => \I1.BITCNTl0r_net_1\, B => \I1.N_1376_i_0\, C
         => \I1.N_604\, Y => \I1.N_1199\);
    
    \I2.un1_tdc_res_36_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl416r, Y => 
        \I2.N_4617_i_0\);
    
    \I2.SUB9_1_ADD_18x18_fast_I115_Y\ : OR2
      port map(A => \I2.N457_adt_net_69532_\, B => \I2.N334\, Y
         => \I2.N457\);
    
    \I2.N477_adt_net_301898_\ : AND2
      port map(A => \I2.N299_0\, B => \I2.N346_0_542\, Y => 
        \I2.N477_adt_net_301898__net_1\);
    
    TDCDB_padl23r : IB33
      port map(PAD => TDCDB(23), Y => TDCDB_cl23r);
    
    \I1.REG_1_234\ : MUX2H
      port map(A => \REGl333r\, B => \I1.REG_74l333r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y => 
        \I1.REG_1_234_net_1\);
    
    \I1.REG_1_281\ : MUX2H
      port map(A => \REGl380r\, B => \I1.REG_74l380r_net_1\, S
         => \I1.N_50_0_ADT_NET_1409__282\, Y => 
        \I1.REG_1_281_net_1\);
    
    \I2.DT_TEMP_7l19r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854240__net_1\, B => 
        \I2.DT_SRAMl19r_net_1\, Y => \I2.DT_TEMP_7l19r_net_1\);
    
    \I2.FID_7_0_ivl29r\ : AO21
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl29r_net_1\, 
        C => \I2.FID_7l29r_adt_net_18653_\, Y => \I2.FID_7l29r\);
    
    \I2.STATE1_ns_a3_i_o3l12r\ : NAND2
      port map(A => \I2.STATE1L7R_632\, B => \I2.N_3883\, Y => 
        \I2.N_3889\);
    
    \I2.OFFSET_565\ : MUX2L
      port map(A => \I2.OFFSETl5r_net_1\, B => \I2.OFFSET_37l5r\, 
        S => \I2.UN1_NWPIPE7_2_297\, Y => \I2.OFFSET_565_net_1\);
    
    \I2.CRC32_12_il13r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_115_i_i_0\, Y => 
        \I2.N_3930\);
    
    \I2.WREi_8_i_i_a2_1\ : OR3
      port map(A => \I2.STATE2l5r_net_1\, B => 
        \I2.STATE2l2r_adt_net_855212__net_1\, C => 
        \I2.WPAGEe_adt_net_855060__net_1\, Y => 
        \I2.WREi_8_i_i_a2_1_net_1\);
    
    \I2.PIPE5_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_702_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl26r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I15_P0N_i_o3\ : OR2
      port map(A => \I2.RAMDT4L12R_798\, B => 
        \I2.PIPE4_DTl15r_net_1\, Y => \I2.N_32_0\);
    
    \I3.VDBOFFA_50_2528\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal6r_net_1\, Y => 
        \I3.VDBoffa_50_adt_net_163548_\);
    
    \I3.REG_1_218\ : MUX2L
      port map(A => VDB_inl5r, B => REGl411r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_218_0\);
    
    \I2.REG_1_n13_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => REGl45r, Y => \I2.REG_1_n13_0_net_1\);
    
    \I5.DATAl7r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12_ivl1r_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => REGl118r);
    
    \I3.REGMAPl14r_1628\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un57_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL14R_735\);
    
    REGl296r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_197_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl296r\);
    
    \I5.N_155_0_adt_net_983_\ : AO21FTT
      port map(A => \I5.COMMANDl0r_net_1\, B => 
        \I5.N_75_adt_net_8973_\, C => \I5.sstate1l11r_net_1\, Y
         => \I5.N_155_0_adt_net_983__net_1\);
    
    \I5.un1_SENS_ADDR_1_I_1\ : NOR2FT
      port map(A => \I5.SENS_ADDRl0r_net_1\, B => 
        \I5.REG_2_sqmuxa_0_adt_net_975__net_1\, Y => 
        \I5.DWACT_ADD_CI_0_TMPl0r\);
    
    \I3.REG_1_269\ : MUX2H
      port map(A => REGl88r, B => \I3.N_1634\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_269_0\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I62_Y_1677\ : AND2FT
      port map(A => \I2.LSRAM_OUTl9r\, B => \I2.PIPE7_DTL9R_696\, 
        Y => \I2.N312_0_adt_net_86445_\);
    
    \I1.N_317_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_317_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_317_Rd1__net_1\);
    
    VAD_padl7r : IOB33PH
      port map(PAD => VAD(7), A => \I3.VADml7r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl7r);
    
    \I2.PIPE5_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_704_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl28r_net_1\);
    
    \I3.VDBi_57_iv_0l5r\ : OR3
      port map(A => \I3.VDBi_57l5r_adt_net_143854_\, B => 
        \I3.VDBi_57l5r_adt_net_143862_\, C => 
        \I3.VDBi_57l5r_adt_net_143863_\, Y => \I3.VDBi_57l5r\);
    
    \I3.VDBOFFB_30_IV_0L3R_2426\ : AND2
      port map(A => \REGl304r\, B => \I3.REGMAPl35r_net_1\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162528_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I136_Y_0_o2_m4_4\ : AOI21
      port map(A => \I2.N_45_1_105\, B => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_N_6_i_adt_net_56545_\, C
         => \I2.ADD_21x21_fast_I136_Y_0_o2_m4_2_i_adt_net_56602_\, 
        Y => \I2.ADD_21x21_fast_I136_Y_0_o2_m4_4_adt_net_56769_\);
    
    \I1.REG_74_0_ivl340r\ : AO21
      port map(A => \REGl340r\, B => \I1.N_209\, C => 
        \I1.REG_74l340r_adt_net_117228_\, Y => 
        \I1.REG_74l340r_net_1\);
    
    \I3.PIPEBl10r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_89_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl10r_net_1\);
    
    \I2.REG_1_C3_I_1744\ : AND2
      port map(A => \I2.un8_evread_1_adt_net_855780__net_1\, B
         => \I2.N_122\, Y => \I2.N_3832_adt_net_101536_\);
    
    \I3.PULSE_330\ : AO21
      port map(A => \I3.N_311_adt_net_854752__net_1\, B => 
        \I3.N_116_adt_net_134828_\, C => 
        \I3.PULSE_330_adt_net_134909_\, Y => \I3.PULSE_330_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I174_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l4r_net_1\, B => 
        \I2.PIPE4_DTL4R_478\, Y => \I2.ADD_21x21_fast_I174_Y_0\);
    
    \I3.STATE1_408\ : OR2
      port map(A => \I3.STATE1_ipl7r\, B => 
        \I3.N_1174_adt_net_1495__net_1\, Y => \I3.N_1174\);
    
    \I2.G_EVNT_NUM_n2_i_0_a2\ : NOR2
      port map(A => \I2.N_186\, B => \I2.G_EVNT_NUMl2r_net_1\, Y
         => \I2.N_316_i\);
    
    \I1.REG_74_0_ivl382r\ : AO21
      port map(A => \REGl382r\, B => \I1.N_257\, C => 
        \I1.REG_74l382r_adt_net_111835_\, Y => \I1.REG_74l382r\);
    
    \I1.PAGECNT_n4_0_0_x2\ : XOR2FT
      port map(A => \I1.PAGECNTl4r_adt_net_835120_Rd1__net_1\, B
         => \I1.N_308_Rd1__net_1\, Y => \I1.N_394_i_i_0_i\);
    
    VDB_padl22r : IOB33PH
      port map(PAD => VDB(22), A => \I3.VDBml22r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl22r);
    
    \I3.VDBi_31l11r\ : MUX2L
      port map(A => \I3.REGl144r\, B => \I3.VDBi_20l11r\, S => 
        \I3.REGMAPl17r_adt_net_854288__net_1\, Y => 
        \I3.VDBi_31l11r_net_1\);
    
    \I2.N_4283_i_0_a2_m1_e_0_663\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854444__net_1\, 
        B => \I2.TEMPF_adt_net_855740__net_1\, Y => 
        \I2.N_4283_I_0_41\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I152_Y_0_2711\ : NAND3
      port map(A => \I2.N502_i_0_adt_net_490246_\, B => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_adt_net_56806_\, C => 
        \I2.N502_i_0_adt_net_490398_\, Y => 
        \I2.N498_0_adt_net_598321_\);
    
    \I2.STATE1l4r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_il14r_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.STATE1l4r_net_1\);
    
    \I3.VDBi_40l4r\ : MUX2L
      port map(A => \I3.N_342\, B => \I3.N_136\, S => 
        \I3.N_354_0_adt_net_855368__net_1\, Y => 
        \I3.VDBi_40l4r_net_1\);
    
    \I1.N_41_9_adt_net_3739_\ : NAND2
      port map(A => \I1.REG_15_SQMUXA_275\, B => 
        \I1.REG_16_SQMUXA_94\, Y => 
        \I1.N_41_9_adt_net_3739__net_1\);
    
    \I3.UN7_RONLY_0_A2_0_A3_2638\ : NOR2FT
      port map(A => \I3.WRITES_8\, B => \I3.VASl12r_net_1\, Y => 
        \I3.un7_ronly_0_a2_0_a3_adt_net_165586_\);
    
    \I1.REG_29_sqmuxa_adt_net_855520_\ : BFR
      port map(A => \I1.REG_29_sqmuxa\, Y => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\);
    
    \I3.REG_1_I_S_I_IL4R_1040\ : NOR2
      port map(A => \I3.REG2l4r_net_1\, B => \I3.REG3L4R_432\, Y
         => \I3.N_203_adt_net_24459_\);
    
    \I1.PAGECNTL5R_2876\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_322_adt_net_854384__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL5R_308\);
    
    \I3.REG_1_205\ : MUX2L
      port map(A => VDB_inl24r, B => \I3.REGl157r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\, Y => 
        \I3.REG_1_205_0\);
    
    DTE_padl28r : IOB33PH
      port map(PAD => DTE(28), A => \I2.DTE_1l28r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl28r);
    
    REGl343r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_244_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl343r\);
    
    \I2.PIPE4_DTl0r_1536\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL0R_643\);
    
    \I2.CRC32_12_i_0_m2l10r\ : MUX2L
      port map(A => \I2.DT_TEMPl10r_net_1\, B => 
        \I2.DT_SRAMl10r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854440__net_1\, Y => 
        \I2.N_227_i_i\);
    
    \I2.N_3234_adt_net_855652_\ : BFR
      port map(A => \I2.N_3234\, Y => 
        \I2.N_3234_adt_net_855652__net_1\);
    
    \I5.COMMAND_47\ : MUX2H
      port map(A => \I5.COMMANDl10r_net_1\, B => 
        \I5.COMMAND_4l10r_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.COMMAND_47_net_1\);
    
    \I1.REG_1_181\ : MUX2H
      port map(A => \REGl280r\, B => \I1.REG_74l280r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\, Y => 
        \I1.REG_1_181_net_1\);
    
    VDB_padl26r : IOB33PH
      port map(PAD => VDB(26), A => \I3.VDBml26r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl26r);
    
    \I3.VDBOFFA_31_IV_0L3R_2570\ : AND2
      port map(A => \REGl280r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        Y => \I3.VDBoffa_31l3r_adt_net_164048_\);
    
    \I5.sstate1se_11_i_0_m4\ : MUX2L
      port map(A => \I5.sstate1l2r_net_1\, B => 
        \I5.sstate1l1r_net_1\, S => TICKL0R_558, Y => \I5.N_95\);
    
    \I2.TDCDASl8r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl8r, Q => 
        \I2.TDCDASl8r_net_1\);
    
    REGl322r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_223_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl322r\);
    
    RAMAD_padl2r : OB33PH
      port map(PAD => RAMAD(2), A => RAMAD_cl2r);
    
    VAD_padl21r : OTB33PH
      port map(PAD => VAD(21), A => \I3.VADml21r\, EN => 
        NOEAD_c_i_0);
    
    \I3.REG3l2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_127_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l2r_net_1\);
    
    \I3.VDBoffa_31_iv_0l7r\ : AND2
      port map(A => \REGl212r\, B => 
        \I3.REGMAPl23r_adt_net_855016__net_1\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163264_\);
    
    \I2.PIPE9_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_286_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl17r_net_1\);
    
    \I2.resyn_0_I2_TRGCNT_n2_0\ : XOR2
      port map(A => \I2.TRGCNTl2r_net_1\, B => 
        \I2.un9_tdctrgi_i_0\, Y => \I2.TRGCNT_n2_0\);
    
    \I1.N_1193_adt_net_133987_\ : AO21
      port map(A => \I1.sstatel3r_net_1\, B => REGl90r, C => 
        \I1.sstatel9r_net_1\, Y => 
        \I1.N_1193_adt_net_133987__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I152_Y\ : XOR2FT
      port map(A => \I2.N448_i\, B => 
        \I2.ADD_18x18_fast_I152_Y_0\, Y => \I2.SUB9_1l15r\);
    
    \I2.LEAD_FLAG6_640\ : AO21
      port map(A => \I2.N_4532_adt_net_1157__net_1\, B => 
        \I2.N_4532_adt_net_64252_\, C => 
        \I2.LEAD_FLAG6_640_adt_net_64292_\, Y => 
        \I2.LEAD_FLAG6_640_net_1\);
    
    \I2.majority_reg_i_0l1r\ : OR2
      port map(A => \I2.N_3877_adt_net_4723_\, B => 
        \I2.N_3877_adt_net_4725_\, Y => \I2.N_3877\);
    
    \I2.TRGSERVL1R_2953\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l1r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVL1R_470\);
    
    \I2.PIPE7_DTL27R_2798\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_91\);
    
    \I2.un1_STATE3_12_i\ : OR2
      port map(A => \I2.N_2989_adt_net_92424_\, B => 
        \I2.N_2989_adt_net_92425_\, Y => \I2.N_2989\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__2751\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__27\);
    
    \I3.VDBil12r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_352_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil12r_net_1\);
    
    \I3.VDBi_350\ : MUX2L
      port map(A => \I3.VDBil10r_net_1\, B => \I3.VDBi_57l10r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_350_net_1\);
    
    \I2.DTE_21_1_IV_0L10R_1303\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.DTE_2_1l10r_net_1\, C
         => \I2.DTE_21_1l10r_adt_net_38515_\, Y => 
        \I2.DTE_21_1l10r_adt_net_38526_\);
    
    \I3.VDBi_57l2r_adt_net_145306_\ : AO21
      port map(A => REGl50r, B => \I3.N_2044\, C => 
        \I3.VDBi_57l2r_adt_net_145295__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145306__net_1\);
    
    \I2.CRC32_12_il21r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_58_i_0_i_0\, Y => 
        \I2.N_3938\);
    
    \I2.DTO_16_1_IVL23R_1102\ : AO21
      port map(A => \I2.N_182_adt_net_1007__net_1\, B => 
        \I2.DT_SRAMl23r_net_1\, C => 
        \I2.DTO_16_1l23r_adt_net_30114_\, Y => 
        \I2.DTO_16_1l23r_adt_net_30115_\);
    
    \I3.REG_1l412r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_219_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl412r);
    
    \I2.STATE2l4r_adt_net_855692_\ : BFR
      port map(A => \I2.STATE2l4r_net_1\, Y => 
        \I2.STATE2l4r_adt_net_855692__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I184_Y\ : XOR2FT
      port map(A => \I2.N_40_0\, B => 
        \I2.ADD_21x21_fast_I184_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l14r\);
    
    \I2.OFFSET_37_12l0r\ : MUX2L
      port map(A => \REGl341r\, B => \I2.N_715\, S => 
        \I2.PIPE7_DTL26R_356\, Y => \I2.N_723\);
    
    \I1.REG_74_0_ivl187r\ : AO21
      port map(A => \REGl187r\, B => \I1.N_57_268\, C => 
        \I1.REG_74l187r_adt_net_131699_\, Y => \I1.REG_74l187r\);
    
    \I2.CHA_DATA8\ : DFFC
      port map(CLK => CLK_c, D => \I2.CHA_DATA8_502_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.CHA_DATA8_net_1\);
    
    \I2.OFFSET_37_26l7r\ : MUX2L
      port map(A => \REGl228r\, B => \I2.N_834\, S => 
        \I2.PIPE7_DTL26R_360\, Y => \I2.N_842\);
    
    \I2.REG_1_c1_i_o2\ : AND2
      port map(A => REGL32R_388, B => REGL33R_389, Y => 
        \I2.N_3844\);
    
    \I1.N_50_0_ADT_NET_1409__2871\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__200\, B => 
        \I1.N_50_0_ADT_NET_109751__258\, Y => 
        \I1.N_50_0_ADT_NET_1409__293\);
    
    \I3.VDBOFFB_30_IV_0L0R_2488\ : AO21
      port map(A => \REGl389r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l0r_adt_net_163118_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163125_\);
    
    \I2.PIPE5_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_686_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl10r_net_1\);
    
    \I1.SSTATEL10R_3005\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_43_i_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL10R_759\);
    
    \I3.REG_1_170\ : MUX2L
      port map(A => VDB_inl21r, B => REGl69r, S => 
        \I3.N_1935_adt_net_855320__net_1\, Y => \I3.REG_1_170_0\);
    
    \I1.REG_74_2_i_a2_0l404r\ : OR2FT
      port map(A => \I1.N_232_1_296\, B => 
        \I1.N_1366_adt_net_112007_\, Y => \I1.N_1366\);
    
    \I2.PIPE7_DTL26R_2896\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_350\);
    
    \I3.VDBml6r\ : MUX2L
      port map(A => \I3.VDBil6r_net_1\, B => \I3.N_148\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml6r_net_1\);
    
    \I2.PIPE5_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_700_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl24r_net_1\);
    
    \I2.DTO_16_1l7r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l7r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l7r_Rd1__net_1\);
    
    \I3.REGMAPL31R_3019\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un136_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAPL31R_773\);
    
    \I1.REG_74_0_ivl276r\ : AO21
      port map(A => \REGl276r\, B => 
        \I1.N_145_adt_net_854768__net_1\, C => 
        \I1.REG_74l276r_adt_net_123302_\, Y => 
        \I1.REG_74l276r_net_1\);
    
    MWOK_pad : GL33
      port map(PAD => MWOK, GL => MWOK_c);
    
    \I5.REG_1l435r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_18_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl435r);
    
    \I2.PIPE3_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl2r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I33_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl12r\, B => 
        \I2.PIPE7_DTL12R_693\, Y => \I2.N267_0\);
    
    \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996_\ : 
        BFR
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__net_1\, Y => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996__net_1\);
    
    \I3.VDBml31r\ : MUX2L
      port map(A => \I3.VDBil31r_net_1\, B => \I3.N_173\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml31r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL9R_1471\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\, B => 
        \I2.PIPE1_DT_30l9r_net_1\, C => 
        \I2.PIPE1_DT_42l9r_adt_net_50183_\, Y => 
        \I2.PIPE1_DT_42l9r_adt_net_50199_\);
    
    \I1.BYTECNT_309\ : MUX2H
      port map(A => \I1.BYTECNTl5r_net_1\, B => \I1.N_75\, S => 
        \I1.N_1383_223\, Y => \I1.BYTECNT_309_net_1\);
    
    \I2.BNCID_VECTROR_1427\ : OA21TTF
      port map(A => \I2.BNCID_VECTror_adt_net_48230__net_1\, B
         => \I2.BNCID_VECTror_adt_net_48231__net_1\, C => 
        \I2.TRGSERVL2R_581\, Y => 
        \I2.BNCID_VECTror_adt_net_48463_\);
    
    \I2.EVNT_WORDl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_723_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl10r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I172_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l2r_net_1\, B => 
        \I2.PIPE4_DTL2R_514\, Y => \I2.ADD_21x21_fast_I172_Y_0\);
    
    \I2.CRC32_12_i_0_x2l30r\ : XOR2FT
      port map(A => \I2.CRC32l30r_net_1\, B => \I2.N_231_i_i\, Y
         => \I2.N_245_i_i_0\);
    
    \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Rd1__net_1\);
    
    \I1.sstatel2r\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_289\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel2r_net_1\);
    
    \I1.REG_74_0_iv_i_a3_0l197r\ : OR3FFT
      port map(A => \I1.N_179\, B => \I1.N_145_12\, C => 
        \I1.N_396\, Y => \I1.N_181\);
    
    \I2.SUB9_1_ADD_18x18_fast_I68_Y\ : AOI21
      port map(A => \I2.N302\, B => \I2.N305\, C => \I2.N301_1\, 
        Y => \I2.N336\);
    
    \I2.ADE_4l12r\ : MUX2L
      port map(A => \I2.RPAGEl12r\, B => \I2.WPAGEl12r_net_1\, S
         => NOESRAME_C_243, Y => \I2.ADE_4l12r_net_1\);
    
    \I2.PIPE2_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl25r_net_1\);
    
    RAMDT_padl2r : IOB33PH
      port map(PAD => RAMDT(2), A => \I1.RAMDT_SPI_1l2r_net_1\, 
        EN => \I1.RAMDT_SPI_E_0\, Y => RAMDT_inl2r);
    
    \I2.ADOl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl1r);
    
    \I5.TEMPDATA_81\ : MUX2L
      port map(A => \I5.TEMPDATAl7r_net_1\, B => REGl132r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_81_net_1\);
    
    \I3.REGMAP_I_0_IL45R_2935\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un206_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL45R_452\);
    
    \I3.VDBml29r\ : MUX2L
      port map(A => \I3.VDBil29r_net_1\, B => \I3.N_171\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml29r_net_1\);
    
    \I2.TDCTRGi\ : DFFC
      port map(CLK => CLK_c, D => \I2.TDCTRGi_266_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => TDCTRG_c);
    
    \I1.N_50_0_adt_net_1409__adt_net_855472_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__21\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I34_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl13r\, B => 
        \I2.PIPE7_DTL13R_692\, Y => \I2.N270_0\);
    
    \I3.STATE1_TR24_I_0_A3_5_2112\ : AND3FFT
      port map(A => \I3.REGMAPl13r_net_1\, B => \I3.N_303\, C => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1577__net_1\, Y => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135633_\);
    
    \I1.REG_74_0_IVL235R_1991\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_9_sqmuxa_adt_net_854724__net_1\, Y => 
        \I1.REG_74l235r_adt_net_127194_\);
    
    \I1.REG_19_sqmuxa_adt_net_855488_\ : BFR
      port map(A => \I1.REG_19_sqmuxa\, Y => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\);
    
    \I2.STATE1l0r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1l2r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1l0r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I151_Y_i_o3_3_i\ : AO21
      port map(A => \I2.PIPE4_DTL11R_408\, B => 
        \I2.PIPE4_DTL12R_510\, C => \I2.RAMDT4L12R_144\, Y => 
        \I2.N_20_i_0\);
    
    \I3.MBLTCYC_1161_1737\ : DFFC
      port map(CLK => CLK_c, D => \I3.MBLTCYC_114_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.MBLTCYC_844\);
    
    \I2.SUB9_1_ADD_18x18_fast_I155_Y\ : XOR2FT
      port map(A => \I2.N439_i\, B => 
        \I2.ADD_18x18_fast_I155_Y_0\, Y => \I2.SUB9_1l18r\);
    
    \I2.STATE5_ns_i_0_1l0r\ : AND3FFT
      port map(A => \I2.STATE5_nsl2r\, B => 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1\, C => \I2.N_4332\, Y => 
        \I2.STATE5_ns_i_0_1_il0r\);
    
    REGl363r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_264_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl363r\);
    
    \I2.PIPE6_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_469_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl15r_net_1\);
    
    \I2.FID_417\ : MUX2H
      port map(A => FID_cl1r, B => \I2.FID_7_0_ivl1r_net_1\, S
         => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        Y => \I2.FID_417_net_1\);
    
    \I2.RAMAD1_667\ : MUX2L
      port map(A => \I2.RAMAD1_12l13r_net_1\, B => 
        \I2.RAMAD1l13r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__170\, Y => 
        \I2.RAMAD1_667_net_1\);
    
    \I2.PIPE5_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_703_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl27r_net_1\);
    
    \I2.PIPE1_DTl6r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_733_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl6r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2696\ : AND2
      port map(A => \I2.PIPE4_DTL19R_634\, B => 
        \I2.PIPE4_DTL17R_636\, Y => 
        \I2.N_152_i_0_adt_net_502367_\);
    
    \I2.PIPE7_DTl6r_1592\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL6R_699\);
    
    \I2.PIPE1_DT_42_1_IVL5R_1490\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl21r_net_1\, Y => 
        \I2.PIPE1_DT_42l5r_adt_net_51167_\);
    
    \I3.VDBi_57l6r_adt_net_143308_\ : AND2
      port map(A => REGl412r, B => \I3.REGMAPl55r_net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143308__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I66_Y_1681\ : AND2FT
      port map(A => \I2.LSRAM_OUTl7r\, B => 
        \I2.PIPE7_DTl7r_net_1\, Y => \I2.N316_i_i_adt_net_86577_\);
    
    \I2.PIPE1_DT_42_1_IVL19R_1395\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040__net_1\, 
        B => \I2.PIPE1_DT_12l19r_net_1\, Y => 
        \I2.PIPE1_DT_42l19r_adt_net_47247_\);
    
    \I2.L2TYPEl11r_1555\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_600_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL11R_662\);
    
    \I3.VDBi_344\ : MUX2L
      port map(A => \I3.VDBil4r_net_1\, B => \I3.VDBi_57l4r\, S
         => \I3.un1_STATE1_13_1_adt_net_1351__net_1\, Y => 
        \I3.VDBi_344_net_1\);
    
    \I1.PAGECNTL7R_2979\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_320_adt_net_854868__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL7R_526\);
    
    \I2.DTO_9_IVL11R_1163\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl11r_net_1\, C => 
        \I2.DTO_9l11r_adt_net_32804_\, Y => 
        \I2.DTO_9l11r_adt_net_32812_\);
    
    \I3.VDBi_57_0_iv_0_0l24r\ : OR2
      port map(A => \I3.VDBi_57l24r_adt_net_138814_\, B => 
        \I3.VDBi_57l24r_adt_net_138815_\, Y => \I3.VDBi_57l24r\);
    
    \I1.REG_1_164\ : MUX2H
      port map(A => \REGl263r\, B => \I1.REG_74l263r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y => 
        \I1.REG_1_164_net_1\);
    
    \I2.PIPE3_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl29r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl29r_net_1\);
    
    \I2.ADEl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl1r);
    
    \I1.REG_74_0_IV_0_O2L253R_1828\ : NOR2
      port map(A => \I1.REG_74_0_iv_0_o2_0_il253r\, B => 
        \I1.N_4867_i\, Y => \I1.N_395_adt_net_113232_\);
    
    \I1.REG_74_0_IVL185R_2049\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l185r_adt_net_131871_\);
    
    \I3.RAMAD_VME_24\ : MUX2H
      port map(A => RAMAD_VMEl0r, B => \I3.VASl1r_net_1\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_24_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I57_Y_0_O2_1547\ : AND2
      port map(A => \I2.RAMDT4L1R_769\, B => 
        \I2.PIPE4_DT_I_IL1R_849\, Y => \I2.N357_adt_net_54538_\);
    
    ASB_pad : GL33
      port map(PAD => ASB, GL => ASB_c);
    
    \I2.resyn_0_I2_N_1186_i_i_a2\ : NAND2FT
      port map(A => TDCTRG_C_570, B => \I2.STATE1l17r_net_1\, Y
         => \I2.N_3794\);
    
    \I3.un2_vsel_1_i_0\ : OR2
      port map(A => \I3.ASBS_net_1\, B => 
        \I3.N_1508_adt_net_135122_\, Y => \I3.N_1508\);
    
    \I3.VDBm_0l29r\ : MUX2L
      port map(A => \I3.PIPEAl29r_net_1\, B => 
        \I3.PIPEBl29r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_171\);
    
    \I3.VAS_65\ : MUX2L
      port map(A => VAD_inl3r, B => \I3.VASl3r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_65_net_1\);
    
    \I3.PIPEA_8_0l7r\ : MUX2L
      port map(A => DPR_cl7r, B => \I3.PIPEA1l7r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855352__net_1\, Y => \I3.N_216\);
    
    \I2.PIPE1_DT_42_1_IVL12R_1448\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl28r_net_1\, Y => 
        \I2.PIPE1_DT_42l12r_adt_net_49438_\);
    
    \I1.REG_1_85\ : MUX2H
      port map(A => \REGl184r\, B => \I1.REG_74l184r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, Y => 
        \I1.REG_1_85_net_1\);
    
    \I3.VDBI_57_IV_0_0L2R_2260\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854360__net_1\, B
         => \I3.VDBoffl2r_net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145362_\);
    
    \I3.VDBi_57_0_iv_0l21r\ : OR2
      port map(A => \I3.VDBi_57l21r_adt_net_139188_\, B => 
        \I3.VDBi_57l21r_adt_net_139189_\, Y => \I3.VDBi_57l21r\);
    
    \I2.STATE1l5r_1484\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3214_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1L5R_591\);
    
    \I2.DTO_1_895\ : MUX2L
      port map(A => \I2.DTO_1l21r_Rd1__net_1\, B => 
        \I2.DTO_16_1l21r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834760_Rd1__net_1\, Y
         => \I2.DTO_1l21r\);
    
    \I2.OFFSET_37_18l4r\ : MUX2L
      port map(A => \REGl249r\, B => \REGl185r\, S => 
        \I2.PIPE7_DTL27R_80\, Y => \I2.N_775\);
    
    \I1.REG_74_0_IVL318R_1898\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l318r_adt_net_119217_\);
    
    \I3.REGMAP_I_0_IL58R_3048\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un235_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL58R_802\);
    
    \I3.REG_1l155r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_203_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl155r\);
    
    \I2.PIPE1_DT_42_1_IVL9R_1466\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl25r_net_1\, Y => 
        \I2.PIPE1_DT_42l9r_adt_net_50179_\);
    
    \I0.BNC_RESerr\ : DFFC
      port map(CLK => CLK_c, D => \I0.BNC_RESerr_1_net_1\, CLR
         => \I0.un4_hwresi_i\, Q => BNC_RES_E);
    
    \I2.resyn_0_I2_BITCNT_940\ : MUX2H
      port map(A => \I2.BITCNT_c0\, B => \I2.BITCNT_n0\, S => 
        \I2.BITCNTe\, Y => \I2.BITCNT_940\);
    
    \I2.END_TDC1_1_SQMUXA_I_O2_1015\ : OR3FTT
      port map(A => \I2.TDCGDB1_net_1\, B => \I2.FIRST_TDC_i_0_i\, 
        C => \I2.un2_tdcgdb1_0_adt_net_830__net_1\, Y => 
        \I2.N_3887_adt_net_21865_\);
    
    \I2.resyn_0_I2_TRGCNT_n1_0\ : XOR2
      port map(A => \I2.TRGCNT_i_0_il1r\, B => 
        \I2.un9_tdctrgi_i_0\, Y => \I2.TRGCNT_n1_0\);
    
    \I2.FIDl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_421_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl5r);
    
    DTO_padl7r : IOB33PH
      port map(PAD => DTO(7), A => \I2.DTO_1l7r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl7r);
    
    \I3.VDBI_29L4R_2720\ : AND2FT
      port map(A => \I3.REGMAPL14R_732\, B => 
        \I3.VDBi_20l4r_adt_net_414785_\, Y => 
        \I3.VDBi_29l4r_adt_net_621825_\);
    
    \I2.DT_SRAMl22r\ : MUX2L
      port map(A => \I2.N_890\, B => \I2.PIPE2_DTl22r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668__net_1\, 
        Y => \I2.DT_SRAMl22r_net_1\);
    
    \I1.REG_74_0_ivl268r\ : AO21
      port map(A => \REGl268r\, B => 
        \I1.N_137_adt_net_854760__net_1\, C => 
        \I1.REG_74l268r_adt_net_124027_\, Y => 
        \I1.REG_74l268r_net_1\);
    
    \I1.PAGECNTl9r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854852__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTl9r_net_1\);
    
    \I2.DTO_1l22r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l22r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l22r_Rd1__net_1\);
    
    \I2.LSRAM_INl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_387_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl3r_net_1\);
    
    \I3.EVREAD_DS_1_sqmuxa_1_i_2\ : AND2FT
      port map(A => \I3.ADACKCYC_net_1\, B => 
        \I3.STATE2l1r_net_1\, Y => \I3.N_1860_2\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I164_Y_2653\ : NAND3FTT
      port map(A => \I2.N321_0\, B => \I2.N317\, C => \I2.N411\, 
        Y => \I2.N495_i_adt_net_202093_\);
    
    \I2.un1_STATE3_12_i_o7\ : OR2
      port map(A => \I2.STATE3l0r_net_1\, B => 
        \I2.STATE3l4r_net_1\, Y => \I2.N_4676\);
    
    \I2.PIPE10_DT_17_i_0l17r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855592__net_1\, B => 
        \I2.PIPE9_DTl17r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l17r_net_1\);
    
    \I2.FID_7_0_IVL12R_968\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl60r, C => 
        \I2.FID_7l12r_adt_net_18175_\, Y => 
        \I2.FID_7l12r_adt_net_18183_\);
    
    \I2.CRC32l23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_818_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l23r_net_1\);
    
    INT_ERRB_pad : IB33
      port map(PAD => INT_ERRB, Y => INT_ERRB_c);
    
    \I1.REG_74_0_ivl320r\ : AO21
      port map(A => \REGl320r\, B => \I1.N_193\, C => 
        \I1.REG_74l320r_adt_net_119045_\, Y => \I1.REG_74l320r\);
    
    \I3.PIPEA_244\ : MUX2L
      port map(A => \I3.PIPEAl13r_net_1\, B => 
        \I3.PIPEA_8l13r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854668__net_1\, Y
         => \I3.PIPEA_244_net_1\);
    
    \I1.LUT_0_sqmuxa_i_0_o2_i_0_834_1235\ : NOR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__186\, B
         => \I1.N_325_500\, Y => \I1.N_328_I_0_497\);
    
    \I2.DTO_16_1_ivl1r\ : OA21FTF
      port map(A => \I2.N_182_ADT_NET_1007__386\, B => 
        \I2.DT_SRAMl1r_net_1\, C => \I2.DTO_16_1_iv_1l1r_net_1\, 
        Y => \I2.DTO_16_1_ivl1r_net_1\);
    
    \I1.REG_22_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_267\, B => \I1.N_243\, Y => 
        \I1.REG_22_sqmuxa\);
    
    \I2.OFFSET_37_13l7r\ : MUX2L
      port map(A => \I2.N_730\, B => \I2.N_714\, S => 
        \I2.PIPE7_DTL25R_683\, Y => \I2.N_738\);
    
    \I3.REG_1l96r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_277_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl96r\);
    
    \I2.PIPE5_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_678_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl2r_net_1\);
    
    \I2.EVNT_NUM_c6\ : AND2
      port map(A => \I2.EVNT_NUMl6r_net_1\, B => 
        \I2.EVNT_NUM_c5_net_1\, Y => \I2.EVNT_NUM_c6_net_1\);
    
    REGl255r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_156_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl255r\);
    
    \I3.REG_1_281\ : MUX2H
      port map(A => VDB_inl9r, B => \I3.REGl100r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_281_0\);
    
    REGl258r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_159_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl258r\);
    
    \I2.PIPE1_DT_42_1_ivl12r\ : OR3
      port map(A => \I2.PIPE1_DT_42l12r_adt_net_49448_\, B => 
        \I2.PIPE1_DT_42l12r_adt_net_49457_\, C => 
        \I2.PIPE1_DT_42l12r_adt_net_49458_\, Y => 
        \I2.PIPE1_DT_42l12r\);
    
    \I2.PIPE5_DT_693\ : MUX2L
      port map(A => \I2.PIPE5_DTl17r_net_1\, B => 
        \I2.PIPE5_DT_6l17r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_693_net_1\);
    
    \I3.REG2_147\ : MUX2L
      port map(A => VDB_inl6r, B => \I3.REG2l6r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG2_147_net_1\);
    
    \I2.N_2828_ADT_NET_1062__ADT_NET_835308_RD1__3003\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2828_adt_net_1062__net_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.N_2828_ADT_NET_1062__ADT_NET_835308_RD1__757\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I200_Y\ : XOR2FT
      port map(A => \I2.N411\, B => \I2.SUB_21x21_fast_I200_Y_0\, 
        Y => \I2.SUB8_2l4r\);
    
    \I2.PIPE1_DT_42_1_IVL0R_1525\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, B => 
        \I2.PIPE1_DT_30l0r_net_1\, C => 
        \I2.PIPE1_DT_42l0r_adt_net_52247_\, Y => 
        \I2.PIPE1_DT_42l0r_adt_net_52249_\);
    
    VDB_padl25r : IOB33PH
      port map(PAD => VDB(25), A => \I3.VDBml25r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl25r);
    
    \I3.REG_1_268\ : MUX2H
      port map(A => REGl87r, B => \I3.N_1633\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_268_0\);
    
    \I2.ADOl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl3r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I35_P0N_1285\ : OR2FT
      port map(A => \I2.LSRAM_OUTl14r\, B => 
        \I2.PIPE7_DTl14r_net_1\, Y => \I2.N273_547\);
    
    \I2.OFFSET_37_22l0r\ : MUX2L
      port map(A => \REGl237r\, B => \REGl173r\, S => 
        \I2.PIPE7_DTL27R_76\, Y => \I2.N_803\);
    
    \I1.REG_74_0_iv_0l176r\ : AO21
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, C => 
        \I1.REG_74l176r_adt_net_132682_\, Y => \I1.REG_74l176r\);
    
    \I2.DTE_21_1_IVL23R_1249\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855196__net_1\, 
        B => \I2.DT_TEMPl23r_net_1\, C => 
        \I2.DTO_16_1l23r_adt_net_30106_\, Y => 
        \I2.DTE_21_1l23r_adt_net_37283_\);
    
    \PULSEl0r_adt_net_854536_\ : BFR
      port map(A => PULSEL0R_756, Y => 
        \PULSEl0r_adt_net_854536__net_1\);
    
    \I1.REG_74_0_ivl226r\ : AO21
      port map(A => \REGl226r\, B => \I1.N_97\, C => 
        \I1.REG_74l226r_adt_net_128136_\, Y => \I1.REG_74l226r\);
    
    \I2.DTO_16_1_ivl14r\ : OR2
      port map(A => \I2.DTO_16_1l14r_adt_net_32209_\, B => 
        \I2.DTO_16_1l14r_adt_net_32210_\, Y => \I2.DTO_16_1l14r\);
    
    \I3.RAMDTSl3r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl3r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl3r_net_1\);
    
    \I2.PIPE6_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_481_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl27r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL15R_1431\ : AND2
      port map(A => \I2.BNCID_VECTrxl11r\, B => 
        \I2.PIPE1_DT_42l15r_adt_net_48714_\, Y => 
        \I2.PIPE1_DT_42l15r_adt_net_48707_\);
    
    \I3.TCNT_n0_0_0_a3_1\ : OR2
      port map(A => \I3.REGMAPl51r_net_1\, B => 
        \I3.REG_1_sqmuxa_3\, Y => \I3.N_1966_1\);
    
    \I2.FID_7_0_IVL20R_951\ : AND2
      port map(A => \I2.DTOSl20r_net_1\, B => \I2.STATE3L2R_413\, 
        Y => \I2.FID_7l20r_adt_net_17380_\);
    
    \I2.OFFSETl1r_1573\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_561_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL1R_680\);
    
    \I3.REG_0_sqmuxa_2_adt_net_855300_\ : BFR
      port map(A => \I3.REG_0_sqmuxa_2\, Y => 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\);
    
    \I2.DTO_1_897\ : MUX2L
      port map(A => \I2.DTO_1l23r_Rd1__net_1\, B => 
        \I2.DTO_16_1l23r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834760_Rd1__net_1\, Y
         => \I2.DTO_1l23r\);
    
    \I5.BITCNT_n0_i\ : OA21FTF
      port map(A => \I5.BITCNT_c0\, B => \I5.N_94\, C => 
        \I5.N_144\, Y => \I5.N_50\);
    
    \I2.PIPE1_DT_42_1_IVL18R_1401\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_341\, B => 
        \I2.EVNT_NUMl2r_net_1\, Y => 
        \I2.PIPE1_DT_42l18r_adt_net_47443_\);
    
    \I3.VDBOFFB_30_IV_0L6R_2374\ : AO21
      port map(A => \REGl339r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l6r_adt_net_161938_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161979_\);
    
    \I1.N_1377_adt_net_1517_\ : AO21
      port map(A => \I1.N_310_Rd1__net_1\, B => 
        \I1.PAGECNTl6r_adt_net_854928__net_1\, C => 
        \I1.N_1377_adt_net_106750__net_1\, Y => 
        \I1.N_1377_adt_net_1517__net_1\);
    
    \I4.un1_lead_flag_1_4_0\ : MUX2L
      port map(A => LEAD_FLAGl5r, B => LEAD_FLAGl1r, S => 
        \I4.bcnt_i_0_il2r_net_1\, Y => \I4.N_4\);
    
    \I3.VDBOFFA_31_IV_0L5R_2543\ : OR2
      port map(A => \I3.VDBoffa_31l5r_adt_net_163691_\, B => 
        \I3.VDBoffa_31l5r_adt_net_163692_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163697_\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855444_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__292\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\);
    
    \I2.DTE_21_1_IV_0_0L7R_1316\ : AND2FT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_289\, B => 
        \I2.DT_SRAMl7r_net_1\, Y => 
        \I2.DTE_21_1l7r_adt_net_38863_\);
    
    \I2.PIPE1_DT_42_1_IVL1R_1516\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl33r_net_1\, C => 
        \I2.PIPE1_DT_42l1r_adt_net_52027_\, Y => 
        \I2.PIPE1_DT_42l1r_adt_net_52043_\);
    
    \I2.PIPE1_DT_42_1_IVL19R_1396\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_341\, B => 
        \I2.EVNT_NUMl3r_net_1\, Y => 
        \I2.PIPE1_DT_42l19r_adt_net_47249_\);
    
    \I3.VDBoffa_31_iv_0l5r\ : AND2
      port map(A => \REGl178r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        Y => \I3.VDBoffa_31l5r_adt_net_163644_\);
    
    \I3.REG_1l97r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_278_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl97r\);
    
    \I1.REG_9_sqmuxa_0_a2_1_0_a2_790\ : OR2
      port map(A => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__490\, 
        B => \I1.REG_74_1_380_M8_I_0_RD1__538\, Y => 
        \I1.N_1169_168\);
    
    \I3.RAMAD_VME_35\ : MUX2H
      port map(A => RAMAD_VMEl11r, B => \I3.REGl94r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_35_net_1\);
    
    \I3.VDBI_57_0_IV_0L20R_2167\ : AND2FT
      port map(A => \I3.N_1917_adt_net_855336__net_1\, B => 
        \I3.REGl153r\, Y => \I3.VDBi_57l20r_adt_net_139281_\);
    
    \I2.PIPE6_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_484_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl30r_net_1\);
    
    \I3.PIPEB_110_2316\ : NOR2FT
      port map(A => \I3.PIPEB_i_0_il31r\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_110_adt_net_159411_\);
    
    \I2.BNCID_VECTrff_3_262_0\ : AO21
      port map(A => \I2.BNCID_VECTrff_3_262_0_a2_0\, B => 
        \I2.BNCID_VECTwa15_1_net_1\, C => \I2.BNCID_VECTro_3\, Y
         => \I2.BNCID_VECTrff_3_262_0_net_1\);
    
    \I3.RAMAD_VME_28\ : MUX2H
      port map(A => RAMAD_VMEl4r, B => \I3.VASl5r_net_1\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_28_net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2535\ : AO21
      port map(A => \REGl242r\, B => \I3.REGMAPl27r_net_1\, C => 
        \I3.VDBoffa_31l5r_adt_net_163644_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163688_\);
    
    \I1.N_299_adt_net_833868_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_299_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.N_299_adt_net_833868_Rd1__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I23_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl2r\, B => \I2.PIPE7_DTL2R_702\, 
        Y => \I2.N237_0\);
    
    \I1.REG_74_0_IVL300R_1918\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l300r_adt_net_120868_\);
    
    \I3.VDBOFFB_30_IV_0L1R_2469\ : AO21
      port map(A => \REGl302r\, B => \I3.REGMAPl35r_net_1\, C => 
        \I3.VDBoffb_30l1r_adt_net_162908_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162934_\);
    
    \I3.VDBI_57_0_IVL14R_2190\ : AND2
      port map(A => \I3.PIPEAl14r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l14r_adt_net_140190_\);
    
    \I2.OFFSET_37_2l4r\ : MUX2L
      port map(A => \REGl385r\, B => \REGl321r\, S => 
        \I2.PIPE7_DTL27R_70\, Y => \I2.N_647\);
    
    \I1.REG_74_0_iv_0l262r\ : AO21
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, C => 
        \I1.REG_74l262r_adt_net_124543_\, Y => \I1.REG_74l262r\);
    
    DTO_padl13r : IOB33PH
      port map(PAD => DTO(13), A => \I2.DTO_1l13r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl13r);
    
    \I2.PIPE1_DT_42_1_IV_2L26R_1368\ : NOR2
      port map(A => REGl430r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855816__net_1\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46173_\);
    
    \I3.REG_44_il88r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_1634_adt_net_150223_\, Y => \I3.N_1634\);
    
    \I3.REG3l1r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG3_126_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l1r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I35_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl14r\, B => 
        \I2.PIPE7_DTL14R_691\, Y => \I2.N273\);
    
    \I2.DTO_16_1_IV_0_0L16R_1137\ : AO21
      port map(A => \I2.N_197_153\, B => \I2.DT_SRAMl16r_net_1\, 
        C => \I2.DTO_16_1l16r_adt_net_31708_\, Y => 
        \I2.DTO_16_1l16r_adt_net_31718_\);
    
    \I3.EVREAD_DS_124\ : MUX2H
      port map(A => \I3.EVREAD_DS_net_1\, B => \I3.N_1861\, S => 
        \I3.un1_EVREAD_DS_1_sqmuxa_1_net_1\, Y => 
        \I3.EVREAD_DS_124_net_1\);
    
    \I1.REG_74_0_ivl219r\ : AO21
      port map(A => \REGl219r\, B => \I1.N_89_165\, C => 
        \I1.REG_74l219r_adt_net_128862_\, Y => \I1.REG_74l219r\);
    
    \I2.PIPE1_DT_42_1_IVL4R_1496\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl20r_net_1\, Y => 
        \I2.PIPE1_DT_42l4r_adt_net_51414_\);
    
    \I2.CRC32l22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_817_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l22r_net_1\);
    
    \I1.sstate_tr18_0_a2_0_a4\ : AND2FT
      port map(A => \I1.N_604\, B => 
        \I1.sstate_ns_il5r_adt_net_107266_\, Y => 
        \I1.sstate_ns_il5r\);
    
    \I2.DTO_9_IV_0L31R_1062\ : AND2FT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl31r_net_1\, Y => 
        \I2.DTO_9l31r_adt_net_27894_\);
    
    \I3.PIPEA1l13r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_311_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l13r_net_1\);
    
    \I2.un7_bnc_id_1_I_48\ : AND2
      port map(A => \I2.BNC_IDl7r_net_1\, B => \I2.N_24_1\, Y => 
        \I2.DWACT_FINC_El4r\);
    
    \I1.REG_74_0_IV_0_0L245R_1981\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l245r_adt_net_126207_\);
    
    \I3.REG_1_162\ : MUX2L
      port map(A => VDB_inl13r, B => REGl61r, S => 
        \I3.N_1935_adt_net_855328__net_1\, Y => \I3.REG_1_162_0\);
    
    \I3.REG_0_sqmuxa_2_adt_net_855304_\ : BFR
      port map(A => \I3.REG_0_sqmuxa_2\, Y => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\);
    
    DTE_padl22r : IOB33PH
      port map(PAD => DTE(22), A => \I2.DTE_1l22r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl22r);
    
    \I1.N_310_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_310_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_310_Rd1__net_1\);
    
    REGl209r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_110_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl209r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I24_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl3r\, B => \I2.PIPE7_DTL3R_701\, 
        Y => \I2.N240_0\);
    
    \I2.STATE1l15r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_i_0_il16r\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1_i_0_il15r\);
    
    \I3.REG_1_166\ : MUX2L
      port map(A => VDB_inl17r, B => REGl65r, S => 
        \I3.N_1935_adt_net_855324__net_1\, Y => \I3.REG_1_166_0\);
    
    FID_padl28r : OB33PH
      port map(PAD => FID(28), A => FID_cl28r);
    
    \I2.TDCDASl13r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl13r, Q => 
        \I2.TDCDASl13r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I138_Y_0_a2_0_2\ : OAI21
      port map(A => \I2.PIPE4_DTL10R_850\, B => 
        \I2.PIPE4_DTL9R_845\, C => \I2.RAMDT4L5R_813\, Y => 
        \I2.N_112_2\);
    
    \I3.UN1_STATE2_15_1_ADT_NET_1342__2856\ : OR2
      port map(A => \I3.STATE2_nsl0r_adt_net_136048_\, B => 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\, Y => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854680_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854680__net_1\);
    
    \I2.PIPE7_DTl25r_1574\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL25R_681\);
    
    \I3.TCNT4_i_0_il2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT4_386_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT4_i_0_il2r_net_1\);
    
    \I1.REG_74_0_ivl349r\ : AO21
      port map(A => \REGl349r\, B => \I1.N_225\, C => 
        \I1.REG_74l349r_adt_net_116203_\, Y => \I1.REG_74l349r\);
    
    \I2.EVNT_NUM_n6\ : NOR2
      port map(A => EV_RES_c, B => \I2.EVNT_NUM_n6_tz_i\, Y => 
        \I2.EVNT_NUM_n6_net_1\);
    
    \I3.REG2l405r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG2_228_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l405r_net_1\);
    
    \I2.PIPE4_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl31r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl31r_net_1\);
    
    \I2.DTE_21_1_IV_0L19R_1264\ : AND2
      port map(A => \I2.DT_SRAMl19r_net_1\, B => 
        \I2.N_199_0_ADT_NET_1054__36\, Y => 
        \I2.DTE_21_1l19r_adt_net_37713_\);
    
    \I2.EVNT_NUM_n4_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl4r_net_1\, B => 
        \I2.EVNT_NUM_c3_net_1\, Y => \I2.EVNT_NUM_n4_tz_i\);
    
    \I2.RAMAD1_668\ : MUX2L
      port map(A => \I2.RAMAD1_12l14r_net_1\, B => 
        \I2.RAMAD1l14r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__170\, Y => 
        \I2.RAMAD1_668_net_1\);
    
    \I1.REG_74_0_IVL401R_1788\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_30_sqmuxa_adt_net_854376__net_1\, Y => 
        \I1.REG_74l401r_adt_net_110014_\);
    
    \I2.PIPE2_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl28r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl28r_net_1\);
    
    \I2.DTO_16_1_IV_0_0L26R_1083\ : AND2
      port map(A => \I2.DTO_1l26r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l26r_adt_net_29428_\);
    
    \I3.TCNT2_395\ : MUX2H
      port map(A => \I3.TCNT2l1r_net_1\, B => \I3.TCNT2_n1_net_1\, 
        S => TICKl0r, Y => \I3.TCNT2_395_net_1\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_adt_net_803__net_1\, Y
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\);
    
    \I2.DTO_16_1_IV_0L20R_1117\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855676__net_1\, B => 
        \I2.DTO_9l20r\, Y => \I2.DTO_16_1l20r_adt_net_30778_\);
    
    \I3.VDBi_20_ivl10r\ : AO21
      port map(A => \I3.VDBi_20l12r_adt_net_140770_\, B => 
        \I3.N_2261\, C => \I3.VDBi_20l10r_adt_net_141609_\, Y => 
        \I3.VDBi_20l10r\);
    
    \I3.UN12_TCNT3_2640\ : NOR2
      port map(A => \I3.TCNT3_i_0_il0r_net_1\, B => 
        \I3.TCNT3l7r_net_1\, Y => \I3.un12_tcnt3_adt_net_165616_\);
    
    \I2.DTO_16_1_IVL22R_1109\ : AO21
      port map(A => \I2.N_182_adt_net_1007__net_1\, B => 
        \I2.DT_SRAMl22r_net_1\, C => 
        \I2.DTO_16_1l22r_adt_net_30360_\, Y => 
        \I2.DTO_16_1l22r_adt_net_30361_\);
    
    \I2.LSRAM_IN_399\ : MUX2L
      port map(A => \I2.PIPE5_DTl15r_net_1\, B => 
        \I2.LSRAM_INl15r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_399_net_1\);
    
    \I2.un78_pipe5_dt_3\ : XOR2
      port map(A => \I2.un78_pipe5_dt_1_net_1\, B => 
        \I2.un78_pipe5_dt_0_net_1\, Y => 
        \I2.un78_pipe5_dt_3_net_1\);
    
    \I2.PIPE8_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_540_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl12r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2555\ : AO21
      port map(A => \REGl225r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.VDBoffa_31l4r_adt_net_163842_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163880_\);
    
    \I3.VDBOFFB_30_IV_0L1R_2472\ : OR3
      port map(A => \I3.VDBoffb_30l1r_adt_net_162935_\, B => 
        \I3.VDBoffb_30l1r_adt_net_162929_\, C => 
        \I3.VDBoffb_30l1r_adt_net_162930_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162939_\);
    
    NPRSFIF_pad : OB33PH
      port map(PAD => NPRSFIF, A => NMRSFIF_c_c);
    
    \I2.PIPE5_DT_6_0l15r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l15r\, B => 
        \I2.un27_pipe5_dt0l15r\, S => 
        \I2.dataout_0_adt_net_855804__net_1\, Y => \I2.N_1084\);
    
    \I2.CRC32l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_798_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l3r_net_1\);
    
    \I1.BYTECNTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_311_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTl3r_net_1\);
    
    \I2.LSRAM_INl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_410_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl26r_net_1\);
    
    DPR_padl19r : IB33
      port map(PAD => DPR(19), Y => DPR_cl19r);
    
    \I3.VDBi_57_0_iv_0l27r\ : OR2
      port map(A => \I3.VDBi_57l27r_adt_net_138440_\, B => 
        \I3.VDBi_57l27r_adt_net_138441_\, Y => \I3.VDBi_57l27r\);
    
    \I3.REG_1_158\ : MUX2L
      port map(A => VDB_inl9r, B => REGl57r, S => 
        \I3.N_1935_adt_net_855328__net_1\, Y => \I3.REG_1_158_0\);
    
    \I2.SUB8l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_508_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l5r_net_1\);
    
    \I2.SRAM_EVNT_C2_I_1747\ : NOR2
      port map(A => \I2.N_3858\, B => \I2.N_128_1\, Y => 
        \I2.N_3827_adt_net_101792_\);
    
    \I2.OFFSET_37_28l4r\ : MUX2L
      port map(A => \I2.N_847\, B => \I2.N_799\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_855\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0_o2_1_726\ : OR2
      port map(A => \I2.N_128_0\, B => 
        \I2.N_74_ADT_NET_55281__326\, Y => \I2.N_74_104\);
    
    \I2.L2SERV_920\ : MUX2H
      port map(A => \I2.RPAGEl14r\, B => \I2.L2SERV_n2_net_1\, S
         => \I2.L2SERVe\, Y => \I2.L2SERV_920_net_1\);
    
    \I2.DTE_1_847\ : MUX2L
      port map(A => \I2.DTE_1l7r_Rd1__net_1\, B => 
        \I2.DTE_21_1l7r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, Y => 
        \I2.DTE_1l7r\);
    
    REGl323r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_224_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl323r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I91_Y_0_a4\ : AND2FT
      port map(A => \I2.N_28_0\, B => 
        \I2.N_2358_tz_tz_adt_net_854956__net_1\, Y => \I2.N_93_0\);
    
    \I2.MIC_REG2_312_adt_net_855644_\ : BFR
      port map(A => \I2.MIC_REG2_312_net_1\, Y => 
        \I2.MIC_REG2_312_adt_net_855644__net_1\);
    
    \I3.VDBOFFB_30_IV_0L0R_2480\ : AND2
      port map(A => \REGl301r\, B => \I3.REGMAPl35r_net_1\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163098_\);
    
    \I2.un1_STATE1_22_1\ : AO21FTT
      port map(A => \I2.N_3272_345\, B => \I2.N_3277\, C => 
        \I2.STATE1l13r_net_1\, Y => \I2.un1_STATE1_22\);
    
    REGl301r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_202_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl301r\);
    
    \I3.VDBi_57l2r_adt_net_145295_\ : AND3FFT
      port map(A => \I3.N_2017\, B => 
        \I3.REGMAPl9r_adt_net_854324__net_1\, C => 
        \I3.VDBi_57l2r_adt_net_1614__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145295__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I33_Y\ : AO21TTF
      port map(A => \I2.SUB8l11r_adt_net_855580__net_1\, B => 
        \I2.SUB8l12r_net_1\, C => \I2.N295_adt_net_68996_\, Y => 
        \I2.N298\);
    
    \I2.DTESl4r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl4r, Q => 
        \I2.DTESl4r_net_1\);
    
    \I1.REG_1_112\ : MUX2H
      port map(A => \REGl211r\, B => \I1.N_144\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_112_net_1\);
    
    REGl190r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_91_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl190r\);
    
    \I1.REG_74_0_iv_i_a2l204r\ : AO21
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\, C => 
        \I1.N_1343_adt_net_130189_\, Y => \I1.N_1343\);
    
    \I1.REG_74_0_ivl379r\ : AO21
      port map(A => \REGl379r\, B => \I1.N_249\, C => 
        \I1.REG_74l379r_adt_net_112571_\, Y => \I1.REG_74l379r\);
    
    \I5.sstate1l7r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el6r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l7r_net_1\);
    
    \I2.ADO_3l4r\ : MUX2L
      port map(A => \I2.WOFFSETl5r\, B => \I2.ROFFSETl5r_net_1\, 
        S => NOESRAME_C_243, Y => \I2.ADO_3l4r_net_1\);
    
    \I1.REG_74_0_IVL261R_1962\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, Y => 
        \I1.REG_74l261r_adt_net_124629_\);
    
    \I2.WPAGE_c2\ : NAND2
      port map(A => \I2.WPAGEl14r_net_1\, B => 
        \I2.WPAGE_c1_net_1\, Y => \I2.WPAGE_c2_net_1\);
    
    \I2.DTE_1_856\ : MUX2L
      port map(A => \I2.DTE_1l16r_Rd1__net_1\, B => 
        \I2.DTE_21_1l16r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\, Y => 
        \I2.DTE_1l16r\);
    
    \I1.BITCNT_n2_i_i_m4\ : AO21TTF
      port map(A => \I1.N_1376_i_0\, B => \I1.N_389_i_i_0\, C => 
        \I1.N_604\, Y => \I1.N_415\);
    
    \I2.LSRAM_IN_385\ : MUX2L
      port map(A => \I2.PIPE5_DTl1r_net_1\, B => 
        \I2.LSRAM_INl1r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_385_net_1\);
    
    \I2.PIPE9_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_284_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl15r_net_1\);
    
    \I2.N_4090_i_0_m2\ : MUX2L
      port map(A => \I2.PIPE10_DTl18r_net_1\, B => 
        \I2.PIPE5_DTl18r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854224__net_1\, Y => 
        \I2.N_202_i\);
    
    \I2.CRC32_12_i_0_m2l27r\ : OAI21TTF
      port map(A => \I2.N_4647\, B => 
        \I2.N_4667_1_adt_net_1046__adt_net_854436__net_1\, C => 
        \I2.N_230_i_i_adt_net_41076_\, Y => \I2.N_230_i_i\);
    
    \I2.ADO_3l8r\ : MUX2L
      port map(A => \I2.WOFFSETl9r\, B => \I2.ROFFSETl9r_net_1\, 
        S => NOESRAME_C_243, Y => \I2.ADO_3l8r_net_1\);
    
    REGl347r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_248_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl347r\);
    
    \I2.OFFSET_37_2l0r\ : MUX2L
      port map(A => \REGl381r\, B => \REGl317r\, S => 
        \I2.PIPE7_DTL27R_74\, Y => \I2.N_643\);
    
    \I2.OFFSET_37_23l7r\ : MUX2L
      port map(A => \REGl276r\, B => \REGl212r\, S => 
        \I2.PIPE7_DTL27R_87\, Y => \I2.N_818\);
    
    \I3.TCNT2_392\ : MUX2H
      port map(A => \I3.TCNT2_i_0_il4r_net_1\, B => 
        \I3.TCNT2_n4_net_1\, S => TICKl0r, Y => 
        \I3.TCNT2_392_net_1\);
    
    \I1.REG_74_0_IV_0L360R_1847\ : AND2
      port map(A => \FBOUTl3r\, B => \I1.REG_25_sqmuxa\, Y => 
        \I1.REG_74l360r_adt_net_114869_\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2515\ : AND2
      port map(A => \REGl275r\, B => \I3.REGMAPl31r_net_1\, Y => 
        \I3.N_2070_adt_net_163474_\);
    
    \I2.SUB8l20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_523_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l20r_net_1\);
    
    \I1.REG_74_0_iv_0l365r\ : AO21
      port map(A => \REGl365r\, B => \I1.N_660\, C => 
        \I1.REG_74l365r_adt_net_113912_\, Y => \I1.REG_74l365r\);
    
    \I3.un5_noemic_0_a2_i\ : NAND3
      port map(A => \I3.LWORDS_net_1\, B => \I3.N_277\, C => 
        \I3.REGMAPl10r_net_1\, Y => NOEMIC_c);
    
    \I1.REG_74_0_IV_0L180R_2054\ : AND2
      port map(A => \REGl180r\, B => \I1.N_49_267\, Y => 
        \I1.REG_74l180r_adt_net_132338_\);
    
    \I3.VDBi_341\ : MUX2L
      port map(A => \I3.VDBil1r_net_1\, B => \I3.VDBi_57l1r\, S
         => \I3.un1_STATE1_13_1_adt_net_1351__net_1\, Y => 
        \I3.VDBi_341_net_1\);
    
    \I3.PIPEB_104\ : AO21
      port map(A => DPR_cl25r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\, 
        C => \I3.PIPEB_104_adt_net_159663_\, Y => 
        \I3.PIPEB_104_net_1\);
    
    \I2.L2TYPE_4_IL9R_1626\ : AND2
      port map(A => \I2.L2TYPE_i_0_il9r\, B => 
        \I2.N_4443_adt_net_67572_\, Y => 
        \I2.N_4443_adt_net_67615_\);
    
    \I3.un6_tcnt1\ : AND3FFT
      port map(A => \I3.TCNT1l2r_net_1\, B => \I3.TCNT1l0r_net_1\, 
        C => \I3.un6_tcnt1_adt_net_134944_\, Y => 
        \I3.un6_tcnt1_net_1\);
    
    \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844_\ : BFR
      port map(A => \I2.MIC_REG1_1_sqmuxa_0\, Y => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\);
    
    \I3.REG_1_189\ : MUX2L
      port map(A => VDB_inl8r, B => \I3.REGl141r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, Y => 
        \I3.REG_1_189_0\);
    
    \I1.REG_74_0_IV_0L367R_1834\ : AND2
      port map(A => \FBOUTl2r\, B => \I1.N_593\, Y => 
        \I1.REG_74l367r_adt_net_113740_\);
    
    \I2.SUB8_1_sqmuxa_0_adt_net_855152_\ : BFR
      port map(A => \I2.SUB8_1_sqmuxa_0\, Y => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855152__net_1\);
    
    \I2.MIC_ERR_REGSl40r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_369_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl40r_net_1\);
    
    \I2.DTO_1_889\ : MUX2L
      port map(A => \I2.DTO_1l15r_Rd1__net_1\, B => 
        \I2.DTO_16_1l15r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834768_Rd1__net_1\, Y
         => \I2.DTO_1l15r\);
    
    \I5.COMMAND_51\ : MUX2H
      port map(A => \I5.COMMANDl14r_net_1\, B => 
        \I5.COMMAND_4l14r_net_1\, S => \I5.sstate1l13r_net_1\, Y
         => \I5.COMMAND_51_net_1\);
    
    \I2.FID_7_0_IVL17R_958\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl65r, C => 
        \I2.FID_7l17r_adt_net_17705_\, Y => 
        \I2.FID_7l17r_adt_net_17713_\);
    
    \I1.REG_74_13_388_m8_i_a4\ : NOR3
      port map(A => \I1.PAGECNTl6r_adt_net_854924__net_1\, B => 
        \I1.PAGECNTl5r_net_1\, C => 
        \I1.REG_74_12_300_N_13_Rd1__net_1\, Y => 
        \I1.REG_74_13_388_N_16_adt_net_109531_\);
    
    \I3.VDBOFFB_30_IV_0L3R_2432\ : AO21
      port map(A => \REGl312r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        C => \I3.VDBoffb_30l3r_adt_net_162524_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162553_\);
    
    \I1.REG_74_12_348_m9_i\ : OR3FTT
      port map(A => \I1.N_232_1\, B => 
        \I1.REG_74_12_348_m9_i_adt_net_115422_\, C => 
        \I1.REG_74_12_348_m9_i_adt_net_115430_\, Y => 
        \I1.REG_74_12_348_m9_i_net_1\);
    
    \I1.REG_74_5_404_m1_e_0\ : NOR2FT
      port map(A => \I1.PAGECNT_0l8r_adt_net_834720_Rd1__net_1\, 
        B => \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__362\, Y => 
        \I1.REG_74_5_404_m1_e_0_net_1\);
    
    \I1.N_223_adt_net_854844_\ : BFR
      port map(A => \I1.N_223\, Y => 
        \I1.N_223_adt_net_854844__net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__3078\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__832\);
    
    \I2.RAMAD_4_0l1r\ : MUX2H
      port map(A => \I2.RAMAD1l1r_net_1\, B => RAMAD_VMEl1r, S
         => \REG_i_il5r_adt_net_855560__net_1\, Y => \I2.N_528\);
    
    \I2.DT_TEMP_786\ : MUX2H
      port map(A => \I2.DT_TEMPl25r_net_1\, B => 
        \I2.DT_TEMP_7l25r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_786_net_1\);
    
    REGl300r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_201_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl300r\);
    
    \I3.VDBI_57_0_IVL14R_2191\ : AND3FTT
      port map(A => \I3.N_1905_1_adt_net_855384__net_1\, B => 
        \I3.N_354_0_adt_net_855368__net_1\, C => \I3.N_352\, Y
         => \I3.VDBi_57l14r_adt_net_140192_\);
    
    \I2.I_1342_G_1\ : XOR2FT
      port map(A => \I2.SUB8l10r_net_1\, B => \I2.OFFSETL7R_671\, 
        Y => \I2.G_1\);
    
    \I2.un7_bnc_id_1_I_55\ : AND2
      port map(A => \I2.N_14\, B => \I2.BNC_IDl9r_net_1\, Y => 
        \I2.N_11_1\);
    
    \I2.STATE3l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl6r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3l7r_net_1\);
    
    \I3.REG_1l115r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_296_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl115r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I202_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl6r\, B => 
        \I2.PIPE7_DTl6r_net_1\, Y => \I2.SUB_21x21_fast_I202_Y_0\);
    
    \I2.OFFSET_37_14l5r\ : MUX2L
      port map(A => \I2.N_736\, B => \I2.N_688\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_744\);
    
    \I1.SBYTE_8_I_0L7R_1755\ : OA21TTF
      port map(A => \I1.N_603_i\, B => \FBOUTl6r\, C => 
        \I1.N_337\, Y => \I1.N_1194_adt_net_106064_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2697\ : OA21
      port map(A => \I2.RAMDT4L12R_829\, B => 
        \I2.N_152_i_0_adt_net_502367_\, C => 
        \I2.ADD_21x21_fast_I140_Y_0_a2_0_0_0\, Y => 
        \I2.N_152_i_0_adt_net_502543_\);
    
    RAMAD_padl7r : OB33PH
      port map(PAD => RAMAD(7), A => RAMAD_cl7r);
    
    \I3.VDBOFFB_30_IV_0L4R_2415\ : AO21
      port map(A => \REGl337r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l4r_adt_net_162338_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162364_\);
    
    \I3.N_1463_i_adt_net_1279_\ : OR2
      port map(A => \I3.EVREAD_DS_729\, B => \I3.N_1896\, Y => 
        \I3.N_1463_i_adt_net_1279__net_1\);
    
    \I2.UN1_STATE1_39_6_1530\ : OAI21FTF
      port map(A => \I2.TDCGDA1_net_1\, B => \I2.STATE1_ns_1l7r\, 
        C => \I2.un1_STATE1_39_6_i_adt_net_52471_\, Y => 
        \I2.un1_STATE1_39_6_i_adt_net_52473_\);
    
    \I2.CRC32_12_il28r\ : NOR2
      port map(A => \I2.N_2867_1_adt_net_854964__net_1\, B => 
        \I2.N_19_i_0_i_0\, Y => \I2.N_3945\);
    
    \I5.sstate1se_7_0_0_o4\ : NAND2
      port map(A => \I5.BITCNTl2r_net_1\, B => \I5.N_65\, Y => 
        \I5.N_67\);
    
    \I3.PIPEA1_12l17r\ : AND2
      port map(A => DPR_cl17r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854500__net_1\, Y => 
        \I3.PIPEA1_12l17r_net_1\);
    
    \I2.DT_TEMP_788\ : MUX2H
      port map(A => \I2.DT_TEMPl27r_net_1\, B => 
        \I2.DT_TEMP_7l27r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_788_net_1\);
    
    \I2.CRC32l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_795_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l0r_net_1\);
    
    \I3.VDBi_40_sn_m2_0\ : NOR2
      port map(A => \I3.REGMAPL57R_807\, B => 
        \I3.REGMAP_I_0_IL58R_802\, Y => \I3.N_354_0\);
    
    \I2.DTE_2_1_0l11r\ : XOR2
      port map(A => \I2.CRC32l19r_net_1\, B => 
        \I2.CRC32l7r_net_1\, Y => \I2.DTE_2_1_0l11r_net_1\);
    
    \I2.PIPE7_DTl25r_1579\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL25R_686\);
    
    \I5.DATAl10r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l10r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl127r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I176_Y\ : AND2FT
      port map(A => \I2.LSRAM_OUTl19r\, B => 
        \I2.PIPE7_DTl19r_net_1\, Y => \I2.N475_adt_net_87372_\);
    
    \I1.REG_74_0_IVL391R_1799\ : NOR2FT
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, Y => 
        \I1.REG_74l391r_adt_net_110956_\);
    
    \I2.BNCID_VECT_tile_DOUTl4r\ : MUX2L
      port map(A => \I2.DIN_REG1l4r\, B => \I2.DOUT_TMPl4r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl4r\);
    
    \I2.BNCID_VECT_tile_DOUTl6r\ : MUX2L
      port map(A => \I2.DIN_REG1l6r\, B => \I2.DOUT_TMPl6r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl6r\);
    
    \I3.EVREADi_1125\ : DFFC
      port map(CLK => CLK_c, D => \I3.EVREADi_225_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => EVREAD_387);
    
    \I1.BITCNTlde_i_a2_0_o2_0\ : OR2
      port map(A => \I1.sstate_nsl4r\, B => \I1.sstate_nsl6r\, Y
         => \I1.N_349_Ra1_\);
    
    \I1.PAGECNTl6r_adt_net_854932_\ : BFR
      port map(A => \I1.PAGECNTl6r_net_1\, Y => 
        \I1.PAGECNTl6r_adt_net_854932__net_1\);
    
    \I3.TCNT3_n5\ : XOR2
      port map(A => \I3.TCNT3l5r_net_1\, B => \I3.TCNT3_c4\, Y
         => \I3.TCNT3_n5_net_1\);
    
    \I2.PIPE1_DT_42_1_iv_2l27r\ : OR2
      port map(A => \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46038_\, 
        B => \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46039_\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il27r\);
    
    \I3.STATE1_ns_0_iv_0l1r\ : OR2
      port map(A => \I3.STATE1_nsl1r_adt_net_134332_\, B => 
        \I3.STATE1_nsl1r_adt_net_134337_\, Y => \I3.STATE1_nsl1r\);
    
    \I5.SDAnoe_83\ : MUX2H
      port map(A => \I5.SDAnoe_net_1\, B => \I5.SDAnoe_8\, S => 
        TICKL0R_3, Y => \I5.SDAnoe_83_net_1\);
    
    \I3.VDBOFFB_30_IV_0L7R_2362\ : AO21
      port map(A => \REGl396r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l7r_adt_net_161788_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161795_\);
    
    \I3.REGMAPL22R_3021\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un91_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL22R_775\);
    
    \I1.REG_74_0_ivl302r\ : AO21
      port map(A => \REGl302r\, B => \I1.N_177\, C => 
        \I1.REG_74l302r_adt_net_120696_\, Y => \I1.REG_74l302r\);
    
    \I3.VDBoffb_30_iv_0_0l5r\ : AND2
      port map(A => \REGl370r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162124_\);
    
    \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149_\ : NOR3FFT
      port map(A => \I2.END_EVNT5_405\, B => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\, C => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_M3_237\, Y => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149__net_1\);
    
    \I3.VDBI_57_0_IVL16R_2182\ : AO21
      port map(A => \I3.VDBil16r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l16r_adt_net_139761_\, Y => 
        \I3.VDBi_57l16r_adt_net_139767_\);
    
    \I3.REG2l3r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG2_144_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l3r_net_1\);
    
    \I3.PULSE_334\ : MUX2L
      port map(A => PULSEL4R_15, B => \I3.N_55\, S => 
        \I3.N_1409_adt_net_854744__net_1\, Y => 
        \I3.PULSE_334_net_1\);
    
    \I2.TOKINAi_325\ : OA21TTF
      port map(A => TOKINA_c, B => \I2.STATE1l13r_net_1\, C => 
        \I2.STATE1l12r_adt_net_855176__net_1\, Y => 
        \I2.TOKINAi_325_net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_45410_\ : OAI21TTF
      port map(A => \I2.TDCGDA1_net_1\, B => 
        \I2.NWPIPE1_4_sqmuxa_1_0\, C => 
        \I2.un1_STATE1_40_1_adt_net_45381__net_1\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45410__net_1\);
    
    \I1.REG_74_0_IVL182R_2052\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l182r_adt_net_132129_\);
    
    \I1.BITCNT_n1_i_i_x2\ : XOR2
      port map(A => \I1.BITCNTl0r_net_1\, B => 
        \I1.BITCNTl1r_net_1\, Y => \I1.N_387_i_0\);
    
    \I3.VDBOFFA_51_2510\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal7r_net_1\, Y => 
        \I3.VDBoffa_51_adt_net_163358_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I114_Y\ : NOR3
      port map(A => \I2.N332\, B => \I2.I94_un1_Y\, C => 
        \I2.I114_un1_Y\, Y => \I2.N454_i\);
    
    \I3.VASl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_66_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl4r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I172_Y\ : XOR2
      port map(A => \I2.N357\, B => \I2.ADD_21x21_fast_I172_Y_0\, 
        Y => \I2.un27_pipe5_dt0l2r\);
    
    \I1.REG_1_249\ : MUX2H
      port map(A => \REGl348r\, B => \I1.REG_74l348r_net_1\, S
         => \I1.N_50_0_ADT_NET_1409__20\, Y => 
        \I1.REG_1_249_net_1\);
    
    \I2.WOFFSETl1r_adt_net_854992_\ : BFR
      port map(A => \I2.WOFFSETl1r\, Y => 
        \I2.WOFFSETl1r_adt_net_854992__net_1\);
    
    \I2.DTOSl3r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl3r, Q => 
        \I2.DTOSl3r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2429\ : AO21
      port map(A => \REGl384r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l3r_adt_net_162512_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162550_\);
    
    \I2.EVNT_NUMl8r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_955_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl8r_net_1\);
    
    N_1_I3_TCNT2_c5 : AND2
      port map(A => \I3.TCNT2l5r_net_1\, B => \I3.TCNT2_c4\, Y
         => \N_1.I3.TCNT2_c5\);
    
    \I2.ROFFSET_n3_tz\ : XOR2FT
      port map(A => \I2.ROFFSETl3r_net_1\, B => 
        \I2.ROFFSET_c2_net_1\, Y => \I2.ROFFSET_n3_tz_i\);
    
    \I2.FID_7_IVL3R_1727\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl51r, C => 
        \I2.STATE3l9r_net_1\, Y => \I2.FID_7l3r_adt_net_93258_\);
    
    \I3.REG_1l83r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_264_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl83r);
    
    \I2.TRGSERVl1r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l1r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVl1r_net_1\);
    
    \I3.un1_singcyc8_i_0\ : AO21
      port map(A => \I3.N_1918\, B => \I3.STATE1_ipl5r\, C => 
        \I3.N_80\, Y => \I3.N_1509\);
    
    \I3.PIPEA_238\ : MUX2L
      port map(A => \I3.PIPEAl7r_net_1\, B => 
        \I3.PIPEA_8l7r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854676__net_1\, Y
         => \I3.PIPEA_238_net_1\);
    
    \I2.DTO_16_1_IV_0L28R_1075\ : NOR2
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608__net_1\, 
        B => \I2.DT_TEMPl28r_net_1\, Y => 
        \I2.DTO_16_1_iv_0l28r_adt_net_28950_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I25_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl4r\, B => 
        \I2.PIPE7_DTl4r_net_1\, Y => \I2.N243_0\);
    
    \I2.majority_reg_i_0l2r\ : OAI21TTF
      port map(A => \I2.MIC_REG3L2R_789\, B => 
        \I2.MIC_REG1L2R_464\, C => \I2.N_3876_adt_net_4861_\, Y
         => \I2.N_3876\);
    
    \I2.DTE_cl_0_sqmuxa_2_0_a2_0_a2_0_909\ : OR2FT
      port map(A => \I2.N_4241_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, Y => 
        \I2.DTE_CL_0_SQMUXA_2_0_287\);
    
    \I2.DTE_21_1l28r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l28r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l28r_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2541\ : AO21
      port map(A => \REGl266r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        C => \I3.VDBoffa_31l5r_adt_net_163668_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163694_\);
    
    TDCDB_padl28r : IB33
      port map(PAD => TDCDB(28), Y => TDCDB_cl28r);
    
    \I2.SUB9_1_ADD_18x18_fast_I124_Y\ : AO21
      port map(A => \I2.N284\, B => \I2.N434_adt_net_69748_\, C
         => \I2.N434_adt_net_69831_\, Y => \I2.N434\);
    
    REGl367r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_268_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl367r\);
    
    \I2.PIPE1_DT_12l18r\ : MUX2L
      port map(A => \I2.TDCDASl18r_net_1\, B => 
        \I2.TDCDASl16r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, Y
         => \I2.PIPE1_DT_12l18r_net_1\);
    
    REGl182r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_83_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl182r\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I178_Y_2704\ : NAND3FTT
      port map(A => \I2.N479_adt_net_296182__net_1\, B => 
        \I2.N501_i_adt_net_88539_\, C => \I2.N355_0\, Y => 
        \I2.N479_adt_net_538220_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I204_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl8r\, B => 
        \I2.PIPE7_DTl8r_net_1\, Y => \I2.SUB_21x21_fast_I204_Y_0\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_a2_1\ : NAND3FFT
      port map(A => \I2.RAMDT4l10r_net_1\, B => 
        \I2.PIPE4_DTl3r_adt_net_854544__net_1\, C => \I2.N_67\, Y
         => \I2.N_107_0_adt_net_320361_\);
    
    \I1.REG_74_0_ivl189r\ : AO21
      port map(A => \REGl189r\, B => \I1.N_65\, C => 
        \I1.REG_74l189r_adt_net_131527_\, Y => \I1.REG_74l189r\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__2835\ : NOR3FFT
      port map(A => \I2.END_EVNT5_406\, B => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\, C => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m3_net_1\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__184\);
    
    \I2.PIPE1_DT_42_1_IVL10R_1460\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl26r_net_1\, Y => 
        \I2.PIPE1_DT_42l10r_adt_net_49932_\);
    
    \I3.PIPEB_4l30r\ : NAND2FT
      port map(A => DPR_cl30r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855280__net_1\, 
        Y => \I3.PIPEB_4l30r_net_1\);
    
    \I2.RAMDT4L10R_3012\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl10r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L10R_766\);
    
    \I2.PIPE4_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl7r_net_1\);
    
    \I2.DTO_9_ivl15r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl15r_net_1\, 
        C => \I2.DTO_9l15r_adt_net_31896_\, Y => \I2.DTO_9l15r\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I137_Y_I_2707\ : OR3FFT
      port map(A => \I2.N_59_0\, B => \I2.N_96_0_adt_net_469923_\, 
        C => \I2.N522_0_adt_net_329219_\, Y => 
        \I2.N_40_0_adt_net_577252_\);
    
    \I1.REG_74_0_iv_0_o2l372r\ : NAND3FFT
      port map(A => \I1.N_396\, B => \I1.N_395\, C => 
        \I1.REG_74_i_o2_i_0l364r_net_1\, Y => \I1.N_660\);
    
    \I2.PIPE9_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_280_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl11r_net_1\);
    
    \I2.DTO_1_898\ : MUX2L
      port map(A => \I2.DTO_1l24r_Rd1__net_1\, B => 
        \I2.DTO_16_1l24r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834756_Rd1__net_1\, Y
         => \I2.DTO_1l24r\);
    
    \I2.STATE3l2r_1151\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_ns_il11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3L2R_413\);
    
    \I2.N_4667_1_adt_net_1046_\ : OAI21FTF
      port map(A => \I2.N_4261_303\, B => \I2.N_4283_I_0_40\, C
         => \I2.STATE2L2R_589\, Y => 
        \I2.N_4667_1_adt_net_1046__net_1\);
    
    \I5.SBYTE_70\ : MUX2H
      port map(A => \I5.SBYTEl5r_net_1\, B => \I5.N_24\, S => 
        \I5.N_406\, Y => \I5.SBYTE_70_net_1\);
    
    \I3.REG_1_ml73r\ : AND2
      port map(A => REGl73r, B => 
        \I3.REGMAPl9r_adt_net_854324__net_1\, Y => 
        \I3.VDBi_20l25r\);
    
    \I3.PIPEA1_308\ : MUX2L
      port map(A => \I3.PIPEA1l10r_net_1\, B => 
        \I3.PIPEA1_12l10r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__253\, Y => 
        \I3.PIPEA1_308_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I120_Y_0\ : AO21FTT
      port map(A => \I2.N537_i\, B => \I2.N531_adt_net_59960_\, C
         => \I2.N_140\, Y => \I2.N531\);
    
    FID_padl14r : OB33PH
      port map(PAD => FID(14), A => FID_cl14r);
    
    \I2.STATEe_1284\ : OR2
      port map(A => \I2.STATEe_ipl1r\, B => \I2.N_3450\, Y => 
        \I2.N_3453\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I14_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L12R_827\, B => 
        \I2.PIPE4_DTL14R_640\, Y => \I2.N_57_0\);
    
    TDCDRYB_pad : IB33
      port map(PAD => TDCDRYB, Y => TDCDRYB_c);
    
    DTE_padl26r : IOB33PH
      port map(PAD => DTE(26), A => \I2.DTE_1l26r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl26r);
    
    \I3.VDBoffa_31_iv_0l2r\ : AND2
      port map(A => \REGl207r\, B => 
        \I3.REGMAPl23r_adt_net_855016__net_1\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164214_\);
    
    \I2.DTE_21_1_IV_0L9R_1306\ : AND2
      port map(A => \I2.DTE_1l9r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1l9r_adt_net_38627_\);
    
    \I3.REGMAPl0r_1615\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un2_reg_ads_0_a2_0_a3_net_1\, Q => \I3.REGMAPL0R_722\);
    
    \I1.NCS0\ : DFFS
      port map(CLK => CLK_c, D => \I1.NCS0_56_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.NCS0_net_1\);
    
    \I3.VDBI_57_0_IV_0_0L8R_2221\ : AND3FFT
      port map(A => \I3.N_2014\, B => \I3.N_1917\, C => 
        \I3.REGl141r\, Y => \I3.VDBi_57l8r_adt_net_142723_\);
    
    \I2.PIPE1_DT_42_1_iv_1l25r\ : OAI21TTF
      port map(A => \I2.TDCDASl25r_net_1\, B => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        C => \I2.PIPE1_DT_42_1_iv_1_il25r_adt_net_46311_\, Y => 
        \I2.PIPE1_DT_42_1_iv_1_il25r\);
    
    \I1.REG_74_0_IV_0L191R_2043\ : AND2
      port map(A => \REGl191r\, B => \I1.N_65_92\, Y => 
        \I1.REG_74l191r_adt_net_131355_\);
    
    \I2.TRGCNTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGCNT_n2\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGCNTl2r_net_1\);
    
    \I2.STATE1_ns_i_i_a3l15r\ : AND2FT
      port map(A => \I2.N_3279_0_adt_net_855224__net_1\, B => 
        \I2.ERR_WORDS_RDY_net_1\, Y => \I2.N_154\);
    
    \I2.PIPE4_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl28r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl28r_net_1\);
    
    \I1.PAGECNT_n9_i_i\ : OAI21
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_854520__net_1\, 
        B => \I1.N_404_i_i_0_i\, C => \I1.N_473\, Y => 
        \I1.N_1380\);
    
    \I3.UN1_NRDMEBI_2_SQMUXA_3_2308\ : AND3FTT
      port map(A => \I3.STATE2l2r_net_1\, B => 
        \I3.NRDMEBi_0_sqmuxa_net_1\, C => 
        \I3.un1_NRDMEBi_2_sqmuxa_3_0_adt_net_153527_\, Y => 
        \I3.un1_NRDMEBi_2_sqmuxa_3_adt_net_153598_\);
    
    \I2.L2RF3\ : DFFS
      port map(CLK => CLK_c, D => \I2.L2RF2_i_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L2RF3_i\);
    
    \I1.REG_74_0_ivl329r\ : AO21
      port map(A => \REGl329r\, B => \I1.N_201\, C => 
        \I1.REG_74l329r_adt_net_118174_\, Y => \I1.REG_74l329r\);
    
    \I1.REG_74_0_iv_0l372r\ : AO21
      port map(A => \REGl372r\, B => \I1.N_660\, C => 
        \I1.REG_74l372r_adt_net_113310_\, Y => \I1.REG_74l372r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I71_Y\ : NAND2
      port map(A => \I2.N243_0\, B => \I2.N246_0\, Y => 
        \I2.N321_0\);
    
    \I2.DTOSl26r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl26r, Q => 
        \I2.DTOSl26r_net_1\);
    
    \I2.DTO_1l12r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l12r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l12r_Rd1__net_1\);
    
    \I3.VDBOFFB_30_IV_0L7R_2365\ : OR3
      port map(A => \I3.VDBoffb_30l7r_adt_net_161797_\, B => 
        \I3.VDBoffb_30l7r_adt_net_161793_\, C => 
        \I3.VDBoffb_30l7r_adt_net_161794_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161800_\);
    
    \I2.resyn_0_I2_TRGCNT_n4_0\ : XOR2
      port map(A => \I2.TRGCNTl4r_net_1\, B => 
        \I2.un9_tdctrgi_i_0\, Y => \I2.TRGCNT_n4_0\);
    
    \I3.VDBil28r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_368_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil28r_net_1\);
    
    \I1.REG_1_246\ : MUX2H
      port map(A => \REGl345r\, B => \I1.REG_74l345r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_246_net_1\);
    
    \I3.un224_reg_ads_0_a2_3_a2_0\ : NAND2
      port map(A => \I3.VASl5r_net_1\, B => \I3.VASl3r_net_1\, Y
         => \I3.N_558\);
    
    \I2.un2_evnt_word_I_13\ : XOR2
      port map(A => \I2.WOFFSETl3r_adt_net_854988__net_1\, B => 
        \I2.DWACT_FINC_E_0l0r\, Y => \I2.I_13_1\);
    
    \I3.REG3l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_130_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l5r_net_1\);
    
    \I2.DTO_1_880\ : MUX2L
      port map(A => \I2.DTO_1l6r_Rd1__net_1\, B => 
        \I2.DTO_16_1l6r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834776_Rd1__net_1\, Y
         => \I2.DTO_1l6r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I0_CO1_i_o2\ : NAND2
      port map(A => \I2.RAMDT4L7R_443\, B => \I2.PIPE4_DTL0R_411\, 
        Y => \I2.N_85_0\);
    
    \I2.SUB9_1_ADD_18x18_fast_I53_Y\ : NOR3FFT
      port map(A => \I2.N271\, B => \I2.N268\, C => \I2.N290\, Y
         => \I2.N321\);
    
    \I2.LEADSRAM.M0\ : RAM256x9SST
      generic map(MEMORYFILE => "LEAD_SRAM_M0.mem")

      port map(DO8 => \I2.LSRAM_OUTl8r\, DO7 => \I2.LSRAM_OUTl7r\, 
        DO6 => \I2.LSRAM_OUTl6r\, DO5 => \I2.LSRAM_OUTl5r\, DO4
         => \I2.LSRAM_OUTl4r\, DO3 => \I2.LSRAM_OUTl3r\, DO2 => 
        \I2.LSRAM_OUTl2r\, DO1 => \I2.LSRAM_OUTl1r\, DO0 => 
        \I2.LSRAM_OUTl0r\, WPE => OPEN, RPE => OPEN, DOS => OPEN, 
        WADDR7 => \GND\, WADDR6 => \GND\, WADDR5 => \GND\, WADDR4
         => \GND\, WADDR3 => \GND\, WADDR2 => 
        \I2.LSRAM_WADDRl2r_net_1\, WADDR1 => 
        \I2.LSRAM_WADDRl1r_net_1\, WADDR0 => 
        \I2.LSRAM_WADDRl0r_net_1\, RADDR7 => \GND\, RADDR6 => 
        \GND\, RADDR5 => \GND\, RADDR4 => \GND\, RADDR3 => \GND\, 
        RADDR2 => \I2.LSRAM_RADDRl2r_net_1\, RADDR1 => 
        \I2.LSRAM_RADDRl1r_net_1\, RADDR0 => 
        \I2.LSRAM_RADDRl0r_net_1\, DI8 => \I2.LSRAM_INl8r_net_1\, 
        DI7 => \I2.LSRAM_INl7r_net_1\, DI6 => 
        \I2.LSRAM_INl6r_net_1\, DI5 => \I2.LSRAM_INl5r_net_1\, 
        DI4 => \I2.LSRAM_INl4r_net_1\, DI3 => 
        \I2.LSRAM_INl3r_net_1\, DI2 => \I2.LSRAM_INl2r_net_1\, 
        DI1 => \I2.LSRAM_INl1r_net_1\, DI0 => 
        \I2.LSRAM_INl0r_net_1\, WRB => \I2.LSRAM_WR_net_1\, RDB
         => \I2.LSRAM_RD_net_1\, WBLKB => \GND\, RBLKB => \GND\, 
        PARODD => \GND\, WCLKS => CLK_c, RCLKS => CLK_c, DIS => 
        \GND\);
    
    \I2.DT_SRAM_0l10r\ : MUX2L
      port map(A => \I2.PIPE10_DTl10r_net_1\, B => 
        \I2.PIPE5_DTl10r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854224__net_1\, Y => 
        \I2.N_878\);
    
    \I2.ADEl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl7r);
    
    GA_padl2r : IB33
      port map(PAD => GA(2), Y => GA_cl2r);
    
    REGl289r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_190_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl289r\);
    
    \I3.VDBOFFA_31_IV_0L3R_2572\ : AO21
      port map(A => \REGl192r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.VDBoffa_31l3r_adt_net_164028_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164069_\);
    
    \I2.PIPE1_DT_42_1_IVL6R_1485\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        B => \I2.PIPE1_DT_12l6r_net_1\, Y => 
        \I2.PIPE1_DT_42l6r_adt_net_50924_\);
    
    \I2.L2TYPE_4_il9r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855716__net_1\, B => 
        \I2.N_4443_adt_net_67572_\, C => 
        \I2.N_4443_adt_net_67615_\, Y => \I2.N_4443\);
    
    \I3.REG_1_209\ : MUX2L
      port map(A => VDB_inl28r, B => \I3.REGl161r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\, Y => 
        \I3.REG_1_209_0\);
    
    \I2.BITCNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.BITCNT_939\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.BITCNTl1r_net_1\);
    
    \I3.TICKil0r_1449\ : DFFC
      port map(CLK => CLK_c, D => \I3.un6_tcnt1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TICKL0R_556);
    
    \I1.REG_74_0_IVL293R_1925\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l293r_adt_net_121470_\);
    
    \I1.N_193_adt_net_118660_\ : NAND3FFT
      port map(A => \I1.N_41_9_adt_net_3739__net_1\, B => 
        \I1.N_193_adt_net_118653__net_1\, C => \I1.N_273_9\, Y
         => \I1.N_193_adt_net_118660__net_1\);
    
    \I1.REG_74_0_IV_0_0L249R_1977\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l249r_adt_net_125863_\);
    
    SP0_pad : OB33PH
      port map(PAD => SP0, A => \GND\);
    
    VAD_padl20r : OTB33PH
      port map(PAD => VAD(20), A => \I3.VADml20r\, EN => 
        NOEAD_c_i_0);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I32_P0N_1759\ : OR2FT
      port map(A => \I2.LSRAM_OUTl11r\, B => 
        \I2.PIPE7_DTL11R_694\, Y => \I2.N264_0_866\);
    
    \I3.VDBI_31L1R_2717\ : AO21
      port map(A => \I3.VDBi_31l1r_adt_net_506111_\, B => 
        \I3.VDBi_31l1r_adt_net_506164_\, C => 
        \I3.VDBi_31l1r_adt_net_614331_\, Y => 
        \I3.VDBi_31l1r_net_1\);
    
    \I2.un1_tdc_res_47_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl407r, Y => 
        \I2.N_4628_i_0\);
    
    \I2.resyn_0_I2_FID_434\ : MUX2H
      port map(A => FID_cl18r, B => \I2.FID_7l18r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\, 
        Y => \I2.FID_434\);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854676_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854676__net_1\);
    
    \I2.FID_7_0_IVL7R_1719\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl55r, C => 
        \I2.FID_7l7r_adt_net_92833_\, Y => 
        \I2.FID_7l7r_adt_net_92841_\);
    
    \I1.REG_74_0_IV_0_0L247R_1979\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l247r_adt_net_126035_\);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854248_\ : BFR
      port map(A => \I2.WR_SRAM_2_adt_net_748__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854248__net_1\);
    
    \I3.REG_1_273\ : MUX2H
      port map(A => VDB_inl1r, B => \I3.REGl92r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_273_0\);
    
    \I2.G_EVNT_NUM_n5_i_0\ : NOR3
      port map(A => EV_RES_C_569, B => \I2.N_319\, C => 
        \I2.N_4672\, Y => \I2.N_4345\);
    
    \I2.DTO_16_1_iv_0l20r\ : OR2
      port map(A => \I2.DTO_16_1l20r_adt_net_30793_\, B => 
        \I2.DTO_16_1l20r_adt_net_30794_\, Y => \I2.DTO_16_1l20r\);
    
    \I2.PIPE1_DT_42_1_IVL10R_1463\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl42r_net_1\, C => 
        \I2.PIPE1_DT_42l10r_adt_net_49932_\, Y => 
        \I2.PIPE1_DT_42l10r_adt_net_49950_\);
    
    \I3.PULSE_46_0_iv_0_0l9r\ : AO21
      port map(A => PULSEl9r, B => 
        \I3.N_311_adt_net_854748__net_1\, C => 
        \I3.PULSE_46l9r_adt_net_146747_\, Y => \I3.PULSE_46l9r\);
    
    \I2.REG_1l45r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n13_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl45r);
    
    \I2.un1_STATE2_15_i_0_a2_1_i\ : NAND2
      port map(A => \I2.STATE2l5r_net_1\, B => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__57\, Y => 
        \I2.N_4641\);
    
    \I1.REG_74_0_IV_0_0L250R_1976\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l250r_adt_net_125777_\);
    
    \I2.PIPE1_DT_42_1_IVL4R_1498\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl0r\, Y => 
        \I2.PIPE1_DT_42l4r_adt_net_51424_\);
    
    \I1.REG_74_0_IVL295R_1923\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l295r_adt_net_121298_\);
    
    \I3.VDBOFFB_30_IV_0L2R_2450\ : AO21
      port map(A => \REGl327r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l2r_adt_net_162714_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162743_\);
    
    \I3.VDBi_40l12r\ : MUX2L
      port map(A => \I3.N_350\, B => \I3.N_1857\, S => 
        \I3.N_354_0_adt_net_855368__net_1\, Y => 
        \I3.VDBi_40l12r_net_1\);
    
    \I2.PIPE8_DT_559\ : MUX2L
      port map(A => \I2.PIPE8_DTl31r_net_1\, B => \I2.N_4418\, S
         => \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_559_net_1\);
    
    \I2.L2SERV_n2\ : XOR2
      port map(A => \I2.RPAGEl14r\, B => \I2.L2SERV_c1_net_1\, Y
         => \I2.L2SERV_n2_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I9_P0N_i_o3\ : OR2
      port map(A => \I2.RAMDT4L12R_144\, B => 
        \I2.PIPE4_DTL9R_471\, Y => \I2.N_13_1\);
    
    \I2.OFFSET_37_24l5r\ : MUX2L
      port map(A => \I2.N_816\, B => \I2.N_808\, S => 
        \I2.PIPE7_DTL26R_357\, Y => \I2.N_824\);
    
    \I2.EVNT_NUM_n11\ : XOR2
      port map(A => \I2.N_1232\, B => \I2.N_1233\, Y => 
        \I2.EVNT_NUM_n11_net_1\);
    
    \I2.OFFSET_37_19l0r\ : MUX2L
      port map(A => \REGl277r\, B => \REGl213r\, S => 
        \I2.PIPE7_DTl27r_net_1\, Y => \I2.N_779\);
    
    \I5.REG_2_sqmuxa_0_adt_net_975_\ : NAND2
      port map(A => \I5.AIR_CHAIN_net_1\, B => 
        \I5.sstate2_5_sqmuxa\, Y => 
        \I5.REG_2_sqmuxa_0_adt_net_975__net_1\);
    
    \I2.N_4529_adt_net_1136_\ : AO21
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_215\, C
         => LEAD_FLAGl6r, Y => \I2.N_4529_adt_net_1136__net_1\);
    
    \I3.PIPEA1_302\ : MUX2L
      port map(A => \I3.PIPEA1l4r_net_1\, B => 
        \I3.PIPEA1_12l4r_net_1\, S => 
        \I3.un1_STATE2_15_1_adt_net_1342__net_1\, Y => 
        \I3.PIPEA1_302_net_1\);
    
    \I2.DTO_16_1_IV_0_0L6R_1192\ : AO21
      port map(A => \I2.N_457\, B => \I2.DTE_2_1l6r_net_1\, C => 
        \I2.DTO_16_1l6r_adt_net_33910_\, Y => 
        \I2.DTO_16_1l6r_adt_net_33921_\);
    
    REGl381r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_282_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl381r\);
    
    \I3.PIPEB_106\ : AO21
      port map(A => DPR_cl27r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\, 
        C => \I3.PIPEB_106_adt_net_159579_\, Y => 
        \I3.PIPEB_106_net_1\);
    
    \I2.STATE3l3r_1153\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3L3R_415\);
    
    \I3.un121_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_639\, B => \I3.N_553\, Y => 
        \I3.un121_reg_ads_0_a2_0_a3_net_1\);
    
    \I1.SBYTE_8_0_i_a2l3r\ : OR2
      port map(A => \I1.sstatel2r_net_1\, B => 
        \I1.sstatel9r_net_1\, Y => \I1.N_602_i\);
    
    \I3.VDBil24r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_364_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil24r_net_1\);
    
    \I3.VAS_74\ : MUX2L
      port map(A => VAD_inl12r, B => \I3.VASl12r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_74_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I121_Y_i_a3_0\ : AO21
      port map(A => \I2.RAMDT4L5R_819\, B => 
        \I2.PIPE4_DTl5r_adt_net_854412__net_1\, C => 
        \I2.N_107_adt_net_276024_\, Y => 
        \I2.ADD_21x21_fast_I121_Y_i_a3_0_i\);
    
    \I3.STATE1_0l8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl2r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl8r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I185_Y\ : XOR2
      port map(A => \I2.N507\, B => \I2.ADD_21x21_fast_I185_Y_0\, 
        Y => \I2.un27_pipe5_dt0l15r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I147_Y_0\ : XOR2FT
      port map(A => \I2.SUB8l11r_adt_net_855580__net_1\, B => 
        \I2.N_3547_i_i\, Y => \I2.ADD_18x18_fast_I147_Y_0\);
    
    \I2.OFFSET_37_16l1r\ : MUX2L
      port map(A => \REGl262r\, B => \REGl198r\, S => 
        \I2.PIPE7_DTL27R_84\, Y => \I2.N_756\);
    
    \I2.STATE1_ns_i_o2l15r\ : AND2
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\, 
        B => \I2.STATE1l9r_net_1\, Y => \I2.N_3280\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I101_Y\ : AOI21
      port map(A => \I2.N313_1\, B => \I2.N316_i_i\, C => 
        \I2.N312_0\, Y => \I2.N355_0\);
    
    \I1.REG_1_162\ : MUX2H
      port map(A => \REGl261r\, B => \I1.REG_74l261r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855452__net_1\, Y => 
        \I1.REG_1_162_net_1\);
    
    FBOUTl4r : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_62_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \FBOUTl4r\);
    
    \I2.L2SERVl2r_1508\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_920_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL14R_615\);
    
    \I2.DTE_1l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_840_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l0r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I138_Y_0_a2\ : AND3FTT
      port map(A => \I2.N_74_i_0_i\, B => \I2.N_52\, C => 
        \I2.N_100_adt_net_58424_\, Y => \I2.N_100\);
    
    \I2.TOKOUT_FL_674_1590\ : AND3FFT
      port map(A => \I2.PIPE1_DT_1_sqmuxa\, B => \I2.N_3890\, C
         => \I2.TOKOUT_FL_674_adt_net_1115__net_1\, Y => 
        \I2.TOKOUT_FL_674_adt_net_61319_\);
    
    \I3.VDBI_20_IVL14R_2189\ : NOR2FT
      port map(A => REGl46r, B => \I3.N_2033\, Y => 
        \I3.VDBi_20l14r_adt_net_140054_\);
    
    \I1.REG_1_248\ : MUX2H
      port map(A => \REGl347r\, B => \I1.REG_74l347r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_248_net_1\);
    
    \I2.DTESl0r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl0r, Q => 
        \I2.DTESl0r_net_1\);
    
    \I2.PIPE6_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_467_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl13r_net_1\);
    
    \I2.PIPE5_DT_690\ : MUX2L
      port map(A => \I2.PIPE5_DTl14r_net_1\, B => 
        \I2.PIPE5_DT_6l14r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_690_net_1\);
    
    \I2.STATE1_ns_a3_1l7r\ : OR2
      port map(A => \I2.END_TDC1_0_sqmuxa_1_net_1\, B => 
        \I2.NWPIPE1_4_sqmuxa_1_0\, Y => \I2.STATE1_ns_1l7r\);
    
    \I2.STATE3_0_sqmuxa_0_a7_1\ : AND3
      port map(A => \I2.DTES_i_0_il30r\, B => \I2.DTESl28r_net_1\, 
        C => \I2.STATE3_0_sqmuxa_1_0_adt_net_24559_\, Y => 
        \I2.STATE3_0_sqmuxa_1_0\);
    
    \I2.DTOSl6r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl6r, Q => 
        \I2.DTOSl6r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I154_Y\ : XOR2FT
      port map(A => \I2.N442_i\, B => 
        \I2.ADD_18x18_fast_I154_Y_0\, Y => \I2.SUB9_1l17r\);
    
    \I2.DTOSl19r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl19r, Q => 
        \I2.DTOSl19r_net_1\);
    
    RAMAD_padl16r : OB33PH
      port map(PAD => RAMAD(16), A => RAMAD_cl16r);
    
    \I2.PIPE1_DT_42_1_IVL19R_1399\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\, B => 
        \I2.PIPE1_DT_30l19r_net_1\, C => 
        \I2.PIPE1_DT_42l19r_adt_net_47247_\, Y => 
        \I2.PIPE1_DT_42l19r_adt_net_47262_\);
    
    \I3.VDBOFFB_30_IV_0L6R_2380\ : AO21
      port map(A => \REGl395r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l6r_adt_net_161978_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161985_\);
    
    \I2.DTE_21_1l4r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l4r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l4r_Rd1__net_1\);
    
    \I5.DATA_12l14r\ : MUX2L
      port map(A => REGl131r, B => \I5.SBYTEl6r_net_1\, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l14r_net_1\);
    
    \I2.BNCID_VECTra15_1\ : AND2
      port map(A => \I2.TRGSERVL0R_465\, B => \I2.TRGSERVL1R_468\, 
        Y => \I2.BNCID_VECTra15_1_net_1\);
    
    \I2.PIPE6_DT_469\ : MUX2H
      port map(A => \I2.PIPE5_DTl15r_net_1\, B => 
        \I2.PIPE6_DTl15r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_469_net_1\);
    
    \I2.PIPE3_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl1r_net_1\);
    
    \I2.ROFFSET_c9\ : AND2
      port map(A => \I2.ROFFSETl9r_net_1\, B => 
        \I2.ROFFSET_c8_net_1\, Y => \I2.ROFFSET_c9_net_1\);
    
    \I5.SDAnoe_8_0\ : AO21
      port map(A => \I5.N_70\, B => \I5.SDAnoe_8_adt_net_9739_\, 
        C => \I5.SDAnoe_8_adt_net_991__net_1\, Y => \I5.SDAnoe_8\);
    
    \I3.VAS_66\ : MUX2L
      port map(A => VAD_inl4r, B => \I3.VASl4r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_66_net_1\);
    
    \I3.VDBoffb_53\ : OR3
      port map(A => \I3.VDBoffb_53_adt_net_162980_\, B => 
        \I3.VDBoffb_30l1r_adt_net_162939_\, C => 
        \I3.VDBoffb_30l1r_adt_net_162940_\, Y => 
        \I3.VDBoffb_53_net_1\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854460_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854472__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854460__net_1\);
    
    \I3.N_1910_0_adt_net_854336_\ : BFR
      port map(A => \I3.N_1910_0\, Y => 
        \I3.N_1910_0_adt_net_854336__net_1\);
    
    \I3.VDBOFFA_31_IV_0L7R_2505\ : AO21
      port map(A => \REGl172r\, B => \I3.REGMAPl18r_net_1\, C => 
        \I3.VDBoffa_31l7r_adt_net_163288_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163314_\);
    
    \I2.OFFSET_37_10l2r\ : MUX2L
      port map(A => \I2.N_701\, B => \I2.N_693\, S => 
        \I2.PIPE7_DTL26R_354\, Y => \I2.N_709\);
    
    \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__2753\ : OAI21TTF
      port map(A => \I2.N_176_i_adt_net_855708__net_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, C => 
        \I2.N_4667_1_ADT_NET_1046__33\, Y => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\);
    
    \I3.VDBOFFA_31_IV_0L0R_2622\ : AND2
      port map(A => \REGl253r\, B => \I3.REGMAPl29r_net_1\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164610_\);
    
    \I2.L2TYPEl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_597_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl8r_net_1\);
    
    \I2.PIPE7_DTL27R_2777\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_70\);
    
    REGl398r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_299_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl398r\);
    
    \I2.RAMADl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l8r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl8r);
    
    \I3.VDBOFFA_31_IV_0L4R_2551\ : AND2
      port map(A => \REGl281r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        Y => \I3.VDBoffa_31l4r_adt_net_163854_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I211_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl15r\, B => 
        \I2.PIPE7_DTl15r_net_1\, Y => 
        \I2.SUB_21x21_fast_I211_Y_0\);
    
    \I2.PIPE1_DT_729\ : MUX2L
      port map(A => \I2.PIPE1_DTl2r_net_1\, B => 
        \I2.PIPE1_DT_42l2r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854588__net_1\, 
        Y => \I2.PIPE1_DT_729_net_1\);
    
    \I3.VDBi_363\ : MUX2L
      port map(A => \I3.VDBil23r_net_1\, B => \I3.VDBi_57l23r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_363_net_1\);
    
    \I3.VDBoffl5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_121_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl5r_net_1\);
    
    \I2.MIC_ERR_REGSl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_342_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl13r_net_1\);
    
    REGl380r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_281_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl380r\);
    
    \I3.un47_reg_ads_0_a2_0_a2_993\ : OR2FT
      port map(A => \I3.WRITES_8\, B => \I3.N_546_374\, Y => 
        \I3.N_547_371\);
    
    \I2.RAMDT4l0r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl0r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l0r_net_1\);
    
    \I2.N_3877_adt_net_855268_\ : BFR
      port map(A => \I2.N_3877\, Y => 
        \I2.N_3877_adt_net_855268__net_1\);
    
    \I2.L2TYPEl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_589_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl0r_net_1\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l4r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl4r_net_1\, Q => 
        \I2.DIN_REG1l4r\);
    
    \I2.RESYN_0_I2_LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_949\ : OR3FFT
      port map(A => \I2.PIPE4_DTl31r_net_1\, B => 
        \I2.NWPIPE5_net_1\, C => \I2.NWPIPE4_575\, Y => 
        \I2.N_4524_adt_net_16803_\);
    
    \I3.UN2_VSEL_1_I_0_A2_2102\ : OR3
      port map(A => AMB_c_i_0_il5r, B => AMB_cl4r, C => 
        \I3.N_2055_adt_net_134991_\, Y => 
        \I3.N_2055_adt_net_134992_\);
    
    \I3.REGMAPl3r_1631\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un17_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL3R_738\);
    
    \I2.MIC_ERR_REGSl46r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_375_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl46r_net_1\);
    
    \I2.DTO_9_iv_0l23r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl23r_net_1\, 
        C => \I2.DTO_9l23r_adt_net_30048_\, Y => \I2.DTO_9l23r\);
    
    \I3.VDBoff_116\ : MUX2L
      port map(A => \I3.VDBoffl0r_net_1\, B => \I3.N_2064\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_116_net_1\);
    
    \I2.MIC_REG2_312\ : MUX2H
      port map(A => \I2.MIC_REG2l3r_adt_net_834020_Rd1__net_1\, B
         => \I2.MIC_REG2_i_0_il4r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_net_1\, Y => 
        \I2.MIC_REG2_312_net_1\);
    
    \I3.PIPEAl21r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_252_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl21r_net_1\);
    
    \I2.ROFFSET_n3\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855700__net_1\, B => 
        \I2.ROFFSET_n3_tz_i\, Y => \I2.ROFFSET_n3_net_1\);
    
    \I2.un1_tdc_res_27_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl415r, Y => 
        \I2.N_4608_i_0\);
    
    \I2.DT_TEMP_780\ : MUX2H
      port map(A => \I2.DT_TEMPl19r_net_1\, B => 
        \I2.DT_TEMP_7l19r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_780_net_1\);
    
    \I2.PIPE9_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_289_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl20r_net_1\);
    
    \I3.STATE1_0l9r_1610\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL9R_717\);
    
    \I2.MIC_REG2_315\ : MUX2L
      port map(A => \I2.MIC_REG2l7r_net_1\, B => 
        \I2.MIC_REG2l6r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG2_315_net_1\);
    
    TOKINA_pad : OB33PH
      port map(PAD => TOKINA, A => TOKINA_c);
    
    REGl193r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_94_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl193r\);
    
    \I5.REG_1_41\ : MUX2L
      port map(A => \I5.SENS_ADDRl0r_net_1\, B => REGl428r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_41_net_1\);
    
    \I5.COMMAND_14\ : MUX2H
      port map(A => \I5.COMMANDl2r_net_1\, B => 
        \I5.COMMAND_4l2r_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.COMMAND_14_net_1\);
    
    \I3.VDBi_23l1r_adt_net_145532_\ : NOR3
      port map(A => GA_cl1r, B => \I3.N_1907_266\, C => 
        \I3.N_2042\, Y => \I3.VDBi_23l1r_adt_net_145532__net_1\);
    
    VDB_padl21r : IOB33PH
      port map(PAD => VDB(21), A => \I3.VDBml21r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl21r);
    
    \I2.ROFFSETl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_909_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl9r_net_1\);
    
    \I3.REGMAPL39R_2800\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un176_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL39R_112\);
    
    \I2.CRC32l15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_810_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l15r_net_1\);
    
    \I3.REG_1_282\ : MUX2L
      port map(A => VDB_inl0r, B => REGl101r, S => 
        \I3.N_318_adt_net_855888__net_1\, Y => \I3.REG_1_282_0\);
    
    \I3.VDBOFFA_31_IV_0L7R_2496\ : AND2
      port map(A => \REGl252r\, B => \I3.REGMAPl28r_net_1\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163280_\);
    
    \I1.N_347_adt_net_854792_\ : BFR
      port map(A => \I1.N_347\, Y => 
        \I1.N_347_adt_net_854792__net_1\);
    
    \I2.DT_SRAM_0l11r\ : MUX2L
      port map(A => \I2.PIPE10_DTl11r_net_1\, B => 
        \I2.PIPE5_DTl11r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, Y => 
        \I2.N_879\);
    
    \I1.REG_74_0_IV_0L221R_2006\ : AND2
      port map(A => \REGl221r\, B => \I1.N_97\, Y => 
        \I1.REG_74l221r_adt_net_128566_\);
    
    \I1.REG_16_sqmuxa_adt_net_855456_\ : BFR
      port map(A => \I1.REG_16_sqmuxa\, Y => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\);
    
    \I2.PIPE5_DT_6_0l16r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l16r\, B => 
        \I2.un27_pipe5_dt0l16r\, S => 
        \I2.dataout_0_adt_net_855804__net_1\, Y => \I2.N_1085\);
    
    \I2.DTE_21_1_IV_2L1R_1342\ : OAI21TTF
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855208__net_1\, 
        B => \I2.DT_TEMPl1r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39583_\, Y => 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39592_\);
    
    \I1.REG_74_0_IV_I_A2L210R_2024\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, Y => 
        \I1.N_1349_adt_net_129673_\);
    
    \I3.TICKi_0l0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.un6_tcnt1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TICKL0R_2);
    
    \I2.PIPE8_DT_16_0l19r\ : MUX2H
      port map(A => \I2.PIPE8_DTl19r_net_1\, B => 
        \I2.PIPE7_DTl19r_net_1\, S => 
        \I2.N_565_0_adt_net_855736__net_1\, Y => \I2.N_585\);
    
    \I2.PIPE4_DTl11r_1147_1734\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL11R_841\);
    
    \I2.DTE_21_1_IV_0L6R_1321\ : AND2
      port map(A => \I2.DT_SRAMl6r_net_1\, B => 
        \I2.N_199_0_ADT_NET_1054__36\, Y => 
        \I2.DTE_21_1l6r_adt_net_38971_\);
    
    REGl327r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_228_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl327r\);
    
    \I3.VDBOFFB_30_IV_0L4R_2416\ : AO21
      port map(A => \REGl393r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l4r_adt_net_162358_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162365_\);
    
    \I3.REG_1l82r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_263_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl82r);
    
    \I3.PULSE_46_0_iv_0_0l5r\ : AO21
      port map(A => PULSEL5R_16, B => 
        \I3.N_311_adt_net_854752__net_1\, C => 
        \I3.PULSE_46l5r_adt_net_147097_\, Y => \I3.PULSE_46l5r\);
    
    \I3.VDBOFFB_30_IV_0L4R_2404\ : AND2
      port map(A => \REGl377r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162322_\);
    
    \I2.un13_start_giro_i_i_a2\ : NAND2
      port map(A => \I2.START_GIRO_net_1\, B => \I2.N_3850\, Y
         => \I2.N_128_1\);
    
    \I5.REG_1l447r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_30_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl447r);
    
    \I1.sstatel6r_1607\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl4r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL6R_714\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l2r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl2r_net_1\, Q => 
        \I2.DIN_REG1_0l2r\);
    
    TDCDA_padl6r : IB33
      port map(PAD => TDCDA(6), Y => TDCDA_cl6r);
    
    \I2.DTESl5r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl5r, Q => 
        \I2.DTESl5r_net_1\);
    
    \I3.PIPEAl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_232_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl1r_net_1\);
    
    \I1.REG_1_104\ : MUX2H
      port map(A => \REGl203r\, B => \I1.N_1342\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_104_net_1\);
    
    \I3.PIPEBl26r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_105_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl26r_net_1\);
    
    \I2.TDCDBSl8r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl8r, Q => 
        \I2.TDCDBSl8r_net_1\);
    
    \I2.RAMDT4L12R_2813\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_141\);
    
    \I2.PIPE5_DT_6_dl17r\ : MUX2L
      port map(A => \I2.PIPE4_DTl17r_net_1\, B => 
        \I2.un27_pipe5_dt1l17r\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855616__net_1\, Y => 
        \I2.PIPE5_DT_6_dl17r_net_1\);
    
    \I2.EVNT_NUMlde_i_a2\ : NOR2
      port map(A => EV_RES_c, B => \I2.STATE1l17r_net_1\, Y => 
        \I2.N_3770\);
    
    \I2.PIPE7_DTl13r_1585\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl13r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL13R_692\);
    
    \I1.REG_74_2_4L228R_1852\ : XOR2
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__761\, B
         => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854396__net_1\, 
        Y => \I1.REG_74_2_4_il228r_adt_net_115255_\);
    
    \I3.PIPEA_8l18r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854468__net_1\, B => 
        \I3.N_227\, Y => \I3.PIPEA_8l18r_net_1\);
    
    \I2.SUB9l18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_586_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l18r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I153_Y_I_O4_1565\ : AO21
      port map(A => \I2.PIPE4_DTL17R_636\, B => 
        \I2.PIPE4_DTl13r_net_1\, C => \I2.RAMDT4L12R_793\, Y => 
        \I2.N_33_0_adt_net_55957_\);
    
    \I3.REG_44_il90r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_1636_adt_net_150083_\, Y => \I3.N_1636\);
    
    \I1.ISCK_53\ : MUX2L
      port map(A => \F_SCK_c\, B => \I1.sstate_nsl9r\, S => 
        \I1.ISCK_0_sqmuxa\, Y => \I1.ISCK_53_net_1\);
    
    \I3.un7_noe32ri_0_i_a3\ : OA21FTT
      port map(A => \I3.N_290\, B => \I3.LWORDS_net_1\, C => 
        NOEAD_c, Y => NOE32R_c);
    
    \I2.OFFSET_37_18l3r\ : MUX2L
      port map(A => \REGl248r\, B => \REGl184r\, S => 
        \I2.PIPE7_DTL27R_82\, Y => \I2.N_774\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I3_P0N_i_o3\ : OR2
      port map(A => \I2.RAMDT4L3R_765\, B => 
        \I2.PIPE4_DTl3r_adt_net_854548__net_1\, Y => \I2.N_28\);
    
    \I5.REG_1l428r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_41_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl428r);
    
    \I2.PIPE8_DT_21l16r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl16r\, B => 
        \I2.PIPE8_DT_16l16r_net_1\, S => \I2.NWPIPE7_net_1\, Y
         => \I2.PIPE8_DT_21l16r_net_1\);
    
    \I2.I_1339_ca_0_and2\ : AND2FT
      port map(A => \I2.OFFSETL4R_675\, B => \I2.SUB8L7R_704\, Y
         => \I2.N_3541_i_i\);
    
    \I2.PIPE1_DT_42_1_IVL16R_1413\ : OAI21FTF
      port map(A => REGl420r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855816__net_1\, C => 
        \I2.PIPE1_DT_42l16r_adt_net_47833_\, Y => 
        \I2.PIPE1_DT_42l16r_adt_net_47850_\);
    
    \I2.DTE_1_850\ : MUX2L
      port map(A => \I2.DTE_1l10r_Rd1__net_1\, B => 
        \I2.DTE_21_1l10r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, Y => 
        \I2.DTE_1l10r\);
    
    \I2.DTE_21_1_IV_0_0L22R_1254\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l22r\, C
         => \I2.DTE_21_1l22r_adt_net_37394_\, Y => 
        \I2.DTE_21_1l22r_adt_net_37395_\);
    
    \I2.DT_TEMP_791\ : MUX2H
      port map(A => \I2.DT_TEMPl30r_net_1\, B => 
        \I2.DT_TEMP_7l30r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_791_net_1\);
    
    \I2.BNCID_VECT_tile_0_WADDR_REG1l3r\ : DFF
      port map(CLK => CLK_c, D => \I2.TRGARRl3r_net_1\, Q => 
        \I2.WADDR_REG1l3r\);
    
    \I2.DTO_16_1_IV_0L13R_1154\ : AO21
      port map(A => \I2.N_457\, B => \I2.N_44_i_0\, C => 
        \I2.DTO_16_1l13r_adt_net_32384_\, Y => 
        \I2.DTO_16_1l13r_adt_net_32395_\);
    
    REGl219r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_120_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl219r\);
    
    \I2.un1_STATE1_40_1_adt_net_812_\ : OR3
      port map(A => \I2.N_3798\, B => 
        \I2.un1_STATE1_40_1_adt_net_45409__net_1\, C => 
        \I2.un1_STATE1_40_1_adt_net_45413__net_1\, Y => 
        \I2.un1_STATE1_40_1_adt_net_812__net_1\);
    
    \I2.STATE3_NSL12R_1045\ : AND2
      port map(A => \I2.STATE3L3R_416\, B => 
        \I2.STOP_RDSRAM_net_1\, Y => 
        \I2.STATE3_nsl12r_adt_net_24672_\);
    
    \I2.ADO_3l10r\ : MUX2L
      port map(A => \I2.WOFFSETl11r\, B => \I2.ROFFSETl11r_net_1\, 
        S => NOESRAME_C_243, Y => \I2.ADO_3l10r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L3R_2568\ : AND2
      port map(A => \REGl248r\, B => \I3.REGMAPl28r_net_1\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164040_\);
    
    \I3.PIPEBl23r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_102_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl23r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I61_Y\ : NAND2
      port map(A => \I2.N294\, B => \I2.N298\, Y => \I2.N329\);
    
    \I1.REG_74l188r_891\ : OR2
      port map(A => \I1.REG_4_sqmuxa\, B => 
        \I1.N_65_ADT_NET_1433__217\, Y => \I1.N_57_269\);
    
    \I2.LEADSRAM.M1\ : RAM256x9SST
      generic map(MEMORYFILE => "LEAD_SRAM_M1.mem")

      port map(DO8 => \I2.LSRAM_OUTl17r\, DO7 => 
        \I2.LSRAM_OUTl16r\, DO6 => \I2.LSRAM_OUTl15r\, DO5 => 
        \I2.LSRAM_OUTl14r\, DO4 => \I2.LSRAM_OUTl13r\, DO3 => 
        \I2.LSRAM_OUTl12r\, DO2 => \I2.LSRAM_OUTl11r\, DO1 => 
        \I2.LSRAM_OUTl10r\, DO0 => \I2.LSRAM_OUTl9r\, WPE => OPEN, 
        RPE => OPEN, DOS => OPEN, WADDR7 => \GND\, WADDR6 => 
        \GND\, WADDR5 => \GND\, WADDR4 => \GND\, WADDR3 => \GND\, 
        WADDR2 => \I2.LSRAM_WADDRl2r_net_1\, WADDR1 => 
        \I2.LSRAM_WADDRl1r_net_1\, WADDR0 => 
        \I2.LSRAM_WADDRl0r_net_1\, RADDR7 => \GND\, RADDR6 => 
        \GND\, RADDR5 => \GND\, RADDR4 => \GND\, RADDR3 => \GND\, 
        RADDR2 => \I2.LSRAM_RADDRl2r_net_1\, RADDR1 => 
        \I2.LSRAM_RADDRl1r_net_1\, RADDR0 => 
        \I2.LSRAM_RADDRl0r_net_1\, DI8 => \I2.LSRAM_INl17r_net_1\, 
        DI7 => \I2.LSRAM_INl16r_net_1\, DI6 => 
        \I2.LSRAM_INl15r_net_1\, DI5 => \I2.LSRAM_INl14r_net_1\, 
        DI4 => \I2.LSRAM_INl13r_net_1\, DI3 => 
        \I2.LSRAM_INl12r_net_1\, DI2 => \I2.LSRAM_INl11r_net_1\, 
        DI1 => \I2.LSRAM_INl10r_net_1\, DI0 => 
        \I2.LSRAM_INl9r_net_1\, WRB => \I2.LSRAM_WR_net_1\, RDB
         => \I2.LSRAM_RD_net_1\, WBLKB => \GND\, RBLKB => \GND\, 
        PARODD => \GND\, WCLKS => CLK_c, RCLKS => CLK_c, DIS => 
        \GND\);
    
    \I5.REG_1l434r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_17_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl434r);
    
    \I3.REG2_144\ : MUX2L
      port map(A => VDB_inl3r, B => \I3.REG2l3r_net_1\, S => 
        \I3.REG3_0_sqmuxa\, Y => \I3.REG2_144_net_1\);
    
    \I2.REG_1_n4_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855784__net_1\, B
         => REGl36r, Y => \I2.REG_1_n4_0_net_1\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2198\ : AO21
      port map(A => REGl45r, B => \I3.N_403_1\, C => 
        \I3.VDBi_57l13r_adt_net_140582_\, Y => 
        \I3.VDBi_57l13r_adt_net_140593_\);
    
    \I3.VDBm_0l15r\ : MUX2L
      port map(A => \I3.PIPEAl15r_net_1\, B => 
        \I3.PIPEBl15r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_157\);
    
    \I2.TRGARRl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGARR_3l3r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGARRl3r_net_1\);
    
    \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092_\ : BFR
      port map(A => \I2.un3_tdcgda1_1_adt_net_821__net_1\, Y => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092__net_1\);
    
    \I2.PIPE1_DT_42_1_IVL10R_1462\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl6r\, Y => 
        \I2.PIPE1_DT_42l10r_adt_net_49942_\);
    
    \I2.OFFSET_37_29l0r\ : MUX2L
      port map(A => \I2.N_851\, B => \I2.N_739\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l0r\);
    
    \I2.PIPE5_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_677_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl1r_net_1\);
    
    \I3.N_1905_1_adt_net_855376_\ : BFR
      port map(A => \I3.N_1905_1\, Y => 
        \I3.N_1905_1_adt_net_855376__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I40_Y\ : AND2
      port map(A => \I2.G_1_0\, B => \I2.N305_adt_net_70150_\, Y
         => \I2.N305\);
    
    \I1.REG_1_217\ : MUX2H
      port map(A => \REGl316r\, B => \I1.REG_74l316r_net_1\, S
         => \I1.N_50_0_ADT_NET_1409__295\, Y => 
        \I1.REG_1_217_net_1\);
    
    \I2.SUB8l3r_1603\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_506_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8L3R_710\);
    
    \I2.WOFFSET_13_0l0r\ : OAI21TTF
      port map(A => 
        \I2.WOFFSETl0r_adt_net_854636__adt_net_855712__net_1\, B
         => \I2.N_2864_0_adt_net_854264__net_1\, C => 
        \I2.WPAGEe_adt_net_855060__net_1\, Y => 
        \I2.WOFFSET_13l0r\);
    
    \I2.resyn_0_I2_FID_426\ : MUX2H
      port map(A => FID_cl10r, B => \I2.FID_7l10r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\, 
        Y => \I2.FID_426\);
    
    \I2.DTE_1l28r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l28r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l28r_Rd1__net_1\);
    
    \I2.PHASE_863\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_C_241);
    
    \I2.DT_SRAM_IL27R_1077\ : NOR2FT
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__27\, B => 
        \I2.DT_SRAM_0_il27r_net_1\, Y => 
        \I2.N_4647_adt_net_29104_\);
    
    \I5.REG_1l436r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_19_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl436r);
    
    \I2.PIPE1_DT_42_1_IVL0R_1523\ : OAI21TTF
      port map(A => GA_cl0r, B => \I2.N_3238\, C => 
        \I2.PIPE1_DT_42l0r_adt_net_52246_\, Y => 
        \I2.PIPE1_DT_42l0r_adt_net_52247_\);
    
    \I2.PIPE8_DT_16_0l15r\ : MUX2H
      port map(A => \I2.PIPE8_DTl15r_net_1\, B => 
        \I2.PIPE7_DTl15r_net_1\, S => 
        \I2.N_565_0_adt_net_855736__net_1\, Y => \I2.N_581\);
    
    \I1.un1_sbyte13_i_i_i_o2\ : OR2FT
      port map(A => \I1.sstatel3r_net_1\, B => PULSEl6r, Y => 
        \I1.N_329\);
    
    \I2.DT_TEMPl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_776_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl15r_net_1\);
    
    \I2.DTE_21_1_IV_0_0L17R_1224\ : AO21
      port map(A => \I2.DT_TEMPl17r_net_1\, B => \I2.N_4038\, C
         => \I2.DTE_21_1l17r_adt_net_36146_\, Y => 
        \I2.DTE_21_1l17r_adt_net_36153_\);
    
    \I2.OFFSET_37_26l1r\ : MUX2L
      port map(A => \REGl222r\, B => \I2.N_828\, S => 
        \I2.PIPE7_DTl26r_net_1\, Y => \I2.N_836\);
    
    \I3.REG_1_277\ : MUX2H
      port map(A => VDB_inl5r, B => \I3.REGl96r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_277_0\);
    
    \I2.LSRAM_IN_403\ : MUX2L
      port map(A => \I2.PIPE5_DTl19r_net_1\, B => 
        \I2.LSRAM_INl19r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_403_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I110_un1_Y\ : AND3
      port map(A => \I2.N466\, B => 
        \I2.I110_un1_Y_adt_net_71212_\, C => \I2.N333\, Y => 
        \I2.I110_un1_Y\);
    
    \I2.PIPE5_DT_6l16r\ : MUX2L
      port map(A => \I2.PIPE4_DTl16r_net_1\, B => \I2.N_1085\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\, Y
         => \I2.PIPE5_DT_6l16r_net_1\);
    
    \I2.DTO_9_IVL15R_1138\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        B => \I2.DTE_2_1l15r_net_1\, Y => 
        \I2.DTO_9l15r_adt_net_31888_\);
    
    \I2.PIPE7_DTL26R_2897\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_351\);
    
    \I2.SUB9_1_ADD_18x18_fast_I0_CO1\ : AND2
      port map(A => \I2.ca\, B => \I2.G_1_5\, Y => \I2.N225\);
    
    \I2.DTE_21_1_IV_0L28R_1236\ : OAI21FTF
      port map(A => \I2.STATE2l3r_net_1\, B => 
        \I2.DTO_9_iv_ml28r_adt_net_857__net_1\, C => 
        \I2.DTE_21_1l28r_adt_net_36758_\, Y => 
        \I2.DTE_21_1l28r_adt_net_36759_\);
    
    \I3.REG_1_208\ : MUX2L
      port map(A => VDB_inl27r, B => \I3.REGl160r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\, Y => 
        \I3.REG_1_208_0\);
    
    \I2.PIPE1_DT_42_1_IVL20R_1391\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_340\, B => 
        \I2.EVNT_NUMl4r_net_1\, Y => 
        \I2.PIPE1_DT_42l20r_adt_net_47055_\);
    
    \I2.PIPE1_DT_42_1_IVL6R_1488\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855228__net_1\, B => 
        \I2.MIC_ERR_REGSl6r_net_1\, C => 
        \I2.PIPE1_DT_42l6r_adt_net_50938_\, Y => 
        \I2.PIPE1_DT_42l6r_adt_net_50939_\);
    
    \I2.DTE_21_1_iv_0l24r\ : AO21
      port map(A => \I2.DTE_1l24r_Rd1__net_1\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835180_Rd1__net_1\, 
        C => \I2.DTE_21_1l24r_adt_net_37175_Rd1__net_1\, Y => 
        \I2.DTE_21_1l24r_Rd1_\);
    
    \I3.PIPEAl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_235_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl4r_net_1\);
    
    \I3.REGMAPl9r_adt_net_854320_\ : BFR
      port map(A => \I3.REGMAPL9R_783\, Y => 
        \I3.REGMAPl9r_adt_net_854320__net_1\);
    
    \I2.PIPE10_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_631_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl26r_net_1\);
    
    \I2.OFFSET_37_8l5r\ : MUX2L
      port map(A => \REGl362r\, B => \REGl298r\, S => 
        \I2.PIPE7_DTL27R_69\, Y => \I2.N_696\);
    
    \I2.PIPE9_DT_286\ : MUX2L
      port map(A => \I2.PIPE9_DTl17r_net_1\, B => 
        \I2.PIPE8_DTl17r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_286_net_1\);
    
    REGl311r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_212_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl311r\);
    
    \I2.RAMAD_4l12r\ : MUX2L
      port map(A => \I2.N_539\, B => 
        \I1.PAGECNTl4r_adt_net_835120_Rd1__net_1\, S => 
        LOAD_RES_1, Y => \I2.RAMAD_4l12r_net_1\);
    
    \I1.BITCNT_317\ : MUX2L
      port map(A => \I1.BITCNTl0r_net_1\, B => \I1.N_1199\, S => 
        \I1.N_68\, Y => \I1.BITCNT_317_net_1\);
    
    \I3.VDBOFFA_31_IV_0L0R_2623\ : AND2
      port map(A => \REGl277r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        Y => \I3.VDBoffa_31l0r_adt_net_164614_\);
    
    \I2.PIPE1_DT_30l18r\ : MUX2L
      port map(A => \I2.TDCDBSl18r_net_1\, B => 
        \I2.TDCDBSl16r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, Y
         => \I2.PIPE1_DT_30l18r_net_1\);
    
    \I2.PIPE1_DT_12l20r\ : MUX2L
      port map(A => \I2.TDCDASl20r_net_1\, B => 
        \I2.TDCDASl18r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092__net_1\, Y
         => \I2.PIPE1_DT_12l20r_net_1\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855432_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__22\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\);
    
    \I2.OFFSET_37_20l2r\ : MUX2L
      port map(A => \I2.N_781\, B => \I2.N_773\, S => 
        \I2.PIPE7_DTL26R_359\, Y => \I2.N_789\);
    
    \I3.PIPEA1_12l4r\ : AND2
      port map(A => DPR_cl4r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854508__net_1\, Y => 
        \I3.PIPEA1_12l4r_net_1\);
    
    \I1.PAGECNT_n2_0_0_o2\ : AND2
      port map(A => \I1.PAGECNT_326_202\, B => 
        \I1.PAGECNT_327_203\, Y => \I1.N_300_Ra1_\);
    
    \I2.STATE5l3r\ : DFFS
      port map(CLK => CLK_c, D => \I2.STATE5_ns_i_0l0r_net_1\, 
        SET => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.STATE5l3r_net_1\);
    
    \I3.VDBI_57_IV_0_0L0R_2284\ : AND2
      port map(A => \I3.N_2036\, B => 
        \I3.VDBi_57l0r_adt_net_1621__net_1\, Y => 
        \I3.VDBi_57l0r_adt_net_146601_\);
    
    \I3.VDBI_57_0_IV_0_0L24R_2156\ : AND2
      port map(A => \I3.PIPEAl24r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l24r_adt_net_138807_\);
    
    \I2.PIPE8_DT_21l26r\ : MUX2H
      port map(A => \I2.PIPE7_DTl26r_net_1\, B => 
        \I2.LSRAM_OUTl26r\, S => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l26r_net_1\);
    
    \I2.DTO_16_1_IV_0_0L16R_1134\ : AND2
      port map(A => \I2.N_4671_adt_net_854596__net_1\, B => 
        \I2.DT_TEMPl16r_net_1\, Y => 
        \I2.DTO_16_1l16r_adt_net_31706_\);
    
    \I3.REGMAP_i_0_il32r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un141_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il32r_net_1\);
    
    \I2.DTO_1_904\ : MUX2L
      port map(A => \I2.DTO_1l30r_net_1\, B => 
        \I2.DTO_16_1_ivl30r_net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => \I2.DTO_1_904_net_1\);
    
    \I3.PIPEA_i_0l31r\ : INV
      port map(A => CLEAR_STAT, Y => CLEAR_STAT_i_0);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I181_Y\ : XOR2
      port map(A => \I2.N519_0\, B => 
        \I2.ADD_21x21_fast_I181_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l11r\);
    
    \I5.SBYTE_9_il3r\ : MUX2L
      port map(A => \I5.COMMANDl11r_net_1\, B => 
        \I5.SBYTEl2r_net_1\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.N_20\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I110_UN1_Y_1664\ : AND2FT
      port map(A => \I2.N290\, B => \I2.N294\, Y => 
        \I2.I110_un1_Y_adt_net_71212_\);
    
    \I2.PIPE2_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl8r_net_1\);
    
    \I1.REG_15_sqmuxa_adt_net_1457_\ : OR3
      port map(A => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__197\, 
        B => \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Rd1__net_1\, C
         => \I1.REG_15_sqmuxa_adt_net_109461_Rd1__net_1\, Y => 
        \I1.REG_15_sqmuxa_adt_net_1457__net_1\);
    
    REGl245r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_146_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl245r\);
    
    REGl248r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_149_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl248r\);
    
    \I2.PIPE7_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl15r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl15r_net_1\);
    
    \I2.N_4644_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4644\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4644_Rd1__net_1\);
    
    \I1.SSTATE_NS_0_IV_0_I_M2L3R_1767\ : AND2FT
      port map(A => \I1.N_321_adt_net_855540__net_1\, B => 
        \I1.sstatel8r_net_1\, Y => \I1.N_420_i_adt_net_107486_\);
    
    \I3.VDBOFFA_31_IV_0L5R_2530\ : AND2
      port map(A => \REGl202r\, B => \I3.REGMAPl22r_net_1\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163652_\);
    
    \I2.DTO_16_1_IVL14R_1147\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855680__net_1\, B => 
        \I2.DTO_9l14r\, Y => \I2.DTO_16_1l14r_adt_net_32194_\);
    
    \I3.un1_NOEDTKi_0_sqmuxa_0_o3\ : OR2
      port map(A => \I3.un1_NOEDTKi_0_sqmuxa_adt_net_4101__net_1\, 
        B => \I3.un1_NOEDTKi_0_sqmuxa_adt_net_159270_\, Y => 
        \I3.un1_NOEDTKi_0_sqmuxa\);
    
    \I2.G_EVNT_NUM_i_0_il0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_934_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUM_i_0_il0r_net_1\);
    
    \I2.CRC32_12_i_x2l12r\ : XOR2FT
      port map(A => \I2.CRC32l12r_net_1\, B => \I2.N_3957_i_i\, Y
         => \I2.N_116_i_i_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I16_G0N_0_a2\ : AND2
      port map(A => \I2.RAMDT4L5R_819\, B => 
        \I2.PIPE4_DTl16r_net_1\, Y => \I2.N307\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I94_Y\ : NAND2
      port map(A => \I2.N305_0\, B => \I2.N309_0\, Y => \I2.N348\);
    
    \I2.DTO_9_ivl7r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl7r_net_1\, 
        C => \I2.DTO_9l7r_adt_net_33668_\, Y => \I2.DTO_9l7r\);
    
    \I1.SSTATE_NS_1_IV_0_0L7R_1769\ : OAI21TTF
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.N_329\, C => \I1.sstate_nsl7r_adt_net_107573_\, Y => 
        \I1.sstate_nsl7r_adt_net_107578_\);
    
    FBOUTl1r : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_59_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \FBOUTl1r\);
    
    \I2.PIPE10_DT_617\ : MUX2L
      port map(A => \I2.PIPE10_DTl12r_net_1\, B => 
        \I2.PIPE9_DTl12r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_617_net_1\);
    
    \I1.PAGECNTl3r_adt_net_835116_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.PAGECNT_324_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNTl3r_adt_net_835116_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L0R_2626\ : AO21
      port map(A => \REGl189r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.VDBoffa_31l0r_adt_net_164598_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164639_\);
    
    \I3.REG_1l133r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_181_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl133r\);
    
    REGl310r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_211_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl310r\);
    
    \I5.DATA_12l9r\ : MUX2L
      port map(A => REGl126r, B => \I5.SBYTEl1r_net_1\, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l9r_net_1\);
    
    \I2.PIPE10_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_635_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl30r_net_1\);
    
    \I2.DT_SRAMl20r\ : MUX2L
      port map(A => \I2.N_888\, B => \I2.PIPE2_DTl20r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668__net_1\, 
        Y => \I2.DT_SRAMl20r_net_1\);
    
    \I3.PIPEA_8_0l8r\ : MUX2L
      port map(A => DPR_cl8r, B => \I3.PIPEA1l8r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855352__net_1\, Y => \I3.N_217\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I99_Y_1660\ : AND2
      port map(A => \I2.N308\, B => \I2.N304\, Y => 
        \I2.N463_adt_net_70886_\);
    
    \I2.SUB8_523_2741\ : AOI21TTF
      port map(A => \I2.N288_0\, B => 
        \I2.N475_adt_net_4127__net_1\, C => 
        \I2.SUB8_523_adt_net_566476_\, Y => 
        \I2.SUB8_523_adt_net_670059_\);
    
    \I3.REG_44_i_0l83r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_327\, Y => \I3.N_1629\);
    
    \I5.BITCNTE_0_A2_0_912\ : OA21FTT
      port map(A => \I5.N_77\, B => \I5.N_75\, C => TICKL0R_556, 
        Y => \I5.BITCNTe_adt_net_9456_\);
    
    \I2.LEAD_FLAG6_7_i_0l2r\ : AOI21
      port map(A => \I2.N_217\, B => \I2.N_484\, C => \I2.N_222\, 
        Y => \I2.N_4533_adt_net_64364_\);
    
    \I2.DTO_16_1_IV_0L17R_1130\ : AND2
      port map(A => \I2.N_4671_adt_net_854596__net_1\, B => 
        \I2.DT_TEMPl17r_net_1\, Y => 
        \I2.DTO_16_1l17r_adt_net_31520_\);
    
    \I2.TOKOUTBS_1522\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKOUTBS_3_i_net_1\, 
        Q => \I2.TOKOUTBS_629\);
    
    \I3.STATE1_0l9r_1157\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL9R_419\);
    
    \I2.FID_7_0_IV_0L1R_1732\ : NOR2FT
      port map(A => \I2.STATE3l7r_net_1\, B => REGl49r, Y => 
        \I2.FID_7_0_iv_0l1r_adt_net_93441_\);
    
    \I2.PIPE8_DT_16_0l11r\ : MUX2H
      port map(A => \I2.PIPE8_DTl11r_net_1\, B => 
        \I2.PIPE7_DTl11r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_577\);
    
    \I2.TDCDBSl19r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl19r, Q => 
        \I2.TDCDBSl19r_net_1\);
    
    \I2.DTE_21_1_0_IV_1L30R_1229\ : NOR2
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855192__net_1\, 
        B => \I2.DT_TEMPl30r_net_1\, Y => 
        \I2.DTE_21_1_0_iv_1l30r_adt_net_36505_\);
    
    TDCDB_padl29r : IB33
      port map(PAD => TDCDB(29), Y => TDCDB_cl29r);
    
    \I2.N507_adt_net_347770_\ : OR2FT
      port map(A => \I2.N_112_2\, B => 
        \I2.N507_adt_net_283110__net_1\, Y => 
        \I2.N507_adt_net_347770__net_1\);
    
    \I1.REG_74_5_404_m1_e_0_901\ : NOR2FT
      port map(A => \I1.PAGECNT_0l8r_adt_net_834720_Rd1__net_1\, 
        B => \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__362\, Y => 
        \I1.REG_74_5_404_M1_E_0_279\);
    
    \I3.VDBOFFB_30_IV_0L2R_2447\ : AO21
      port map(A => \REGl383r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l2r_adt_net_162702_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162740_\);
    
    \I1.PAGECNT_319\ : MUX2H
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        B => \I1.N_1379\, S => 
        \I1.PAGECNTe_adt_net_854892__net_1\, Y => 
        \I1.PAGECNT_319_net_1\);
    
    \I3.TCNT4_n2\ : XOR2
      port map(A => \I3.TCNT4_i_0_il2r_net_1\, B => 
        \I3.TCNT4_c1_net_1\, Y => \I3.TCNT4_n2_net_1\);
    
    \I5.sstate2se_0_0\ : AO21FTT
      port map(A => \I5.N_464\, B => \I5.sstate2l4r_net_1\, C => 
        \I5.sstate2_ns_el1r_adt_net_8563_\, Y => 
        \I5.sstate2_ns_el1r\);
    
    \I3.VDBil26r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_366_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil26r_net_1\);
    
    \I3.SINGCYC\ : DFFC
      port map(CLK => CLK_c, D => \I3.SINGCYC_115_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.SINGCYC_net_1\);
    
    \I2.PIPE2_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl5r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl5r_net_1\);
    
    \I2.REG_1_n3_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855784__net_1\, B
         => REGl35r, Y => \I2.REG_1_n3_0_net_1\);
    
    \I2.PIPE8_DT_16l18r\ : AND2
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855164__net_1\, B => 
        \I2.N_584\, Y => \I2.PIPE8_DT_16l18r_net_1\);
    
    \I2.DTE_21_1_IV_0_0L4R_1331\ : AND2
      port map(A => \I2.DT_SRAMl4r_net_1\, B => 
        \I2.N_199_0_ADT_NET_1054__37\, Y => 
        \I2.DTE_21_1l4r_adt_net_39199_\);
    
    \I2.un1_PIPE1_DT_1_sqmuxa_2_0\ : OA21TTF
      port map(A => \I2.un1_PIPE1_DT_1_sqmuxa_2_adt_net_20482_\, 
        B => \I2.N_3902_adt_net_20437_\, C => 
        \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\, Y => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\);
    
    \I1.REG_74_0_ivl281r\ : AO21
      port map(A => \REGl281r\, B => \I1.N_153\, C => 
        \I1.REG_74l281r_adt_net_122635_\, Y => \I1.REG_74l281r\);
    
    \I2.BNCID_VECTROR_1425\ : OR2
      port map(A => \I2.BNCID_VECTror_adt_net_48461_\, B => 
        \I2.BNCID_VECTror_adt_net_48463_\, Y => 
        \I2.BNCID_VECTror_adt_net_48422_\);
    
    \REG_i_il5r_adt_net_855552_\ : BFR
      port map(A => \REG_i_il5r_adt_net_855560__net_1\, Y => 
        \REG_i_il5r_adt_net_855552__net_1\);
    
    \I1.REG_74_0_iv_0_0l255r\ : AO21
      port map(A => \REGl255r\, B => \I1.N_658\, C => 
        \I1.REG_74l255r_adt_net_125228_\, Y => \I1.REG_74l255r\);
    
    \I2.CHB_DATA8_2_I_1693\ : AND2FT
      port map(A => \I2.PIPE7_DTl28r_net_1\, B => \I2.N_4402\, Y
         => \I2.N_4397_adt_net_90034_\);
    
    \I2.L2TYPEl3r_1554\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_592_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL3R_661\);
    
    \I1.REG_1_77\ : MUX2H
      port map(A => \REGl176r\, B => \I1.REG_74l176r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\, Y => 
        \I1.REG_1_77_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2390\ : AND2
      port map(A => \REGl306r\, B => \I3.REGMAPl35r_net_1\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162148_\);
    
    \I2.OFFSET_37_28l3r\ : MUX2L
      port map(A => \I2.N_846\, B => \I2.N_798\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_854\);
    
    \I2.L2TYPE_4_IL0R_1642\ : AND2
      port map(A => \I2.L2TYPEl0r_net_1\, B => 
        \I2.N_4452_adt_net_68713_\, Y => 
        \I2.N_4452_adt_net_68756_\);
    
    \I2.MIC_REG3_319\ : MUX2H
      port map(A => \I2.MIC_REG3l2r_net_1\, B => 
        \I2.MIC_REG3l3r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG3_319_net_1\);
    
    \I2.PIPE5_DT_694\ : MUX2L
      port map(A => \I2.PIPE5_DTl18r_net_1\, B => 
        \I2.PIPE5_DT_6l18r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_694_net_1\);
    
    \I2.I_1341_G_1\ : XOR2FT
      port map(A => \I2.OFFSETL6R_673\, B => \I2.SUB8l9r_net_1\, 
        Y => \I2.G_1_0\);
    
    NOESRAMO_pad : OB33PH
      port map(PAD => NOESRAMO, A => NOESRAMO_c);
    
    \I2.DTE_21_1_iv_0_0_18_m7\ : OR3
      port map(A => \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35891_\, 
        B => \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35904_\, C => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35905_\, Y => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0\);
    
    \I2.PIPE7_DTL27R_2776\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_69\);
    
    \I2.un1_STATE1_21_0_0\ : OR3FTT
      port map(A => \I2.N_3287_i_0\, B => \I2.STATE1l14r_net_1\, 
        C => \I2.N_3890\, Y => \I2.un1_STATE1_21\);
    
    \I3.REG_1_I_S_I_IL4R_1041\ : AOI21
      port map(A => \I3.REG2l4r_net_1\, B => \I3.REG3L4R_431\, C
         => \I3.REG1l4r_net_1\, Y => \I3.N_203_adt_net_24461_\);
    
    \I3.REG_1l73r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_174_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl73r);
    
    \I2.resyn_0_I2_TRGCNT_c1_i\ : OAI21
      port map(A => \I2.un9_tdctrgi_i_0\, B => \I2.N_3765\, C => 
        \I2.N_3796\, Y => \I2.N_3762\);
    
    \I2.OFFSETl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_560_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl0r_net_1\);
    
    \I2.REG_1_c9_i\ : OAI21TTF
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => \I2.N_3853\, C => \I2.N_3838_adt_net_101306_\, Y => 
        \I2.N_3838\);
    
    \I1.REG_7_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_254\, B => \I1.N_243\, Y => 
        \I1.REG_7_sqmuxa\);
    
    \I2.NWPIPE8_0_0\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, 
        SET => CLEAR_STAT_i_0, Q => \I2.NWPIPE8_i_0_i_0_0\);
    
    \I2.G_EVNT_NUM_n10_0_a2_0_0\ : NOR2
      port map(A => EV_RES_C_568, B => \I2.G_EVNT_NUMl10r_net_1\, 
        Y => \I2.G_EVNT_NUM_n10_0_a2_0_0_i\);
    
    \I3.REG_1_171\ : MUX2L
      port map(A => VDB_inl22r, B => REGl70r, S => 
        \I3.N_1935_adt_net_855320__net_1\, Y => \I3.REG_1_171_0\);
    
    \I3.VDBi_55l4r\ : MUX2H
      port map(A => \I3.VDBil4r_net_1\, B => \I3.RAMDTSl4r_net_1\, 
        S => \I3.N_57_i_0_0_adt_net_854688__net_1\, Y => 
        \I3.VDBi_55l4r_net_1\);
    
    \I2.SUB9l15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_583_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9_i_0_il15r\);
    
    \I3.RAMAD_VME_37\ : MUX2H
      port map(A => RAMAD_VMEl13r, B => \I3.REGl96r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_37_net_1\);
    
    \I2.BNCID_VECT_tile_0_WADDR_REG1l1r\ : DFF
      port map(CLK => CLK_c, D => \I2.TRGARRl1r_net_1\, Q => 
        \I2.WADDR_REG1l1r\);
    
    \I2.STATEE_ILLEGAL_1027\ : AND2
      port map(A => \I2.STATEe_ipl2r\, B => \I2.STATEe_ipl3r\, Y
         => \I2.N_3457_ip_adt_net_23071_\);
    
    \I2.PIPE1_DT_42_1_ivl6r\ : OR3
      port map(A => \I2.PIPE1_DT_42l6r_adt_net_50930_\, B => 
        \I2.PIPE1_DT_42l6r_adt_net_50939_\, C => 
        \I2.PIPE1_DT_42l6r_adt_net_50940_\, Y => 
        \I2.PIPE1_DT_42l6r\);
    
    \I3.N_48_i_0_o2\ : NOR3FTT
      port map(A => \I3.N_177_adt_net_134570_\, B => 
        \I3.REGMAP_I_0_IL36R_529\, C => \I3.REGMAPL35R_528\, Y
         => \I3.N_177\);
    
    \I2.BNCID_VECTror_8_tz_0\ : AO21
      port map(A => \I2.BNCID_VECTra13_1_net_1\, B => 
        \I2.BNCID_VECTro_9\, C => 
        \I2.BNCID_VECTror_8_tz_0_i_adt_net_48007_\, Y => 
        \I2.BNCID_VECTror_8_tz_0_i\);
    
    \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_4066_\ : AO21
      port map(A => \I3.VDBil0r_net_1\, B => \I3.N_2048\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146205__net_1\, Y
         => \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_4066__net_1\);
    
    \I3.PIPEA_8_0l17r\ : MUX2L
      port map(A => DPR_cl17r, B => \I3.PIPEA1l17r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855348__net_1\, Y => \I3.N_226\);
    
    \I1.REG_1_154\ : MUX2H
      port map(A => \REGl253r\, B => \I1.REG_74l253r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_154_net_1\);
    
    REGl232r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_133_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl232r\);
    
    \I2.EVNT_NUMl0r_1134\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_963_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUML0R_396\);
    
    \I2.DTO_16_1_IV_1L30R_1068\ : NOR2
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608__net_1\, 
        B => \I2.DT_TEMPl30r_net_1\, Y => 
        \I2.DTO_16_1_iv_1l30r_adt_net_28466_\);
    
    \I1.REG_1_199\ : MUX2H
      port map(A => \REGl298r\, B => \I1.REG_74l298r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\, Y => 
        \I1.REG_1_199_net_1\);
    
    \I2.DT_SRAM_i_m2l13r\ : MUX2L
      port map(A => \I2.N_4046\, B => \I2.PIPE2_DTl13r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.N_4048\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I199_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl3r\, B => 
        \I2.PIPE7_DTl3r_net_1\, Y => \I2.SUB_21x21_fast_I199_Y_0\);
    
    \I3.VDBi_57_0_ivl22r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l22r_net_1\, C
         => \I3.VDBi_57l22r_adt_net_139087_\, Y => 
        \I3.VDBi_57l22r\);
    
    \I2.PIPE4_DTL10R_3037\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL10R_791\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I22_G0N\ : AND2FT
      port map(A => \I2.LSRAM_OUTl1r\, B => \I2.PIPE7_DTL1R_703\, 
        Y => \I2.N233\);
    
    REGl265r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_166_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl265r\);
    
    \I3.REG_1_223\ : MUX2L
      port map(A => VDB_inl10r, B => REGl416r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_223_0\);
    
    \I2.DTO_16_1_IV_0L9R_1176\ : AO21
      port map(A => \I2.N_197_154\, B => \I2.N_4047\, C => 
        \I2.DTO_16_1l9r_adt_net_33242_\, Y => 
        \I2.DTO_16_1l9r_adt_net_33252_\);
    
    REGl268r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_169_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl268r\);
    
    \I2.RAMDT4L5R_2808\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_136\);
    
    \I2.PIPE1_DT_30l11r\ : MUX2L
      port map(A => \I2.TDCDBSl11r_net_1\, B => 
        \I2.TDCDBSl9r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, Y
         => \I2.PIPE1_DT_30l11r_net_1\);
    
    \I2.PIPE9_DT_282\ : MUX2L
      port map(A => \I2.PIPE9_DTl13r_net_1\, B => 
        \I2.PIPE8_DTl13r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_282_net_1\);
    
    \I5.BITCNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.BITCNT_86_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.BITCNT_c0\);
    
    \I1.REG_74_0_IVL297R_1921\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l297r_adt_net_121126_\);
    
    \I2.STATE1_ns_0l5r_adt_net_855812_\ : BFR
      port map(A => \I2.STATE1_ns_0l5r\, Y => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\);
    
    \I1.sstate_ns_0_iv_0_0_o2l2r\ : OR2
      port map(A => \I1.N_317_Rd1__net_1\, B => 
        \I1.N_321_adt_net_105403_\, Y => \I1.N_321\);
    
    \I1.un1_sbyte13_i_i_i_1\ : OR3
      port map(A => \PULSEl0r_adt_net_854532__net_1\, B => 
        \I1.N_598\, C => \I1.un1_sbyte13_i_i_i_1_adt_net_108267_\, 
        Y => \I1.un1_sbyte13_i_i_i_1_net_1\);
    
    \I2.FID_7_0_IVL21R_994\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl69r, C => 
        \I2.FID_7l21r_adt_net_19397_\, Y => 
        \I2.FID_7l21r_adt_net_19405_\);
    
    \I2.ROFFSETe_0_adt_net_27184_\ : OAI21FTF
      port map(A => \I2.STATE3L2R_413\, B => 
        \I2.STOP_RDSRAM_net_1\, C => \I2.N_4676\, Y => 
        \I2.ROFFSETe_0_adt_net_27184__net_1\);
    
    \I2.BNCID_VECTwa13_1\ : NOR2FT
      port map(A => \I2.TRGARRl0r_net_1\, B => 
        \I2.TRGARRl1r_net_1\, Y => \I2.BNCID_VECTwa13_1_net_1\);
    
    \I2.N436_adt_net_1185_\ : OR3FTT
      port map(A => \I2.N268\, B => 
        \I2.SUB8l15r_adt_net_855572__net_1\, C => \I2.N290\, Y
         => \I2.N436_adt_net_1185__net_1\);
    
    \I3.REGMAP_i_0_a2l52r\ : NOR3FFT
      port map(A => \I3.UN1_REGMAP_34_123\, B => 
        \I3.N_638_adt_net_134647_\, C => \I3.N_2017_118\, Y => 
        \I3.N_638\);
    
    \I1.REG_74_0_IVL385R_1808\ : AND2
      port map(A => \FBOUTl4r\, B => \I1.REG_28_sqmuxa\, Y => 
        \I1.REG_74l385r_adt_net_111577_\);
    
    \I2.TDCDBSl31r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl31r, Q => 
        \I2.TDCDBSl31r_net_1\);
    
    \I3.VDBil4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_344_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil4r_net_1\);
    
    \I2.resyn_0_I2_TRGCNT_n3\ : XOR2FT
      port map(A => \I2.N_3763\, B => \I2.TRGCNT_n3_0\, Y => 
        \I2.TRGCNT_n3\);
    
    \I2.DTO_1l19r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l19r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l19r_Rd1__net_1\);
    
    \I3.REG_44_i_a2_0l89r\ : NOR2
      port map(A => VDB_inl6r, B => \I3.N_98\, Y => \I3.N_1673\);
    
    \I5.REG_1_54_924\ : NOR3FTT
      port map(A => \I5.sstate1l13r_net_1\, B => 
        \I5.PULSE_FL_net_1\, C => \I5.PULSE_I2C_net_1\, Y => 
        \I5.REG_1_54_adt_net_11847_\);
    
    REGl339r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_240_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl339r\);
    
    \I2.OFFSET_37_9l1r\ : MUX2L
      port map(A => \REGl390r\, B => \REGl326r\, S => 
        \I2.PIPE7_DTL27R_84\, Y => \I2.N_700\);
    
    \I2.LSRAM_IN_397\ : MUX2L
      port map(A => \I2.PIPE5_DTl13r_net_1\, B => 
        \I2.LSRAM_INl13r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_397_net_1\);
    
    \I2.DTE_1_862\ : MUX2L
      port map(A => \I2.DTE_1l24r_Rd1__net_1\, B => 
        \I2.DTE_21_1l24r_Rd1_\, S => 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\, Y => 
        \I2.DTE_1l24r\);
    
    \I1.ISCK_0_sqmuxa_0_0_a2_1232\ : NAND3FFT
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__862\, B => 
        \I1.N_359\, C => \I1.sstatel4r_net_1\, Y => 
        \I1.N_656_494\);
    
    \I3.un47_reg_ads_0_a2_0_a3\ : NOR3
      port map(A => \I3.N_547\, B => \I3.N_551\, C => 
        \I3.un47_reg_ads_1\, Y => 
        \I3.un47_reg_ads_0_a2_0_a3_net_1\);
    
    DS0B_pad : IB33
      port map(PAD => DS0B, Y => DS0B_c);
    
    \I2.PIPE10_DT_626\ : MUX2L
      port map(A => \I2.PIPE10_DTl21r_net_1\, B => 
        \I2.PIPE9_DTl21r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_626_net_1\);
    
    \I2.PIPE10_DT_609\ : MUX2L
      port map(A => \I2.PIPE10_DTl4r_net_1\, B => 
        \I2.PIPE9_DTl4r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_609_net_1\);
    
    \I2.OFFSETl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_566_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl6r_net_1\);
    
    \I2.MIC_ERR_REGS_340\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl12r_net_1\, B => 
        \I2.MIC_ERR_REGSl11r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\, Y => 
        \I2.MIC_ERR_REGS_340_net_1\);
    
    \I3.VDBI_57_IV_0_0L7R_2232\ : AO21
      port map(A => \I3.VDBil7r_net_1\, B => \I3.N_2048\, C => 
        \I3.VDBi_57l7r_adt_net_143099_\, Y => 
        \I3.VDBi_57l7r_adt_net_143112_\);
    
    \I2.STATE4_ns_i_0_1l1r\ : NOR2
      port map(A => \I2.N_4481\, B => REGl2r, Y => \I2.N_3376_1\);
    
    \I2.N_3287_i_0_a2\ : NAND2
      port map(A => \I2.N_3882\, B => \I2.STATE1L18R_627\, Y => 
        \I2.N_3287_i_0\);
    
    \I2.DT_SRAM_0l23r\ : MUX2L
      port map(A => \I2.PIPE10_DTl23r_net_1\, B => 
        \I2.PIPE5_DTL23R_624\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, Y => 
        \I2.N_891\);
    
    \I2.CRC32_12_0_0_x2l25r\ : XOR2FT
      port map(A => \I2.CRC32l25r_net_1\, B => \I2.N_4349_i_i\, Y
         => \I2.N_42_i_0_i_0\);
    
    \I2.N346_adt_net_69448_\ : OA21
      port map(A => \I2.ca_0_and2\, B => \I2.G_1_4\, C => 
        \I2.N225\, Y => \I2.N346_adt_net_69448__net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I136_Y_0_O2_M4_E_2_1568\ : 
        AND3
      port map(A => \I2.N_57_0\, B => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_2_adt_net_56513_\, C
         => \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_i_1\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_2_adt_net_56515_\);
    
    \I1.REG_74_0_IVL306R_1912\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l306r_adt_net_120352_\);
    
    \I2.RAMAD1_12l8r\ : MUX2L
      port map(A => \I2.TDCDASl6r_net_1\, B => 
        \I2.TDCDBSl6r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855180__net_1\, Y => 
        \I2.RAMAD1_12l8r_net_1\);
    
    \I3.PIPEA_8l28r\ : OR2FT
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854484__net_1\, B => 
        \I3.N_237\, Y => \I3.PIPEA_8l28r_net_1\);
    
    \I3.PIPEA_8_0l9r\ : MUX2L
      port map(A => DPR_cl9r, B => \I3.PIPEA1l9r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855352__net_1\, Y => \I3.N_218\);
    
    \I2.BNC_IDl8r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_45_0\, CLR => 
        \I2.N_4619_i_0\, SET => \I2.N_4612_i_0\, Q => 
        \I2.BNC_IDl8r_net_1\);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854232_\ : BFR
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854248__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854232__net_1\);
    
    \I5.BITCNT_n2_i\ : OA21TTF
      port map(A => \I5.BITCNTl2r_net_1\, B => \I5.N_65\, C => 
        \I5.N_144\, Y => \I5.N_54_adt_net_9598_\);
    
    \I2.un28_sram_empty_14_0\ : MUX2L
      port map(A => \I2.N_632\, B => \I2.N_629\, S => 
        \I2.RPAGEL13R_609\, Y => \I2.N_633\);
    
    \I2.STATE2_ns_i_0_o2_0_0_m7_i\ : AO21
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__488\, B => 
        \I2.N_4273_adt_net_20831_\, C => 
        \I2.N_4273_adt_net_20928_\, Y => \I2.N_4273\);
    
    \I2.CRC32l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_797_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l2r_net_1\);
    
    \I2.FID_7_0_IVL18R_955\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl18r_net_1\, 
        Y => \I2.FID_7l18r_adt_net_17611_\);
    
    \I3.UN221_REG_ADS_0_A2_0_A3_2648\ : NOR2
      port map(A => \I3.VASl12r_net_1\, B => \I3.N_562\, Y => 
        \I3.un221_reg_ads_0_a2_0_a3_adt_net_165933_\);
    
    \I2.LSRAM_INl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_395_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl11r_net_1\);
    
    \I3.TCNT2_391\ : MUX2H
      port map(A => \I3.TCNT2l5r_net_1\, B => \I3.TCNT2_n5_net_1\, 
        S => TICKl0r, Y => \I3.TCNT2_391_net_1\);
    
    \I2.DTE_21_1l22r_adt_net_37395_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.DTE_21_1l22r_adt_net_37395_\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.DTE_21_1l22r_adt_net_37395_Rd1__net_1\);
    
    \I3.UN2_VSEL_1_I_0_A2_2101\ : OR3FFT
      port map(A => IACKB_c, B => AMB_cl3r, C => AMB_cl2r, Y => 
        \I3.N_2055_adt_net_134991_\);
    
    \I1.REG_1_267\ : MUX2H
      port map(A => \REGl366r\, B => \I1.REG_74l366r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_267_net_1\);
    
    \I3.STATE1_NS_1_IV_0L2R_2096\ : NOR3FFT
      port map(A => \I3.N_437\, B => 
        \I3.STATE1_nsl2r_adt_net_1586__net_1\, C => \I3.N_276\, Y
         => \I3.STATE1_nsl2r_adt_net_134784_\);
    
    \I2.DT_TEMP_792\ : MUX2H
      port map(A => \I2.DT_TEMPl31r_net_1\, B => 
        \I2.DT_TEMP_7l31r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_792_net_1\);
    
    \I2.BNCID_VECTrff_2_263_0\ : AO21
      port map(A => \I2.BNCID_VECTrff_3_262_0_a2_0\, B => 
        \I2.BNCID_VECTwa14_1_net_1\, C => \I2.BNCID_VECTro_2\, Y
         => \I2.BNCID_VECTrff_2_263_0_net_1\);
    
    \I2.DTO_16_1_IV_0_0L26R_1082\ : AND2
      port map(A => \I2.N_4671_adt_net_854592__net_1\, B => 
        \I2.DT_TEMPl26r_net_1\, Y => 
        \I2.DTO_16_1l26r_adt_net_29426_\);
    
    \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1\ : OR2
      port map(A => \I1.PAGECNT_325_net_1\, B => 
        \I1.PAGECNT_326_net_1\, Y => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Ra1_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I109_un1_Y\ : AND3
      port map(A => \I2.N463\, B => 
        \I2.I109_un1_Y_adt_net_70914_\, C => \I2.N331\, Y => 
        \I2.I109_un1_Y\);
    
    \I2.G_EVNT_NUM_924\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl10r_net_1\, B => 
        \I2.G_EVNT_NUM_n10\, S => \I2.N_3769\, Y => 
        \I2.G_EVNT_NUM_924_net_1\);
    
    TDCTRG_pad : OB33PH
      port map(PAD => TDCTRG, A => TDCTRG_c);
    
    REGl272r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_173_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl272r\);
    
    \I2.TDCDASl4r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl4r, Q => 
        \I2.TDCDASl4r_net_1\);
    
    \I2.CRC32_12_il16r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_112_i_i_0\, Y => 
        \I2.N_3933\);
    
    \I3.VDBOFFA_31_IV_0L7R_2507\ : OR2
      port map(A => \I3.VDBoffa_31l7r_adt_net_163311_\, B => 
        \I3.VDBoffa_31l7r_adt_net_163312_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163317_\);
    
    \I3.REGMAP_I_0_A2L52R_2093\ : AND3
      port map(A => \I3.N_638_adt_net_134639_\, B => \I3.N_590\, 
        C => \I3.N_1641\, Y => \I3.N_638_adt_net_134644_\);
    
    \I2.DT_TEMP_784\ : MUX2H
      port map(A => \I2.DT_TEMPl23r_net_1\, B => 
        \I2.DT_TEMP_7l23r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_784_net_1\);
    
    \I2.N_3822_adt_net_855588_\ : BFR
      port map(A => \I2.N_3822\, Y => 
        \I2.N_3822_adt_net_855588__net_1\);
    
    \I2.TDCDBSl11r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl11r, Q => 
        \I2.TDCDBSl11r_net_1\);
    
    \I3.VDBI_57_IV_0_0L7R_2227\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854356__net_1\, B
         => \I3.VDBoffl7r_net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_143093_\);
    
    \I2.N_4247_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4247\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4247_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2604\ : AND2
      port map(A => \REGl246r\, B => \I3.REGMAPl28r_net_1\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164420_\);
    
    \I2.CRC32l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_799_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l4r_net_1\);
    
    \I2.PIPE6_DT_480\ : MUX2H
      port map(A => \I2.PIPE5_DTl26r_net_1\, B => 
        \I2.PIPE6_DTl26r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_480_net_1\);
    
    \I2.OFFSET_37_8l2r\ : MUX2L
      port map(A => \REGl359r\, B => \REGl295r\, S => 
        \I2.PIPE7_DTL27R_72\, Y => \I2.N_693\);
    
    \I3.PIPEA_8l7r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854480__net_1\, B => 
        \I3.N_216\, Y => \I3.PIPEA_8l7r_net_1\);
    
    \I2.PIPE8_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_546_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl18r_net_1\);
    
    \I3.VAS_63\ : MUX2L
      port map(A => VAD_inl1r, B => \I3.VASl1r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_63_net_1\);
    
    \I2.PIPE4_DTl11r_1146\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL11R_408\);
    
    \I2.PIPE1_DT_42_1_IVL30R_1353\ : NAND2
      port map(A => \I2.N_3279_0_adt_net_855232__net_1\, B => 
        \I2.PIPE1_DT_42_1l29r\, Y => 
        \I2.PIPE1_DT_42l30r_adt_net_45594_\);
    
    \I3.N_1463_i_1_adt_net_855352_\ : BFR
      port map(A => \I3.N_1463_i_1\, Y => 
        \I3.N_1463_i_1_adt_net_855352__net_1\);
    
    \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__2831\ : OR3FFT
      port map(A => \I2.N_2870\, B => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854628__net_1\, 
        C => \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35789__net_1\, Y
         => \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\);
    
    \I1.BYTECNT_I_0_IL1R_2845\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_313_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.BYTECNT_I_0_IL1R_214\);
    
    \I5.SDAOUT_12_IV_0_921\ : OAI21FTT
      port map(A => \I5.COMMANDl2r_net_1\, B => \I5.N_70\, C => 
        \I5.N_150\, Y => \I5.SDAout_12_adt_net_9916_\);
    
    TDCDB_padl31r : IB33
      port map(PAD => TDCDB(31), Y => TDCDB_cl31r);
    
    \I2.TRGSERV_2_I_11\ : XOR2
      port map(A => \I2.TRGSERVl0r_net_1\, B => 
        \I2.STATE1_i_0_il15r\, Y => 
        \I2.DWACT_ADD_CI_0_partial_sum_1l0r\);
    
    \I2.EVNT_NUM_n10\ : NOR2
      port map(A => EV_RES_c, B => \I2.EVNT_NUM_n10_tz_i\, Y => 
        \I2.EVNT_NUM_n10_net_1\);
    
    \I2.DTO_1_886\ : MUX2L
      port map(A => \I2.DTO_1l12r_Rd1__net_1\, B => 
        \I2.DTO_16_1l12r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834768_Rd1__net_1\, Y
         => \I2.DTO_1l12r\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_A2_1_2674\ : OA21
      port map(A => \I2.N_140_0_ADT_NET_947__327\, B => 
        \I2.N_139_0_adt_net_55124_\, C => \I2.RAMDT4L12R_140\, Y
         => \I2.N_107_0_adt_net_320362_\);
    
    \I2.PIPE1_DT_42_1_ivl21r\ : OR3
      port map(A => \I2.PIPE1_DT_42l21r_adt_net_46861_\, B => 
        \I2.PIPE1_DT_42l21r_adt_net_46873_\, C => 
        \I2.PIPE1_DT_42l21r_adt_net_46874_\, Y => 
        \I2.PIPE1_DT_42l21r\);
    
    \I3.REGMAPl22r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un91_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl22r_net_1\);
    
    \I2.RAMDT4L5R_3062\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_816\);
    
    \I2.DT_TEMPl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_767_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl6r_net_1\);
    
    \I2.OFFSET_37_2l2r\ : MUX2L
      port map(A => \REGl383r\, B => \REGl319r\, S => 
        \I2.PIPE7_DTL27R_72\, Y => \I2.N_645\);
    
    \I3.PIPEA1_12l2r\ : AND2
      port map(A => DPR_cl2r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, Y => 
        \I3.PIPEA1_12l2r_net_1\);
    
    \I3.REGMAPL35R_2981\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un156_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL35R_528\);
    
    \I3.PULSE_46_0_iv_0_il2r\ : AO21
      port map(A => \I3.REGMAPl6r_net_1\, B => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        C => PULSEl2r, Y => \I3.N_122_adt_net_147352_\);
    
    \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__2907\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_320_adt_net_854876__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__361\);
    
    \I2.un1_DTE_1_sqmuxa_2_1_adt_net_4146_\ : NAND2
      port map(A => NOESRAME_C_242, B => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__181\, Y => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_4146__net_1\);
    
    \I1.PAGECNT_319_adt_net_854860_\ : BFR
      port map(A => \I1.PAGECNT_319_net_1\, Y => 
        \I1.PAGECNT_319_adt_net_854860__net_1\);
    
    \I2.SRAM_EVNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SRAM_EVNT_n1_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.SRAM_EVNTl1r_net_1\);
    
    \I2.REG_0l3r_adt_net_848__adt_net_854212_\ : BFR
      port map(A => \I2.REG_0l3r_adt_net_848__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\);
    
    \I2.CRC32l19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_814_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l19r_net_1\);
    
    \I2.PIPE1_DT_30l2r\ : MUX2L
      port map(A => \I2.TDCDBSl2r_net_1\, B => 
        \I2.TDCDBSl0r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, Y
         => \I2.PIPE1_DT_30l2r_net_1\);
    
    \I3.UN6_ASB_NE_2116\ : NOR2
      port map(A => \I3.N_262_i_0\, B => \I3.N_261_i_0\, Y => 
        \I3.un6_asb_NE_adt_net_135785_\);
    
    \I2.MIC_REG2L1R_2989\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_310_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2L1R_536\);
    
    \I2.FIDl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_433\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl17r);
    
    \I2.un1_STATE1_40_1_adt_net_45409_\ : OR3FTT
      port map(A => \I2.STATE1_1_sqmuxa_3\, B => 
        \I2.un1_STATE1_40_1_adt_net_45387__net_1\, C => 
        \I2.un1_STATE1_40_1_adt_net_45406__net_1\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45409__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I69_Y\ : AND2
      port map(A => \I2.N246_0\, B => \I2.N249_0\, Y => 
        \I2.N319_0\);
    
    \I3.PULSE_46_0_iv_i_il4r\ : AO21
      port map(A => \I3.REGMAPl10r_net_1\, B => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        C => \I3.N_55_adt_net_147183_\, Y => \I3.N_55\);
    
    \I1.PAGECNT_n7_i_i\ : OAI21
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_854524__net_1\, 
        B => \I1.N_403_i_i_0_i\, C => \I1.N_473\, Y => 
        \I1.N_1378\);
    
    \I2.CRC32_798\ : MUX2L
      port map(A => \I2.CRC32l3r_net_1\, B => \I2.N_3920\, S => 
        \I2.N_2826_1_adt_net_794__net_1\, Y => 
        \I2.CRC32_798_net_1\);
    
    \I2.N516_adt_net_87903_\ : AND3
      port map(A => \I2.N237_0\, B => 
        \I2.N411_adt_net_194931__net_1\, C => 
        \I2.N411_adt_net_194981__net_1\, Y => 
        \I2.N516_adt_net_87903__net_1\);
    
    \I2.OFFSET_37_3l3r\ : MUX2L
      port map(A => \I2.N_646\, B => \I2.N_638\, S => 
        \I2.PIPE7_DTL26R_349\, Y => \I2.N_654\);
    
    \I3.REG1_136\ : MUX2L
      port map(A => VDB_inl3r, B => \I3.REG1l3r_net_1\, S => 
        \I3.REG3_0_sqmuxa\, Y => \I3.REG1_136_net_1\);
    
    \I3.PIPEB_4l29r\ : NAND2FT
      port map(A => DPR_cl29r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855280__net_1\, 
        Y => \I3.PIPEB_4l29r_net_1\);
    
    \I3.VDBi_57_0_iv_0_a2_i_o3l19r\ : NAND2FT
      port map(A => \I3.N_1905_1\, B => 
        \I3.REGMAPl17r_adt_net_854300__net_1\, Y => \I3.N_1917\);
    
    \I3.UN1_NOEDTKI_0_SQMUXA_1_0_2315\ : OR2
      port map(A => \I3.STATE1_IPL8R_10\, B => 
        \I3.un1_NOEDTKi_0_sqmuxa_1_adt_net_159322_\, Y => 
        \I3.un1_NOEDTKi_0_sqmuxa_1_adt_net_159328_\);
    
    \I2.STATE5l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE5_ns_il1r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.STATE5l2r_net_1\);
    
    \I2.OFFSET_567\ : MUX2L
      port map(A => \I2.OFFSETl7r_net_1\, B => \I2.OFFSET_37l7r\, 
        S => \I2.UN1_NWPIPE7_2_297\, Y => \I2.OFFSET_567_net_1\);
    
    REGl379r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_280_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl379r\);
    
    \I2.STATE5l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE5_nsl3r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.STATE5l0r_net_1\);
    
    \I2.DTO_1l20r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l20r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l20r_Rd1__net_1\);
    
    \I2.UN1_STATE1_38_0_1531\ : AND3FFT
      port map(A => \I2.N_3287_i_0\, B => \I2.STATE1l10r_net_1\, 
        C => \I2.N_3283_adt_net_855064__net_1\, Y => 
        \I2.un1_STATE1_38_adt_net_52557_\);
    
    \I2.DTO_16_1_IV_1L1R_1209\ : NOR2
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620__net_1\, 
        B => \I2.DT_TEMPl1r_net_1\, Y => 
        \I2.DTO_16_1_iv_1l1r_adt_net_35122_\);
    
    \I3.PIPEA_8l3r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854460__net_1\, B => 
        \I3.N_212\, Y => \I3.PIPEA_8l3r_net_1\);
    
    \I3.REG_1l158r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_206_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl158r\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I138_Y_0_A2_1577\ : 
        NOR3FFT
      port map(A => \I2.N357\, B => \I2.N_53\, C => \I2.N_80\, Y
         => \I2.N_100_adt_net_58424_\);
    
    \I1.REG_74_0_ivl336r\ : AO21
      port map(A => \REGl336r\, B => \I1.N_209\, C => 
        \I1.REG_74l336r_adt_net_117572_\, Y => \I1.REG_74l336r\);
    
    \I1.REG_1_280\ : MUX2H
      port map(A => \REGl379r\, B => \I1.REG_74l379r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_280_net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2470\ : AO21
      port map(A => \REGl390r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l1r_adt_net_162928_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162935_\);
    
    \I2.REG_0L3R_ADT_NET_848__2766\ : AO21
      port map(A => \I3.REG1l3r_net_1\, B => \I3.REG2l3r_net_1\, 
        C => \I2.REG_0L3R_ADT_NET_19773_RD1__315\, Y => 
        \I2.REG_0L3R_ADT_NET_848__49\);
    
    \I1.REG_1_271\ : MUX2H
      port map(A => \REGl370r\, B => \I1.REG_74l370r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_271_net_1\);
    
    \I1.BYTECNTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_307_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTl7r_net_1\);
    
    \I3.UN15_ANYCYC_2296\ : AND3
      port map(A => \I3.PIPEAl28r_net_1\, B => 
        \I3.PIPEAl30r_net_1\, C => 
        \I3.un15_anycyc_adt_net_147616_\, Y => 
        \I3.un15_anycyc_adt_net_147611_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I47_Y\ : AND2
      port map(A => \I2.N279\, B => \I2.N282\, Y => \I2.N297_0\);
    
    \I1.REG_3_sqmuxa_0_a2_0_818\ : NAND2FT
      port map(A => \I1.PAGECNTL9R_244\, B => 
        \I1.N_238_Rd1__adt_net_854888__net_1\, Y => 
        \I1.N_254_196\);
    
    \I2.BNCID_VECTrff_15_250_0\ : AO21
      port map(A => \I2.BNCID_VECTwa15_1_net_1\, B => 
        \I2.BNCID_VECTrff_12_253_0_a2_0\, C => 
        \I2.BNCID_VECTro_15\, Y => 
        \I2.BNCID_VECTrff_15_250_0_net_1\);
    
    \I3.REG_1_152\ : MUX2L
      port map(A => VDB_inl3r, B => REGl51r, S => 
        \I3.N_1935_adt_net_855332__net_1\, Y => \I3.REG_1_152_0\);
    
    \I2.DTE_2_1l7r\ : XOR2
      port map(A => \I2.CRC32l3r_net_1\, B => 
        \I2.DTE_2_1_0l7r_net_1\, Y => \I2.DTE_2_1l7r_net_1\);
    
    \I1.REG_74_0_IVL309R_1907\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l309r_adt_net_119991_\);
    
    \I1.REG_74_0_IVL236R_1990\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_9_sqmuxa_adt_net_854724__net_1\, Y => 
        \I1.REG_74l236r_adt_net_127108_\);
    
    ADE_padl14r : OB33PH
      port map(PAD => ADE(14), A => ADE_cl14r);
    
    \I3.N_1905_1_adt_net_855380_\ : BFR
      port map(A => \I3.N_1905_1_adt_net_855384__net_1\, Y => 
        \I3.N_1905_1_adt_net_855380__net_1\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2519\ : AO21
      port map(A => \REGl227r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.N_2070_adt_net_163462_\, Y => 
        \I3.N_2070_adt_net_163500_\);
    
    REGl185r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_86_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl185r\);
    
    \I2.DT_TEMPl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_781_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl20r_net_1\);
    
    \I2.TDCDASl14r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl14r, Q => 
        \I2.TDCDASl14r_net_1\);
    
    FID_padl2r : OB33PH
      port map(PAD => FID(2), A => FID_cl2r);
    
    \I2.TDC_650\ : MUX2H
      port map(A => \I2.TDCl0r_net_1\, B => 
        \I2.RAMAD1_12l13r_net_1\, S => 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_1038__net_1\, Y => 
        \I2.TDC_650_net_1\);
    
    \I3.REG_1_156\ : MUX2L
      port map(A => VDB_inl7r, B => REGl55r, S => 
        \I3.N_1935_adt_net_855328__net_1\, Y => \I3.REG_1_156_0\);
    
    \I2.DTE_21_1_IV_0L5R_1327\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855192__net_1\, 
        B => \I2.DT_TEMPl5r_net_1\, C => 
        \I2.DTE_21_1l5r_adt_net_39083_\, Y => 
        \I2.DTE_21_1l5r_adt_net_39098_\);
    
    \I5.SBYTE_65\ : MUX2H
      port map(A => \I5.SBYTEl0r_net_1\, B => \I5.SBYTE_9l0r\, S
         => \I5.N_406\, Y => \I5.SBYTE_65_net_1\);
    
    \I1.REG_74_22l404r_811\ : OR3FFT
      port map(A => \I1.REG_74_4_i_a2_404_N_4_i\, B => 
        \I1.N_347_adt_net_854792__net_1\, C => \I1.N_396_192\, Y
         => \I1.N_201_9_189\);
    
    \I3.PIPEA_8_0l30r\ : MUX2L
      port map(A => DPR_cl30r, B => \I3.PIPEA1l30r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855356__net_1\, Y => \I3.N_239\);
    
    \I1.REG_74_0_IVL329R_1887\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l329r_adt_net_118174_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I153_Y_i_o3\ : AO21
      port map(A => \I2.PIPE4_DTL11R_410\, B => 
        \I2.PIPE4_DTL12R_512\, C => \I2.RAMDT4L5R_820\, Y => 
        \I2.N_20_i\);
    
    \I2.PIPE3_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl0r_net_1\);
    
    \I2.N_4547_1_adt_net_1209__adt_net_855608_\ : BFR
      port map(A => \I2.N_4547_1_adt_net_1209__net_1\, Y => 
        \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\);
    
    \I1.REG_74_0_ivl183r\ : AO21
      port map(A => \REGl183r\, B => \I1.N_57_269\, C => 
        \I1.REG_74l183r_adt_net_132043_\, Y => \I1.REG_74l183r\);
    
    \I2.ROFFSET_n2_tz\ : XOR2
      port map(A => \I2.ROFFSETl2r_net_1\, B => 
        \I2.ROFFSET_c1_net_1\, Y => \I2.ROFFSET_n2_tz_i\);
    
    \I3.VDBi_57_ivl1r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855384__net_1\, B => 
        \I3.VDBi_43l1r_net_1\, C => 
        \I3.VDBi_57l1r_adt_net_145947_\, Y => \I3.VDBi_57l1r\);
    
    \I3.VDBOFFB_30_IV_0L2R_2443\ : AND2
      port map(A => \REGl311r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        Y => \I3.VDBoffb_30l2r_adt_net_162714_\);
    
    \I2.L2TYPE_592\ : MUX2L
      port map(A => \I2.L2TYPEl3r_net_1\, B => \I2.N_4449\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_592_net_1\);
    
    \I2.RAMAD1_12l3r\ : MUX2L
      port map(A => \I2.TDCDASl1r_net_1\, B => 
        \I2.TDCDBSl1r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855176__net_1\, Y => 
        \I2.RAMAD1_12l3r_net_1\);
    
    \I2.STATE3l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3l1r_net_1\);
    
    RAMDT_padl11r : IOB33PH
      port map(PAD => RAMDT(11), A => \I1.RAMDT_SPI_1l4r_net_1\, 
        EN => \I1.RAMDT_SPI_E_0\, Y => RAMDT_inl11r);
    
    \I3.UN975_REGMAP_3_I_0_O2_I_A2_2085\ : NOR2
      port map(A => \I3.REGMAP_I_0_IL38R_113\, B => 
        \I3.REGMAPL39R_112\, Y => \I3.N_560_adt_net_134484_\);
    
    \I2.PIPE1_DT_42_1_IVL7R_1478\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl23r_net_1\, Y => 
        \I2.PIPE1_DT_42l7r_adt_net_50673_\);
    
    \I1.REG_8_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_268_Rd1__adt_net_854800__net_1\, B => 
        \I1.N_243_167\, Y => \I1.N_12233_i\);
    
    \I3.PIPEAl24r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_255_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl24r_net_1\);
    
    \I1.REG_1_283\ : MUX2H
      port map(A => \REGl382r\, B => \I1.REG_74l382r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_283_net_1\);
    
    \I2.FID_7_0_IVL11R_969\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl11r_net_1\, 
        Y => \I2.FID_7l11r_adt_net_18269_\);
    
    \I3.PIPEB_102\ : AO21
      port map(A => DPR_cl23r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\, 
        C => \I3.PIPEB_102_adt_net_159747_\, Y => 
        \I3.PIPEB_102_net_1\);
    
    \I2.DT_TEMP_787\ : MUX2H
      port map(A => \I2.DT_TEMPl26r_net_1\, B => 
        \I2.DT_TEMP_7l26r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_787_net_1\);
    
    \I2.EVNT_NUM_c1\ : AND2
      port map(A => \I2.EVNT_NUML0R_396\, B => 
        \I2.EVNT_NUML1R_397\, Y => \I2.EVNT_NUM_c1_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I179_Y_2685\ : AND3FFT
      port map(A => \I2.N303_0\, B => \I2.N357_1\, C => 
        \I2.N350_864\, Y => \I2.N481_adt_net_424213_\);
    
    \I1.SSTATE_NS_0_IV_0_0L1R_1771\ : AND3FTT
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.sstatel10r_net_1\, C => \I1.N_328_i_0\, Y => 
        \I1.sstate_nsl1r_adt_net_107663_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I95_Y\ : AO21FTT
      port map(A => \I2.N307_2\, B => \I2.N310_0\, C => 
        \I2.N306_i_i\, Y => \I2.N349\);
    
    \I1.PAGECNTe_adt_net_854892_\ : BFR
      port map(A => \I1.PAGECNTe\, Y => 
        \I1.PAGECNTe_adt_net_854892__net_1\);
    
    \I3.REG_1l94r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_275_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl94r\);
    
    \I2.PIPE8_DT_532\ : MUX2L
      port map(A => \I2.PIPE8_DTl4r_net_1\, B => 
        \I2.PIPE8_DT_21l4r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_532_net_1\);
    
    FID_padl25r : OB33PH
      port map(PAD => FID(25), A => FID_cl25r);
    
    \I2.PIPE1_DT_42_1_IVL7R_1482\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855228__net_1\, B => 
        \I2.MIC_ERR_REGSl7r_net_1\, C => 
        \I2.PIPE1_DT_42l7r_adt_net_50691_\, Y => 
        \I2.PIPE1_DT_42l7r_adt_net_50692_\);
    
    \I1.REG_74_0_IV_0L370R_1831\ : AND2
      port map(A => \FBOUTl5r\, B => \I1.N_593\, Y => 
        \I1.REG_74l370r_adt_net_113482_\);
    
    \I2.PIPE1_DT_42_1_IVL8R_1474\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl4r\, Y => 
        \I2.PIPE1_DT_42l8r_adt_net_50436_\);
    
    \I1.REG_1_171\ : MUX2H
      port map(A => \REGl270r\, B => \I1.REG_74l270r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y => 
        \I1.REG_1_171_net_1\);
    
    \I2.PIPE10_DT_608\ : MUX2L
      port map(A => \I2.PIPE10_DTl3r_net_1\, B => 
        \I2.PIPE9_DTl3r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_608_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I119_Y_I_O4_1585\ : 
        AOI21TTF
      port map(A => \I2.RAMDT4L12R_798\, B => 
        \I2.N_3_adt_net_940__net_1\, C => \I2.N_31_0\, Y => 
        \I2.N_3_0_adt_net_59703_\);
    
    \I3.PIPEA1_309\ : MUX2L
      port map(A => \I3.PIPEA1l11r_net_1\, B => 
        \I3.PIPEA1_12l11r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__253\, Y => 
        \I3.PIPEA1_309_net_1\);
    
    \I1.REG_74l300r\ : NAND2FT
      port map(A => \I1.REG_18_sqmuxa\, B => \I1.REG_74_1l308r\, 
        Y => \I1.N_169\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I154_Y_0_o2\ : OR2FT
      port map(A => \I2.N_8\, B => \I2.N_163_adt_net_1241__net_1\, 
        Y => \I2.N_82_adt_net_496796_\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I100_Y_1663\ : AND2
      port map(A => \I2.N310\, B => \I2.N306\, Y => 
        \I2.N466_adt_net_71184_\);
    
    \I2.UN1_REG80_I_1699\ : NOR2
      port map(A => REGL33R_389, B => REGL34R_563, Y => 
        \I2.N_3824_adt_net_90291_\);
    
    \I1.REG_74_0_IV_0_0L251R_1975\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l251r_adt_net_125691_\);
    
    \I3.REG_1l72r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_173_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl72r);
    
    NDTKIN_pad : OB33PH
      port map(PAD => NDTKIN, A => NDTKIN_c);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I180_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl10r_net_1\, Y => 
        \I2.ADD_21x21_fast_I180_Y_0\);
    
    \I1.LOAD_RESi_0\ : DFFC
      port map(CLK => CLK_c, D => \I1.LOAD_RESi_50_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => LOAD_RES_1);
    
    \I5.COMMAND_4l11r\ : MUX2L
      port map(A => \I5.AIR_WDATAl11r_net_1\, B => REGl112r, S
         => REGl7r, Y => \I5.COMMAND_4l11r_net_1\);
    
    \I1.REG_74_0_IVL311R_1905\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l311r_adt_net_119819_\);
    
    \I2.WOFFSET_13_il4r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_20\, Y => \I2.N_4247\);
    
    \I1.REG_74_8_0_o4_372_m7_i_x2\ : XOR2FT
      port map(A => \I1.N_299_adt_net_833868_Rd1__net_1\, B => 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__adt_net_855516__net_1\, 
        Y => \I1.REG_74_8_0_o4_372_N_9_i\);
    
    \I3.VDBoffa_49\ : OR3
      port map(A => \I3.VDBoffa_49_adt_net_163738_\, B => 
        \I3.VDBoffa_31l5r_adt_net_163699_\, C => 
        \I3.VDBoffa_31l5r_adt_net_163700_\, Y => 
        \I3.VDBoffa_49_net_1\);
    
    \I2.SUB8_517\ : MUX2H
      port map(A => \I2.SUB8l14r_adt_net_855568__net_1\, B => 
        \I2.SUB8_2l14r\, S => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855140__net_1\, Y => 
        \I2.SUB8_517_net_1\);
    
    \I2.resyn_0_I2_TRGCNT_c2_i\ : OAI21TTF
      port map(A => \I2.TRGCNTl2r_net_1\, B => \I2.N_3796\, C => 
        \I2.N_3763_adt_net_16097_\, Y => \I2.N_3763\);
    
    \I2.PIPE1_DT_42_1_IV_2L26R_1369\ : OAI21TTF
      port map(A => REGl446r, B => 
        \I2.N_3234_adt_net_855652__net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46173_\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46178_\);
    
    \I2.TDCGDAi_672\ : MUX2L
      port map(A => TDCGDA_c, B => \I2.un1_STATE1_23_net_1\, S
         => \I2.un1_STATE1_30_net_1\, Y => \I2.TDCGDAi_672_net_1\);
    
    \I0.EV_RESi\ : DFFC
      port map(CLK => CLK_c, D => \I0.EV_RESi_1_net_1\, CLR => 
        \I0.un4_hwresi_i\, Q => EV_RES_c);
    
    \I3.VDBi_57_0_iv_0l20r\ : OR2
      port map(A => \I3.VDBi_57l20r_adt_net_139290_\, B => 
        \I3.VDBi_57l20r_adt_net_139291_\, Y => \I3.VDBi_57l20r\);
    
    \I2.N_565_0_adt_net_855736_\ : BFR
      port map(A => \I2.N_565_0\, Y => 
        \I2.N_565_0_adt_net_855736__net_1\);
    
    \I3.un101_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_582\, B => \I3.N_551\, Y => 
        \I3.un101_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.ROFFSETl2r_1138\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_916_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETL2R_400\);
    
    REGl225r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_126_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl225r\);
    
    \I2.un21_sram_empty_3\ : XOR2
      port map(A => \I2.RPAGEL15R_522\, B => \I2.L2ARRL3R_605\, Y
         => \I2.un21_sram_empty_3_net_1\);
    
    REGl228r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_129_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl228r\);
    
    \I2.DTO_16_1_IV_0L27R_1081\ : AO21FTT
      port map(A => \I2.N_4647\, B => \I2.N_197\, C => 
        \I2.DTO_16_1l27r_adt_net_29242_\, Y => 
        \I2.DTO_16_1l27r_adt_net_29252_\);
    
    \I3.VADm_0_a3l17r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl17r_net_1\, Y => \I3.VADml17r\);
    
    \I3.REG_44_il87r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_1633_adt_net_150293_\, Y => \I3.N_1633\);
    
    VDB_padl20r : IOB33PH
      port map(PAD => VDB(20), A => \I3.VDBml20r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl20r);
    
    \I2.RAMAD1_655\ : MUX2L
      port map(A => \I2.RAMAD1_12l1r_net_1\, B => 
        \I2.RAMAD1l1r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__173\, Y => 
        \I2.RAMAD1_655_net_1\);
    
    \I2.PIPE7_DTL27R_2780\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_73\);
    
    \I1.REG_74_0_IVL178R_2056\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, Y => 
        \I1.REG_74l178r_adt_net_132510_\);
    
    \I1.REG_1_102\ : MUX2H
      port map(A => \REGl201r\, B => \I1.N_1340\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\, Y => 
        \I1.REG_1_102_net_1\);
    
    \I3.PIPEB_85\ : AO21
      port map(A => DPR_cl6r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_85_adt_net_160461_\, Y => 
        \I3.PIPEB_85_net_1\);
    
    \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_1_1_net_1\, Y => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\);
    
    \I2.G_EVNT_NUM_n9_0\ : AND2FT
      port map(A => EV_RES_C_569, B => 
        \I2.G_EVNT_NUM_n9_adt_net_26657_\, Y => 
        \I2.G_EVNT_NUM_n9\);
    
    \I2.PIPE1_DT_12l16r\ : MUX2L
      port map(A => \I2.TDCDASl16r_net_1\, B => 
        \I2.TDCDASl14r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, Y
         => \I2.PIPE1_DT_12l16r_net_1\);
    
    \I2.N_22_i_0_adt_net_855596_\ : BFR
      port map(A => \I2.N_22_i_0\, Y => 
        \I2.N_22_i_0_adt_net_855596__net_1\);
    
    \I1.REG_4_sqmuxa_0_a2_0_0_o2\ : NAND2
      port map(A => \I1.PAGECNT_321_net_1\, B => 
        \I1.PAGECNT_322_net_1\, Y => \I1.N_299_Ra1_\);
    
    \I3.VDBOFFB_30_IV_0L3R_2427\ : AO21
      port map(A => \REGl400r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l3r_adt_net_162504_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162548_\);
    
    \I2.PIPE1_DT_42_1_IVL7R_1483\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855756__net_1\, B => 
        \I2.PIPE1_DT_30l7r_net_1\, C => 
        \I2.PIPE1_DT_42l7r_adt_net_50677_\, Y => 
        \I2.PIPE1_DT_42l7r_adt_net_50693_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I180_UN1_Y_2659\ : NAND3FTT
      port map(A => \I2.N359_adt_net_86622_\, B => 
        \I2.N495_i_adt_net_202032_\, C => 
        \I2.N495_i_adt_net_202093_\, Y => 
        \I2.I180_un1_Y_adt_net_240115_\);
    
    \I2.DTE_21_1_IVL11R_1295\ : AND2FT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_289\, B => 
        \I2.DT_SRAMl11r_net_1\, Y => 
        \I2.DTE_21_1l11r_adt_net_38407_\);
    
    \I3.REGMAPl25r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un106_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl25r_net_1\);
    
    \I2.PIPE6_DT_467\ : MUX2H
      port map(A => \I2.PIPE5_DTl13r_net_1\, B => 
        \I2.PIPE6_DTl13r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_467_net_1\);
    
    \I2.OFFSET_37_18l1r\ : MUX2L
      port map(A => \REGl246r\, B => \REGl182r\, S => 
        \I2.PIPE7_DTL27R_85\, Y => \I2.N_772\);
    
    \I0.TDC_RESI_1_937\ : AND2FT
      port map(A => \I0.COM_SERF1_net_1\, B => COM_SERS, Y => 
        \I0.TDC_RESi_1_adt_net_15858_\);
    
    \I3.PIPEAl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_234_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl3r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I197_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl1r\, B => 
        \I2.PIPE7_DTl1r_net_1\, Y => \I2.SUB_21x21_fast_I197_Y_0\);
    
    \I1.RAMDT_SPI_1l0r\ : DFFC
      port map(CLK => CLK_c, D => \FBOUTl0r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.RAMDT_SPI_1l0r_net_1\);
    
    \I1.REG_74_0_ivl317r\ : AO21
      port map(A => \REGl317r\, B => \I1.N_193\, C => 
        \I1.REG_74l317r_adt_net_119303_\, Y => \I1.REG_74l317r\);
    
    REGl206r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_107_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl206r\);
    
    ADO_padl13r : OB33PH
      port map(PAD => ADO(13), A => ADO_cl13r);
    
    \I2.DTO_16_1l8r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l8r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l8r_Rd1__net_1\);
    
    \I1.REG_74_0_ivl279r\ : AO21
      port map(A => \REGl279r\, B => \I1.N_153\, C => 
        \I1.REG_74l279r_adt_net_122807_\, Y => \I1.REG_74l279r\);
    
    \I3.VDBOFFA_31_IV_0L1R_2614\ : AO21
      port map(A => \REGl182r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.VDBoffa_31l1r_adt_net_164448_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164455_\);
    
    \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108_\ : BFR
      port map(A => \I2.un3_tdcgda1_1_adt_net_821__net_1\, Y => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\);
    
    CLK_pad : GL33
      port map(PAD => CLK, GL => CLK_c);
    
    \I2.G_EVNT_NUM_n6_i_o2_0\ : AND2
      port map(A => \I2.N_4672_552\, B => 
        \I2.G_EVNT_NUMl6r_net_1\, Y => \I2.N_198\);
    
    \I3.un116_reg_ads_0_a2_2_a3\ : NOR2
      port map(A => \I3.N_584\, B => \I3.N_553\, Y => 
        \I3.un116_reg_ads_0_a2_2_a3_net_1\);
    
    \I3.REGMAPl9r_adt_net_854304_\ : BFR
      port map(A => \I3.REGMAPl9r_adt_net_854308__net_1\, Y => 
        \I3.REGMAPl9r_adt_net_854304__net_1\);
    
    \I1.SSTATE_NS_0_IV_0_0_O2L2R_1750\ : OR3FTT
      port map(A => \I1.BYTECNTL3R_434\, B => \I1.BYTECNTL2R_213\, 
        C => \I1.BYTECNT_I_0_IL1R_214\, Y => 
        \I1.N_321_adt_net_105403_\);
    
    \I3.PIPEAl5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_236_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl5r_net_1\);
    
    \I5.SBYTE_9_il5r\ : MUX2L
      port map(A => \I5.COMMANDl13r_net_1\, B => 
        \I5.SBYTEl4r_net_1\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.N_24\);
    
    \I2.PIPE1_DTl29r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_756_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl29r_net_1\);
    
    \I2.STATE3_0_SQMUXA_0_A7_1_1044\ : NOR2
      port map(A => \I2.DTESl31r_net_1\, B => \I2.DTESl29r_net_1\, 
        Y => \I2.STATE3_0_sqmuxa_1_0_adt_net_24559_\);
    
    \I2.MTDIAF1\ : DFFC
      port map(CLK => CLK_c, D => MTDIA_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.MTDIAF1_net_1\);
    
    \I2.BNCID_VECTrff_15\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_15_250_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_15\);
    
    \I1.REG_74_0_IVL387R_1806\ : AND2
      port map(A => \FBOUTl6r\, B => \I1.REG_28_sqmuxa\, Y => 
        \I1.REG_74l387r_adt_net_111405_\);
    
    \I1.N_161_adt_net_1449_\ : OR2
      port map(A => \I1.N_41_8\, B => 
        \I1.N_161_adt_net_121649__net_1\, Y => 
        \I1.N_161_adt_net_1449__net_1\);
    
    \I2.L2TYPE_593\ : MUX2L
      port map(A => \I2.L2TYPEl4r_net_1\, B => \I2.N_4448\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_593_net_1\);
    
    \I2.SUB9l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_569_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l1r_net_1\);
    
    \I2.FID_7_0_IVL15R_962\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl63r, C => 
        \I2.FID_7l15r_adt_net_17893_\, Y => 
        \I2.FID_7l15r_adt_net_17901_\);
    
    \I3.REGMAPl17r_adt_net_854296_\ : BFR
      port map(A => \I3.REGMAPl17r_adt_net_854300__net_1\, Y => 
        \I3.REGMAPl17r_adt_net_854296__net_1\);
    
    \I2.EVNT_NUM_n1\ : XOR2
      port map(A => \I2.N_1211\, B => \I2.N_1213\, Y => 
        \I2.EVNT_NUM_n1_net_1\);
    
    \I2.un2_evnt_word_I_51\ : AND2
      port map(A => \I2.WOFFSETl8r\, B => \I2.DWACT_FINC_E_0l4r\, 
        Y => \I2.N_19\);
    
    \I2.CRC32_1_sqmuxa_0_a2_0_a2_0_660\ : OR2
      port map(A => \I2.WR_SRAM_2_ADT_NET_748__39\, B => 
        \I2.N_4273\, Y => \I2.CRC32_1_SQMUXA_0_38\);
    
    \I2.ADEl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l15r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl15r);
    
    \I3.VDBOFFA_31_IV_0L0R_2631\ : AO21
      port map(A => \REGl245r\, B => \I3.REGMAPl28r_net_1\, C => 
        \I3.VDBoffa_31l0r_adt_net_164618_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164644_\);
    
    \I3.REGMAP_i_0_il36r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un161_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il36r_net_1\);
    
    \I2.PIPE5_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_676_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl0r_net_1\);
    
    \I2.un6_tdcgdb1_0\ : XOR2
      port map(A => \I2.TDCl0r_net_1\, B => \I2.TDCDBSl24r_net_1\, 
        Y => \I2.un6_tdcgdb1_0_net_1\);
    
    \I3.un96_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_585\, B => \I3.N_551\, Y => 
        \I3.un96_reg_ads_0_a2_0_a3_net_1\);
    
    \I1.REG_1_139\ : MUX2H
      port map(A => \REGl238r\, B => \I1.REG_74l238r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\, Y => 
        \I1.REG_1_139_net_1\);
    
    \I1.FCS\ : AND2
      port map(A => \I1.NCS0_net_1\, B => REGl82r, Y => FCS_c);
    
    \I3.VDBi_23_0_a2_1l1r\ : AND2FT
      port map(A => \I3.N_1907_266\, B => \I3.REGMAPL1R_725\, Y
         => \I3.N_2056\);
    
    \I2.DTE_1_841\ : MUX2L
      port map(A => \I2.DTE_1l1r_net_1\, B => 
        \I2.DTE_21_1_iv_i_0l1r\, S => \I2.N_2868_1\, Y => 
        \I2.DTE_1_841_net_1\);
    
    \I2.END_TDC1_1_sqmuxa_i_o3\ : OR2
      port map(A => \I2.TOKOUT_FL_net_1\, B => \I2.TOKOUTBS_163\, 
        Y => \I2.N_3879\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I175_Y\ : XOR2FT
      port map(A => \I2.N537_i_0\, B => 
        \I2.ADD_21x21_fast_I175_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l5r\);
    
    \I2.un1_tdc_res_42_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl412r, Y => 
        \I2.N_4623_i_0\);
    
    \I2.DTOSl30r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl30r, Q => 
        \I2.DTOSl30r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I38_Y\ : AND2
      port map(A => \I2.G_1\, B => \I2.N303_adt_net_69116_\, Y
         => \I2.N303\);
    
    \I2.STATE1_ns_0l11r\ : NAND3FFT
      port map(A => \I2.STATE1_nsl11r_adt_net_23387_\, B => 
        \I2.STATE1_nsl11r_adt_net_23385_\, C => 
        \I2.un1_STATE1_27\, Y => \I2.STATE1_nsl11r\);
    
    \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m2\ : XOR2
      port map(A => \I2.MIC_REG1_304_net_1\, B => 
        \I2.MIC_REG2_312_adt_net_855644__net_1\, Y => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Ra1_\);
    
    \I2.END_EVNT6_267\ : MUX2H
      port map(A => \I2.END_EVNT5_net_1\, B => 
        \I2.END_EVNT6_net_1\, S => END_FLUSH, Y => 
        \I2.END_EVNT6_267_net_1\);
    
    \I2.PIPE9_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_297_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl28r_net_1\);
    
    \I3.REGMAP_I_0_IL32R_3020\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un141_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL32R_774\);
    
    \I2.REG_0l3r_adt_net_19771_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.REG_0l3r_adt_net_19771_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.REG_0l3r_adt_net_19771_Rd1__net_1\);
    
    \I2.PIPE6_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_456_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl2r_net_1\);
    
    \I2.CHAIN_ERR_DIS\ : DFFC
      port map(CLK => CLK_c, D => \I2.CHAIN_ERR_DIS_448_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => REGl26r);
    
    \I2.BNCID_VECTrff_0_265_0_a2_0\ : NOR3FTT
      port map(A => TDCTRG_c, B => \I2.TRGARRl2r_net_1\, C => 
        \I2.TRGARRl3r_net_1\, Y => 
        \I2.BNCID_VECTrff_3_262_0_a2_0\);
    
    \I3.MBLTCYC_114\ : MUX2H
      port map(A => \I3.MBLTCYC_net_1\, B => 
        \I3.un7_cycs_0_a3_0_a3_net_1\, S => \I3.N_80\, Y => 
        \I3.MBLTCYC_114_net_1\);
    
    \I1.REG_74_12_300_M8_I_1908\ : AND2FT
      port map(A => \I1.N_1169_adt_net_854824__net_1\, B => 
        \I1.REG_74_12_300_N_15\, Y => 
        \I1.REG_74_12_300_N_11_adt_net_120111_\);
    
    \I1.REG_74_0_ivl181r\ : AO21
      port map(A => \REGl181r\, B => \I1.N_57\, C => 
        \I1.REG_74l181r_adt_net_132215_\, Y => \I1.REG_74l181r\);
    
    \I2.REG_1_n10\ : XOR2
      port map(A => \I2.N_3838\, B => \I2.REG_1_n10_0_net_1\, Y
         => \I2.REG_1_n10_net_1\);
    
    \I2.DTO_16_1_IV_0_0L19R_1124\ : AO21
      port map(A => \I2.G_EVNT_NUMl3r_net_1\, B => \I2.N_457\, C
         => \I2.DTO_16_1l19r_adt_net_30968_\, Y => 
        \I2.DTO_16_1l19r_adt_net_30979_\);
    
    \I3.VADm_0_a3l5r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl5r_net_1\, Y => \I3.VADml5r\);
    
    \I3.VDBI_57_IV_0L5R_2249\ : OAI21FTF
      port map(A => \FBOUTl5r\, B => \I3.N_2047\, C => 
        \I3.VDBi_57l5r_adt_net_143846_\, Y => 
        \I3.VDBi_57l5r_adt_net_143863_\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2202\ : AO21FTT
      port map(A => \I3.N_1905\, B => 
        \I3.VDBi_57l13r_adt_net_140454_\, C => 
        \I3.VDBi_57l13r_adt_net_140595_\, Y => 
        \I3.VDBi_57l13r_adt_net_140597_\);
    
    \I2.un2_evnt_word_I_30\ : AND2
      port map(A => \I2.WOFFSETl5r\, B => \I2.N_39\, Y => 
        \I2.N_34\);
    
    \I1.BYTECNT_308\ : MUX2H
      port map(A => \I1.BYTECNTl6r_net_1\, B => \I1.N_77\, S => 
        \I1.N_1383_225\, Y => \I1.BYTECNT_308_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2609\ : AO21
      port map(A => \REGl222r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.VDBoffa_31l1r_adt_net_164412_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164450_\);
    
    \I2.DT_TEMPl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_783_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl22r_net_1\);
    
    \I2.FID_7_0_IV_0L5R_1722\ : NOR2FT
      port map(A => \I2.STATE3l7r_net_1\, B => REGl53r, Y => 
        \I2.FID_7_0_iv_0l5r_adt_net_93017_\);
    
    \I2.DTE_21_1_IV_0L21R_1256\ : AO21
      port map(A => \I2.DT_SRAMl21r_net_1\, B => 
        \I2.N_199_0_ADT_NET_1054__37\, C => 
        \I2.DTE_21_1l21r_adt_net_37485_\, Y => 
        \I2.DTE_21_1l21r_adt_net_37496_\);
    
    \I1.REG_1_72\ : MUX2H
      port map(A => \REGl171r\, B => \I1.REG_74l171r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, Y => 
        \I1.REG_1_72_net_1\);
    
    \I2.PIPE5_DT_706\ : MUX2H
      port map(A => \I2.PIPE4_DTl30r_net_1\, B => 
        \I2.PIPE5_DTl30r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_706_net_1\);
    
    \I2.PIPE10_DT_17_i_o3l13r\ : NOR3FTT
      port map(A => \I2.PIPE9_DTL31R_667\, B => 
        \I2.PIPE9_DTL29R_669\, C => \I2.PIPE9_DTL30R_668\, Y => 
        \I2.N_22_i_0\);
    
    \I2.DTE_21_1_iv_0_0l7r\ : AO21
      port map(A => \I2.DTE_1l7r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, C => 
        \I2.DTE_21_1l7r_adt_net_38873_\, Y => \I2.DTE_21_1l7r\);
    
    \I2.N_3_0_adt_net_1070__adt_net_855604_\ : BFR
      port map(A => \I2.N_3_0_adt_net_1070__net_1\, Y => 
        \I2.N_3_0_adt_net_1070__adt_net_855604__net_1\);
    
    \I2.LSRAM_IN_409\ : MUX2L
      port map(A => \I2.PIPE5_DTl25r_net_1\, B => 
        \I2.LSRAM_INl25r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_409_net_1\);
    
    \I5.BITCNT_85\ : MUX2H
      port map(A => \I5.BITCNTl1r_net_1\, B => \I5.N_52\, S => 
        \I5.BITCNTe\, Y => \I5.BITCNT_85_net_1\);
    
    \I2.un1_STATE3_10_1_adt_net_17431_\ : NAND3FFT
      port map(A => \I2.STATE3L3R_415\, B => 
        \I2.STATE3_ns_il7r_net_1\, C => \I2.STATE3_il8r\, Y => 
        \I2.un1_STATE3_10_1_adt_net_17431__net_1\);
    
    \I2.PIPE1_DT_733\ : MUX2L
      port map(A => \I2.PIPE1_DTl6r_net_1\, B => 
        \I2.PIPE1_DT_42l6r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854584__net_1\, 
        Y => \I2.PIPE1_DT_733_net_1\);
    
    \I2.PIPE5_DT_6_0l2r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l2r\, B => 
        \I2.un27_pipe5_dt0l2r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1071\);
    
    \I1.REG_17_sqmuxa_adt_net_855480_\ : BFR
      port map(A => \I1.REG_17_sqmuxa\, Y => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\);
    
    \I2.PIPE7_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl2r_net_1\);
    
    \I2.resyn_0_I2_TRGCNT_n4\ : XOR2FT
      port map(A => \I2.N_3764\, B => \I2.TRGCNT_n4_0\, Y => 
        \I2.TRGCNT_n4\);
    
    REGl334r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_235_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl334r\);
    
    \I1.REG_74_0_iv_0_0l257r\ : AO21
      port map(A => \REGl257r\, B => \I1.N_658\, C => 
        \I1.REG_74l257r_adt_net_125056_\, Y => \I1.REG_74l257r\);
    
    \I1.BITCNT_n2_i_i_o2_647\ : AND2
      port map(A => \I1.BITCNTL0R_805\, B => \I1.BITCNTL1R_260\, 
        Y => \I1.N_324_25\);
    
    \I2.DTO_16_1_IV_1L3R_1204\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.DTO_9_ivl3r_net_1\, C => 
        \I2.DTO_16_1_iv_1l3r_adt_net_34602_\, Y => 
        \I2.DTO_16_1_iv_1l3r_adt_net_34608_\);
    
    \I3.N_57_i_0_0_adt_net_854700_\ : BFR
      port map(A => \I3.N_57_i_0_0\, Y => 
        \I3.N_57_i_0_0_adt_net_854700__net_1\);
    
    \I2.OFFSET_37_4l2r\ : MUX2L
      port map(A => \REGl367r\, B => \REGl303r\, S => 
        \I2.PIPE7_DTL27R_72\, Y => \I2.N_661\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I57_Y_0_o2\ : AO21
      port map(A => \I2.RAMDT4L8R_527\, B => 
        \I2.PIPE4_DT_I_IL1R_474\, C => \I2.N357_0_adt_net_55523_\, 
        Y => \I2.N357_0\);
    
    \I2.END_EVNT6\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT6_267_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.END_EVNT6_net_1\);
    
    VAD_padl8r : IOB33PH
      port map(PAD => VAD(8), A => \I3.VADml8r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl8r);
    
    \I5.TEMPDATAl0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_74_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl0r_net_1\);
    
    \I2.PIPE5_DT_704\ : MUX2L
      port map(A => \I2.PIPE5_DTl28r_net_1\, B => 
        \I2.PIPE5_DT_6l28r\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_704_net_1\);
    
    \I3.TCNT1_i_0_il1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT1_n1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT1_i_0_il1r_net_1\);
    
    \I2.LEAD_FLAG6l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_638_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl1r);
    
    \I1.REG_74_0_iv_i_a3l197r\ : OR2
      port map(A => \I1.N_181\, B => \I1.REG_6_sqmuxa\, Y => 
        \I1.N_182_i\);
    
    \I3.VADm_0_a3l30r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl30r_net_1\, Y => \I3.VADml30r\);
    
    \I3.PIPEA1l6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_304_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l6r_net_1\);
    
    \I2.REG_1l40r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n8_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl40r);
    
    \I2.BNCID_VECTrff_1_264_0\ : AO21
      port map(A => \I2.BNCID_VECTrff_3_262_0_a2_0\, B => 
        \I2.BNCID_VECTwa13_1_net_1\, C => \I2.BNCID_VECTro_1\, Y
         => \I2.BNCID_VECTrff_1_264_0_net_1\);
    
    REGl188r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_89_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl188r\);
    
    \I2.NWPIPE5\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE4_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE5_net_1\);
    
    \I2.SRAM_EVNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SRAM_EVNT_n0_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.SRAM_EVNTl0r_net_1\);
    
    \I1.REG_74_0_ivl214r\ : AO21
      port map(A => \REGl214r\, B => \I1.N_89\, C => 
        \I1.REG_74l214r_adt_net_129292_\, Y => \I1.REG_74l214r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I9_P0N_i_o3\ : OR2
      port map(A => \I2.RAMDT4L5R_821\, B => 
        \I2.PIPE4_DTl9r_net_1\, Y => \I2.N_13_0\);
    
    \I3.PIPEBl0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_79_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl0r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I189_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_799\, B => 
        \I2.PIPE4_DTl19r_net_1\, Y => 
        \I2.ADD_21x21_fast_I189_Y_0_0\);
    
    \I3.VDBOFFB_30_IV_0L6R_2371\ : AND2
      port map(A => \REGl363r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        Y => \I3.VDBoffb_30l6r_adt_net_161954_\);
    
    \I3.REG_1_271\ : MUX2H
      port map(A => REGl90r, B => \I3.N_1636\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_271_0\);
    
    \I2.PIPE5_DT_691\ : MUX2L
      port map(A => \I2.PIPE5_DTl15r_net_1\, B => 
        \I2.PIPE5_DT_6l15r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_691_net_1\);
    
    \I3.TCNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_384_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTl0r_net_1\);
    
    \I1.PAGECNT_n3_0_0_x2\ : XOR2
      port map(A => \I1.PAGECNTl3r_adt_net_835116_Rd1__net_1\, B
         => \I1.N_305_Rd1__net_1\, Y => \I1.N_393_i_i_0_i\);
    
    \I2.OFFSET_37_13l0r\ : MUX2L
      port map(A => \I2.N_723\, B => \I2.N_707\, S => 
        \I2.PIPE7_DTL25R_686\, Y => \I2.N_731\);
    
    \I2.DTO_16_1_iv_0_0l26r\ : OR2
      port map(A => \I2.DTO_16_1l26r_adt_net_29437_\, B => 
        \I2.DTO_16_1l26r_adt_net_29438_\, Y => \I2.DTO_16_1l26r\);
    
    \I2.PIPE9_DT_300\ : MUX2H
      port map(A => \I2.PIPE8_DTl31r_net_1\, B => 
        \I2.PIPE9_DTl31r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_300_net_1\);
    
    \I2.PHASE\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_c);
    
    \I2.END_CHAINB1_0_sqmuxa_i_a2_i_o3_0\ : OR2
      port map(A => REGl26r, B => \I2.N_3876\, Y => 
        \I2.CHAINB_EN244_c_0\);
    
    \I2.REG_1_n8\ : XOR2FT
      port map(A => \I2.N_3836_i_0\, B => \I2.REG_1_n8_0_net_1\, 
        Y => \I2.REG_1_n8_net_1\);
    
    \I1.REG_74_13_0_x2l404r\ : XOR2FT
      port map(A => \I1.PAGECNTl6r_adt_net_854924__net_1\, B => 
        \I1.PAGECNTl5r_net_1\, Y => \I1.N_330_i_0_i\);
    
    \I3.REG1_137\ : MUX2L
      port map(A => VDB_inl4r, B => \I3.REG1l4r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG1_137_net_1\);
    
    \I3.PIPEBl9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_88_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl9r_net_1\);
    
    \I3.N_48_I_0_O2_2088\ : NOR2
      port map(A => \I3.REGMAP_I_0_IL40R_450\, B => 
        \I3.REGMAPL37R_449\, Y => \I3.N_177_adt_net_134570_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I153_Y_i\ : NAND3
      port map(A => \I2.N_20_i\, B => \I2.N_33\, C => \I2.N_86_i\, 
        Y => \I2.N_2\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2514\ : AND2
      port map(A => \REGl251r\, B => \I3.REGMAPl28r_net_1\, Y => 
        \I3.N_2070_adt_net_163470_\);
    
    \I3.PIPEA_257\ : MUX2L
      port map(A => \I3.PIPEAl26r_net_1\, B => 
        \I3.PIPEA_8l26r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854656__net_1\, Y
         => \I3.PIPEA_257_net_1\);
    
    \I2.DTO_16_1_IV_0L24R_1094\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854612__net_1\, 
        B => \I2.DT_TEMPl24r_net_1\, C => 
        \I2.DTO_16_1l24r_adt_net_29860_\, Y => 
        \I2.DTO_16_1l24r_adt_net_29868_\);
    
    \I3.PIPEB_109\ : MUX2H
      port map(A => \I3.PIPEBl30r_net_1\, B => 
        \I3.PIPEB_4l30r_net_1\, S => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_109_net_1\);
    
    \I1.BYTECNTlde_i_a2_i_846\ : AO21
      port map(A => \I1.N_628\, B => 
        \I1.sstate_ns_i_0_a4_0_1l0r_adt_net_107171_\, C => 
        \I1.N_223_226\, Y => \I1.N_1383_224\);
    
    \I2.DTO_16_1_iv_0_0l29r\ : OR2
      port map(A => \I2.DTO_16_1l29r_adt_net_28739_\, B => 
        \I2.DTO_16_1l29r_adt_net_28740_\, Y => \I2.DTO_16_1l29r\);
    
    \I1.REG_74_0_ivl229r\ : AO21
      port map(A => \REGl229r\, B => \I1.N_105\, C => 
        \I1.REG_74l229r_adt_net_127710_\, Y => \I1.REG_74l229r\);
    
    \I3.VDBoffb_30_iv_0l3r\ : AND2
      port map(A => \REGl368r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162504_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_A2_1_2675\ : 
        OR3FFT
      port map(A => \I2.N_28_0\, B => \I2.N_108_0_adt_net_55153_\, 
        C => \I2.N_107_0_adt_net_320362_\, Y => \I2.N_107_0\);
    
    \I2.TRGSERV_2_I_19\ : AND2
      port map(A => \I2.DWACT_ADD_CI_0_TMP_0l0r\, B => 
        \I2.TRGSERVl1r_net_1\, Y => 
        \I2.DWACT_ADD_CI_0_g_array_1_0l0r\);
    
    \I3.PIPEBl25r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_104_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl25r_net_1\);
    
    \I2.OFFSET_37_28l1r\ : MUX2L
      port map(A => \I2.N_844\, B => \I2.N_796\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_852\);
    
    \I3.VDBi_23_0_a2l1r\ : OR2
      port map(A => \I3.N_2018\, B => \I3.REGMAPl3r_net_1\, Y => 
        \I3.N_2031\);
    
    \I1.REG_74_0_IV_I_A2L208R_2026\ : AND2
      port map(A => \REGl208r\, B => \I1.N_183_i_0\, Y => 
        \I1.N_1347_adt_net_129845_\);
    
    \I3.VDBil22r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_362_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil22r_net_1\);
    
    \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854908_\ : BFR
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__831\, Y => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854908__net_1\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854472_\ : BFR
      port map(A => \I3.N_243_4_adt_net_1290__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854472__net_1\);
    
    \I2.LSRAM_RADDRil1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_RADDRi_500\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.LSRAM_RADDRil1r_net_1\);
    
    \I2.SRAM_EVNT_n3\ : XOR2
      port map(A => \I2.N_3827\, B => \I2.SRAM_EVNT_n3_0_net_1\, 
        Y => \I2.SRAM_EVNT_n3_net_1\);
    
    EV_RES_pad : OB33PH
      port map(PAD => EV_RES, A => EV_RES_C_569);
    
    \I2.PIPE6_DT_479\ : MUX2H
      port map(A => \I2.PIPE5_DTl25r_net_1\, B => 
        \I2.PIPE6_DTl25r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_479_net_1\);
    
    \I2.resyn_0_I2_FID_442\ : MUX2H
      port map(A => FID_cl26r, B => \I2.FID_7l26r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\, 
        Y => \I2.FID_442\);
    
    \I5.REG_1_39\ : MUX2L
      port map(A => \I5.TEMPDATAl6r_net_1\, B => REGl426r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_39_net_1\);
    
    \I2.DTE_21_1_IV_0L10R_1299\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855116__net_1\, B => 
        \I2.EVNT_WORDl6r_net_1\, Y => 
        \I2.DTE_21_1l10r_adt_net_38511_\);
    
    \I2.UN1_STATE3_12_I_1712\ : OR3
      port map(A => \I2.STATE3_nsl6r_adt_net_24857_\, B => 
        \I2.N_2989_adt_net_92422_\, C => \I2.STATE3l11r_net_1\, Y
         => \I2.N_2989_adt_net_92425_\);
    
    \I2.RAMAD1l14r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_668_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l14r_net_1\);
    
    REGl374r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_275_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl374r\);
    
    \I1.SBYTE_63\ : MUX2L
      port map(A => \FBOUTl5r\, B => \I1.N_204\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_63_net_1\);
    
    \I3.VDBi_57l8r_adt_net_142588_\ : AND2
      port map(A => REGl414r, B => \I3.REGMAPl55r_net_1\, Y => 
        \I3.VDBi_57l8r_adt_net_142588__net_1\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__2972\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__489\);
    
    \I1.REG_74_12_348_M9_I_1854\ : AND2
      port map(A => \I1.REG_74_2_4_il228r\, B => 
        \I1.REG_74_12_348_m9_i_adt_net_115329_\, Y => 
        \I1.REG_74_12_348_m9_i_adt_net_115422_\);
    
    \I2.DTO_1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_879_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l5r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I152_Y_0_a2\ : OA21
      port map(A => \I2.N_147_0_adt_net_604875_\, B => 
        \I2.N_82_adt_net_496796_\, C => \I2.N_33_adt_net_55021_\, 
        Y => \I2.N_103\);
    
    \I2.STATE1_ns_i_o2l9r\ : OR3
      port map(A => FLUSH, B => \I2.FCNT_c1\, C => 
        \I2.FCNTL2R_600\, Y => \I2.N_3272\);
    
    \I2.RAMDT4L5R_3060\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_814\);
    
    \I3.un1_STATE2_9\ : OAI21FTF
      port map(A => \I3.STATE2l1r_net_1\, B => \I3.N_1861\, C => 
        \I3.un1_STATE2_9_adt_net_154004_\, Y => 
        \I3.un1_STATE2_9_net_1\);
    
    \I5.un1_SENS_ADDR_1_I_9\ : XOR2FT
      port map(A => \I5.SENS_ADDRl0r_net_1\, B => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\, Y
         => \I5.DWACT_ADD_CI_0_partial_suml0r\);
    
    \I1.REG_1_152\ : MUX2H
      port map(A => \REGl251r\, B => \I1.REG_74l251r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_152_net_1\);
    
    \I2.DTE_21_1_IV_0_0L4R_1333\ : AO21
      port map(A => \I2.DT_TEMPl4r_net_1\, B => \I2.N_4038\, C
         => \I2.DTE_21_1l4r_adt_net_39195_\, Y => 
        \I2.DTE_21_1l4r_adt_net_39209_\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854436_\ : BFR
      port map(A => \I2.N_4667_1_adt_net_1046__net_1\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854436__net_1\);
    
    \I3.N_1910_0_adt_net_854344_\ : BFR
      port map(A => \I3.N_1910_0_adt_net_854348__net_1\, Y => 
        \I3.N_1910_0_adt_net_854344__net_1\);
    
    \I2.PIPE6_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_475_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl21r_net_1\);
    
    \I3.VADm_0_a3l15r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl15r_net_1\, Y => \I3.VADml15r\);
    
    \I2.LSRAM_INl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_405_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl21r_net_1\);
    
    \I2.DTO_1l10r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l10r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l10r_Rd1__net_1\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854440_\ : BFR
      port map(A => \I2.N_4667_1_adt_net_1046__net_1\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854440__net_1\);
    
    \I5.AIR_WDATAl10r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_60_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl10r_net_1\);
    
    \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855076_\ : BFR
      port map(A => \I2.un2_tdcgdb1_0_adt_net_830__net_1\, Y => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855076__net_1\);
    
    DTO_padl29r : IOB33PH
      port map(PAD => DTO(29), A => \I2.DTO_1l29r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl29r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I51_Y\ : AND2
      port map(A => \I2.N273\, B => \I2.N276\, Y => \I2.N301_2\);
    
    \I1.REG_74l188r\ : OR2
      port map(A => \I1.REG_4_sqmuxa\, B => 
        \I1.N_65_ADT_NET_1433__217\, Y => \I1.N_57\);
    
    \I2.RAMDT4L12R_3074\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_828\);
    
    \I2.TDCDBSl20r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl20r, Q => 
        \I2.TDCDBSl20r_net_1\);
    
    \I2.DTE_21_1_IVL14R_1278\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855128__net_1\, B => 
        \I2.EVNT_WORDl10r_net_1\, Y => 
        \I2.DTE_21_1l14r_adt_net_38053_\);
    
    \I3.VDBOFFA_31_IV_0L5R_2536\ : AO21
      port map(A => \REGl226r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.VDBoffa_31l5r_adt_net_163648_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163689_\);
    
    \I3.VDBOFFA_31_IV_0L4R_2556\ : AO21
      port map(A => \REGl209r\, B => 
        \I3.REGMAPl23r_adt_net_855012__net_1\, C => 
        \I3.VDBoffa_31l4r_adt_net_163846_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163881_\);
    
    \I2.DTO_16_1_iv_0_a2_2l21r_675\ : AND3
      port map(A => \I2.N_223_54\, B => \I2.N_4182\, C => 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_888__net_1\, Y => 
        \I2.N_196_53\);
    
    \I3.N_1764_adt_net_854352_\ : BFR
      port map(A => \I3.N_1764\, Y => 
        \I3.N_1764_adt_net_854352__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I153_Y_0\ : XOR2FT
      port map(A => \I2.N_3560_i_net_1\, B => 
        \I2.N_3558_i_adt_net_855584__net_1\, Y => 
        \I2.ADD_18x18_fast_I153_Y_0\);
    
    \I2.SUB9_1_ADD_18x18_fast_I58_Y\ : AO21
      port map(A => \I2.N292\, B => \I2.N295\, C => \I2.N291\, Y
         => \I2.N326\);
    
    \I1.REG_74_0_IV_0L194R_2040\ : AND2
      port map(A => \REGl194r\, B => \I1.N_65_92\, Y => 
        \I1.REG_74l194r_adt_net_131097_\);
    
    \I3.un1_STATE1_13_1_adt_net_137890_\ : AND2FT
      port map(A => \I3.N_1905_1_adt_net_855376__net_1\, B => 
        \I3.N_638_117\, Y => 
        \I3.un1_STATE1_13_1_adt_net_137890__net_1\);
    
    \I2.DTO_1l31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_905_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l31r_net_1\);
    
    \I3.PIPEA_241\ : MUX2L
      port map(A => \I3.PIPEAl10r_net_1\, B => 
        \I3.PIPEA_8l10r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854672__net_1\, Y
         => \I3.PIPEA_241_net_1\);
    
    \I2.PIPE8_DT_16_sn_m1_0_a2_0\ : OR2FT
      port map(A => \I2.PIPE7_DTl31r_net_1\, B => 
        \I2.PIPE7_DTl30r_adt_net_855172__net_1\, Y => 
        \I2.N_565_0\);
    
    \I2.FID_7_0_IVL19R_954\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl67r, C => 
        \I2.FID_7l19r_adt_net_17517_\, Y => 
        \I2.FID_7l19r_adt_net_17525_\);
    
    \I2.PIPE7_DTL27R_2787\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_80\);
    
    \I3.TCNTlde_0_a2\ : NOR3FTT
      port map(A => \I3.WRITES_8\, B => \I3.N_1641\, C => 
        \I3.N_276\, Y => \I3.un1_STATE1_10_i_0\);
    
    \I2.PIPE1_DT_42_1_ivl4r\ : OR3
      port map(A => \I2.PIPE1_DT_42l4r_adt_net_51424_\, B => 
        \I2.PIPE1_DT_42l4r_adt_net_51433_\, C => 
        \I2.PIPE1_DT_42l4r_adt_net_51434_\, Y => 
        \I2.PIPE1_DT_42l4r\);
    
    \I3.VDBI_57_0_IV_0L21R_2165\ : AO21
      port map(A => REGl69r, B => \I3.N_1839\, C => 
        \I3.VDBi_57l21r_adt_net_139183_\, Y => 
        \I3.VDBi_57l21r_adt_net_139188_\);
    
    \I2.DTE_21_1_IV_2L1R_1343\ : OAI21TTF
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_290\, B => 
        \I2.DT_SRAMl1r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39592_\, Y => 
        \I2.DTE_21_1_iv_2_il1r_adt_net_39593_\);
    
    REGl286r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_187_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl286r\);
    
    \I3.STATE1_TR24_I_0_O2_1_0_2111\ : NAND2FT
      port map(A => \I3.N_276\, B => \I3.WRITES_8\, Y => 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135386_\);
    
    \I5.SBYTEl1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_66_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl1r_net_1\);
    
    \I1.REG_74_0_IVL226R_2001\ : AND2
      port map(A => \FBOUTl5r\, B => \I1.N_12233_i\, Y => 
        \I1.REG_74l226r_adt_net_128136_\);
    
    \I1.REG_1_221\ : MUX2H
      port map(A => \REGl320r\, B => \I1.REG_74l320r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_221_net_1\);
    
    \I2.un2_evnt_word_I_31\ : XOR2
      port map(A => \I2.WOFFSETl6r\, B => \I2.N_34\, Y => 
        \I2.I_31\);
    
    NOE16R_pad : OB33PH
      port map(PAD => NOE16R, A => NOE16R_c);
    
    \I2.RAMAD1_663\ : MUX2L
      port map(A => \I2.RAMAD1_12l9r_net_1\, B => 
        \I2.RAMAD1l9r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__171\, Y => 
        \I2.RAMAD1_663_net_1\);
    
    \I2.ADE_4l10r\ : MUX2H
      port map(A => \I2.WOFFSETl11r\, B => \I2.ROFFSETl11r_net_1\, 
        S => NOESRAME_c, Y => \I2.ADE_4l10r_net_1\);
    
    \I2.MIC_ERR_REGSl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_336_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl7r_net_1\);
    
    \I2.DTE_1l12r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l12r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l12r_Rd1__net_1\);
    
    \I2.BNCID_VECTrff_1\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_1_264_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_1\);
    
    \I3.TCNT2_393\ : MUX2H
      port map(A => \I3.TCNT2l3r_net_1\, B => \I3.TCNT2_n3_net_1\, 
        S => TICKl0r, Y => \I3.TCNT2_393_net_1\);
    
    \I2.PIPE1_DTl31r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_758_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl31r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I120_Y_0_o2_0_730\ : NAND2
      port map(A => \I2.N_64_0\, B => \I2.N_89_0_111\, Y => 
        \I2.N_72_0_108\);
    
    \I2.PIPE5_DT_6_0l14r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l14r\, B => 
        \I2.un27_pipe5_dt0l14r\, S => 
        \I2.dataout_0_adt_net_855804__net_1\, Y => \I2.N_1083\);
    
    \I3.PIPEBl17r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_96_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl17r_net_1\);
    
    \I2.N_2868_1_adt_net_835996_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2868_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\);
    
    \I2.resyn_0_I2_BITCNTlde_0\ : OR2
      port map(A => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855860__net_1\, B => 
        \I2.ERR_WORDS_RDY_0_sqmuxa\, Y => \I2.BITCNTe\);
    
    \I2.majority_reg_il0r\ : AO21
      port map(A => \I2.MIC_REG3l0r_net_1\, B => 
        \I2.MIC_REG2l0r_net_1\, C => \reg_il0r_adt_net_105174_\, 
        Y => reg_il0r);
    
    \I1.REG_74_0_iv_i_a2l212r\ : AO21
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, C => 
        \I1.N_1350_adt_net_129501_\, Y => \I1.N_1350\);
    
    \I2.CRC32_12_i_x2l14r\ : XOR2FT
      port map(A => \I2.CRC32l14r_net_1\, B => \I2.N_3959_i_i\, Y
         => \I2.N_4026_i_0\);
    
    \I2.CRC32_822\ : MUX2L
      port map(A => \I2.CRC32l27r_net_1\, B => \I2.N_3944\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_822_net_1\);
    
    \I2.N_587_adt_net_1201__adt_net_855164_\ : BFR
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\, Y => 
        \I2.N_587_adt_net_1201__adt_net_855164__net_1\);
    
    \I1.REG_74_0_IVL172R_2062\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l172r_adt_net_133063_\);
    
    \I3.VDBoffb_59\ : OR3
      port map(A => \I3.VDBoffb_59_adt_net_161840_\, B => 
        \I3.VDBoffb_30l7r_adt_net_161799_\, C => 
        \I3.VDBoffb_30l7r_adt_net_161800_\, Y => 
        \I3.VDBoffb_59_net_1\);
    
    \I2.resyn_0_I2_BITCNT_n2_i_o3\ : AND2
      port map(A => \I2.N_4327\, B => \I2.BITCNTl2r_net_1\, Y => 
        \I2.N_4328\);
    
    \I2.FID_7_0_ivl11r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl11r_net_1\, 
        C => \I2.FID_7l11r_adt_net_18277_\, Y => \I2.FID_7l11r\);
    
    \I2.RAMAD1_659\ : MUX2L
      port map(A => \I2.RAMAD1_12l5r_net_1\, B => 
        \I2.RAMAD1l5r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__172\, Y => 
        \I2.RAMAD1_659_net_1\);
    
    \I2.L1AF1\ : DFFC
      port map(CLK => CLK_c, D => L1A_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L1AF1_net_1\);
    
    \I2.PIPE7_DTL26R_2899\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_353\);
    
    \I3.PIPEA1_12l14r\ : AND2
      port map(A => DPR_cl14r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854500__net_1\, Y => 
        \I3.PIPEA1_12l14r_net_1\);
    
    FID_padl22r : OB33PH
      port map(PAD => FID(22), A => FID_cl22r);
    
    \I3.VDBOFFB_30_IV_0L7R_2364\ : OR3
      port map(A => \I3.VDBoffb_30l7r_adt_net_161795_\, B => 
        \I3.VDBoffb_30l7r_adt_net_161789_\, C => 
        \I3.VDBoffb_30l7r_adt_net_161790_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161799_\);
    
    \I2.L2SERVl3r_1257\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_519\);
    
    \I2.PIPE10_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_621_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl16r_net_1\);
    
    \I2.DTO_16_1_IV_0L31R_1066\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855680__net_1\, B => 
        \I2.DTO_9l31r\, C => \I2.DTO_16_1l31r_adt_net_28248_\, Y
         => \I2.DTO_16_1l31r_adt_net_28255_\);
    
    \I2.UN1_STATE2_7_0_1534\ : AND3FTT
      port map(A => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_N_20_i\, B
         => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_net_1\, C => 
        \I2.STATE2l2r_adt_net_855212__net_1\, Y => 
        \I2.un1_STATE2_7_adt_net_53240_\);
    
    \I1.REG_9_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_240\, B => \I1.N_255\, Y => 
        \I1.REG_9_sqmuxa\);
    
    \I3.CLOSEDTK\ : DFFC
      port map(CLK => \I3.N_95\, D => \VCC\, CLR => NOEDTK_c, Q
         => \I3.CLOSEDTK_net_1\);
    
    \I2.FID_7_0_IVL22R_991\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl22r_net_1\, 
        Y => \I2.FID_7l22r_adt_net_19303_\);
    
    \I1.REG_74_0_IV_I_A2L204R_2030\ : AND2
      port map(A => \REGl204r\, B => \I1.N_182_i\, Y => 
        \I1.N_1343_adt_net_130189_\);
    
    \I2.un6_tdcgdb1_2\ : XOR2
      port map(A => \I2.TDCl2r_net_1\, B => \I2.TDCDBSl26r_net_1\, 
        Y => \I2.un6_tdcgdb1_2_net_1\);
    
    \I2.RAMDT4l1r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl1r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l1r_net_1\);
    
    REGl396r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_297_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl396r\);
    
    \I2.PIPE4_DTl17r_1529\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl17r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL17R_636\);
    
    \I2.un1_STATE1_40_1_adt_net_45381_\ : NOR2
      port map(A => \I2.TDCGDB1_net_1\, B => \I2.N_3889\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45381__net_1\);
    
    \I2.DTE_1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_845_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l5r_net_1\);
    
    \I2.RAMAD_4l0r\ : MUX2L
      port map(A => \I2.N_527\, B => \I1.BYTECNTl0r_net_1\, S => 
        LOAD_RES, Y => \I2.RAMAD_4l0r_net_1\);
    
    \I5.REG_1_40\ : MUX2L
      port map(A => \I5.TEMPDATAl7r_net_1\, B => REGl427r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_40_net_1\);
    
    \I2.OFFSET_37_23l0r\ : MUX2L
      port map(A => \REGl269r\, B => \REGl205r\, S => 
        \I2.PIPE7_DTl27r_net_1\, Y => \I2.N_811\);
    
    \I3.RAMAD_VMEl11r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_35_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl11r);
    
    \I3.REG_1_179\ : MUX2L
      port map(A => VDB_inl30r, B => REGl78r, S => 
        \I3.N_1935_adt_net_855316__net_1\, Y => \I3.REG_1_179_0\);
    
    \I2.PIPE3_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl13r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl13r_net_1\);
    
    \I2.DTO_9_IVL24R_1090\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        B => \I2.G_EVNT_NUMl8r_net_1\, Y => 
        \I2.DTO_9l24r_adt_net_29794_\);
    
    \I3.un1_REGMAP_30_0_a2\ : AND3
      port map(A => \I3.un1_REGMAP_30_adt_net_134454_\, B => 
        \I3.un1_REGMAP_30_0_a2_0_net_1\, C => \I3.N_68\, Y => 
        \I3.un1_REGMAP_30\);
    
    \I2.ROFFSET_917\ : MUX2H
      port map(A => \I2.ROFFSETl1r_net_1\, B => 
        \I2.ROFFSET_n1_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_917_net_1\);
    
    \I2.PIPE8_DT_16_0l9r\ : MUX2H
      port map(A => \I2.PIPE8_DTl9r_net_1\, B => 
        \I2.PIPE7_DTl9r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_575\);
    
    \I2.N_199_0_adt_net_1054_\ : OAI21FTT
      port map(A => \I2.STATE2L3R_440\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.DTE_CL_0_SQMUXA_2_0_288\, Y => 
        \I2.N_199_0_adt_net_1054__net_1\);
    
    \I2.RAMADl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l16r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl16r);
    
    \I2.STATEe_1281\ : OR2
      port map(A => \I2.N_3496_adt_net_926__net_1\, B => 
        \I2.STATEel4r_net_1\, Y => \I2.N_3450\);
    
    \I2.FID_7_0_IVL8R_1716\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl8r_net_1\, 
        Y => \I2.FID_7l8r_adt_net_92739_\);
    
    \I2.CRC32l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_796_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l1r_net_1\);
    
    \I1.REG_1_121\ : MUX2H
      port map(A => \REGl220r\, B => \I1.REG_74l220r_net_1\, S
         => \I1.N_50_0_ADT_NET_1409__320\, Y => 
        \I1.REG_1_121_net_1\);
    
    \I2.CRC32_12_i_m2l14r\ : MUX2H
      port map(A => \I2.DT_SRAMl14r_net_1\, B => 
        \I2.DT_TEMPl14r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854432__net_1\, Y => 
        \I2.N_3959_i_i\);
    
    \I1.REG_1_282\ : MUX2H
      port map(A => \REGl381r\, B => \I1.REG_74l381r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_282_net_1\);
    
    \I3.REG_1_ml78r\ : AND2
      port map(A => REGl78r, B => 
        \I3.REGMAPl9r_adt_net_854304__net_1\, Y => 
        \I3.VDBi_20l30r\);
    
    \I3.REG1l7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG1_140_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l7r_net_1\);
    
    \I2.PIPE5_DT_6_0l10r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l10r\, B => 
        \I2.un27_pipe5_dt0l10r\, S => 
        \I2.dataout_0_adt_net_855804__net_1\, Y => \I2.N_1079\);
    
    \I2.EVNT_NUMl4r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_959_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl4r_net_1\);
    
    \I2.ADOl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l15r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl15r);
    
    \I3.VDBi_57_0_iv_2_0_m2l9r\ : MUX2H
      port map(A => \I3.VDBil9r_net_1\, B => \I3.RAMDTSl9r_net_1\, 
        S => \I3.N_57_i_0_0_adt_net_854696__net_1\, Y => 
        \I3.N_92\);
    
    \I2.MIC_ERR_REGS_336\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl8r_net_1\, B => 
        \I2.MIC_ERR_REGSl7r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_336_net_1\);
    
    REGl355r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_256_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl355r\);
    
    \I5.DATA_12l12r\ : MUX2L
      port map(A => REGl129r, B => \I5.SBYTEl4r_net_1\, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l12r_net_1\);
    
    \I5.COMMAND_12\ : MUX2H
      port map(A => \I5.COMMANDl0r_net_1\, B => 
        \I5.COMMAND_4l0r_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.COMMAND_12_net_1\);
    
    \I2.REG_1_C9_I_1740\ : AND2FT
      port map(A => REGl41r, B => \I2.N_129\, Y => 
        \I2.N_3838_adt_net_101306_\);
    
    \I2.RAMAD1l10r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_664_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l10r_net_1\);
    
    INTR2_pad : OB33PH
      port map(PAD => INTR2, A => \GND\);
    
    \I2.PIPE6_DT_459\ : MUX2H
      port map(A => \I2.PIPE5_DTl5r_net_1\, B => 
        \I2.PIPE6_DTl5r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_459_net_1\);
    
    \I2.DT_TEMPl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_777_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl16r_net_1\);
    
    \I2.PIPE10_DT_17_I_A3_2L13R_1612\ : OR3
      port map(A => \I2.N_3822_adt_net_64761_\, B => 
        \I2.SUB9_i_0_il17r\, C => \I2.SUB9l16r_net_1\, Y => 
        \I2.N_3822_adt_net_64765_\);
    
    \I2.DTE_21_1_IVL23R_1250\ : AO21FTT
      port map(A => \I2.DTE_cl_0_sqmuxa_2_0\, B => 
        \I2.DT_SRAMl23r_net_1\, C => 
        \I2.DTE_21_1l23r_adt_net_37283_\, Y => 
        \I2.DTE_21_1l23r_adt_net_37284_\);
    
    \I3.PIPEB_91_2332\ : NOR2FT
      port map(A => \I3.PIPEBl12r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_91_adt_net_160209_\);
    
    \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1577_\ : OR3FFT
      port map(A => \I3.un1_REGMAP_30_adt_net_134453_\, B => 
        \I3.N_68\, C => \I3.STATE1_tr24_i_0_a3_28_tz_i\, Y => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1577__net_1\);
    
    MTDIA_pad : IB33
      port map(PAD => MTDIA, Y => MTDIA_c);
    
    \I1.REG_1_284\ : MUX2H
      port map(A => \REGl383r\, B => \I1.REG_74l383r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y => 
        \I1.REG_1_284_net_1\);
    
    TDCDA_padl22r : IB33
      port map(PAD => TDCDA(22), Y => TDCDA_cl22r);
    
    \I2.PIPE1_DT_42_1_IVL2R_1513\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, B => 
        \I2.PIPE1_DT_30l2r_net_1\, C => 
        \I2.PIPE1_DT_42l2r_adt_net_51837_\, Y => 
        \I2.PIPE1_DT_42l2r_adt_net_51839_\);
    
    \I2.FIDl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_431\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl15r);
    
    \I2.DTE_21_1_0_ivl31r\ : AO21
      port map(A => \I2.DTE_1l31r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\, C => 
        \I2.DTE_21_1l31r_adt_net_36417_\, Y => \I2.DTE_21_1l31r\);
    
    \I2.un1_CHAIN_RDY_1_sqmuxa_i\ : OR3
      port map(A => \I2.STATEe_ipl3r\, B => 
        \I2.STATEe_nsl3r_adt_net_22965_\, C => 
        \I2.N_3494_adt_net_90563_\, Y => \I2.N_3494\);
    
    \I2.PIPE6_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_476_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl22r_net_1\);
    
    \I1.REG_74_8_0L380R_1816\ : AND3FTT
      port map(A => \I1.REG_30_sqmuxa\, B => 
        \I1.REG_29_SQMUXA_219\, C => \I1.N_347\, Y => 
        \I1.N_185_9_adt_net_112166_\);
    
    \I3.VDBi_57_0_ivl30r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l30r_net_1\, C
         => \I3.VDBi_57l30r_adt_net_138039_\, Y => 
        \I3.VDBi_57l30r\);
    
    \I3.VDBi_349\ : MUX2L
      port map(A => \I3.VDBil9r_net_1\, B => \I3.VDBi_57l9r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_349_net_1\);
    
    \I3.PIPEB_95_2328\ : NOR2FT
      port map(A => \I3.PIPEBl16r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_95_adt_net_160041_\);
    
    \I1.NWRLUTi\ : DFFS
      port map(CLK => CLK_c, D => \I1.NWRLUTi_57_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.NWRLUTi_net_1\);
    
    \I1.REG_74_0_IVL343R_1870\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l343r_adt_net_116756_\);
    
    \I2.BITCNTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.BITCNT_935\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.BITCNTl5r_net_1\);
    
    \I2.CRC32l24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_819_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l24r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL7R_1480\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl3r\, Y => 
        \I2.PIPE1_DT_42l7r_adt_net_50683_\);
    
    \I2.DTE_1l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_843_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l3r_net_1\);
    
    \I2.un7_bnc_id_1_I_52\ : XOR2
      port map(A => \I2.N_14\, B => \I2.BNC_IDl9r_net_1\, Y => 
        \I2.I_52_0\);
    
    \I2.un7_tdcgda1_3\ : XOR2
      port map(A => \I2.TDCDASl27r_net_1\, B => \I2.TDCl3r_net_1\, 
        Y => \I2.un7_tdcgda1_3_i_i\);
    
    \I2.SRAM_EVNT_n4_0\ : XOR2FT
      port map(A => \I2.SRAM_EVNTl4r_net_1\, B => \I2.N_128_1\, Y
         => \I2.SRAM_EVNT_n4_0_net_1\);
    
    \I2.OFFSET_37_6l2r\ : MUX2L
      port map(A => \I2.N_669\, B => \I2.N_661\, S => 
        \I2.PIPE7_DTL26R_354\, Y => \I2.N_677\);
    
    \I2.CRC32_820\ : MUX2L
      port map(A => \I2.CRC32l25r_net_1\, B => \I2.N_3942\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_820_net_1\);
    
    \I2.ROFFSET_n12\ : XOR2
      port map(A => \I2.N_1378\, B => \I2.N_1379\, Y => 
        \I2.ROFFSET_n12_net_1\);
    
    \I2.REG_1_c14_i\ : AO21FTT
      port map(A => REGl46r, B => \I2.N_138\, C => 
        \I2.N_3843_adt_net_101094_\, Y => \I2.N_3843\);
    
    \I2.EVNT_NUMl7r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_956_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl7r_net_1\);
    
    \I3.PIPEB_101_2322\ : NOR2FT
      port map(A => \I3.PIPEBl22r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_101_adt_net_159789_\);
    
    \I1.REG_74_0_IVL317R_1899\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l317r_adt_net_119303_\);
    
    \I2.L2SERVl1r_1502\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_921_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL13R_609\);
    
    \I2.PIPE4_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl24r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl24r_net_1\);
    
    \I2.DTE_21_1l15r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l15r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l15r_Rd1__net_1\);
    
    \I2.OFFSET_37_12l4r\ : MUX2L
      port map(A => \REGl345r\, B => \I2.N_719\, S => 
        \I2.PIPE7_DTL26R_357\, Y => \I2.N_727\);
    
    \I3.VDBI_57_IVL1R_2268\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => 
        \I3.VDBi_55l1r_net_1\, C => 
        \I3.VDBi_57l1r_adt_net_145945_\, Y => 
        \I3.VDBi_57l1r_adt_net_145946_\);
    
    \I2.SUB9_568\ : MUX2H
      port map(A => \I2.SUB9l0r_net_1\, B => \I2.SUB8l1r_net_1\, 
        S => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_568_net_1\);
    
    \I2.PIPE2_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl4r_net_1\);
    
    \I3.REG_44_i_a2_0l87r\ : NOR2
      port map(A => VDB_inl4r, B => \I3.N_98\, Y => \I3.N_1669\);
    
    \I1.REG_1_207\ : MUX2H
      port map(A => \REGl306r\, B => \I1.REG_74l306r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_207_net_1\);
    
    \I3.PIPEB_90_2333\ : NOR2FT
      port map(A => \I3.PIPEBl11r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_90_adt_net_160251_\);
    
    \I2.un2_evnt_word_I_55\ : AND2
      port map(A => \I2.N_19\, B => \I2.WOFFSETl9r\, Y => 
        \I2.N_16_1\);
    
    \I1.sstate_ns_i_0_a4_0_1_0l0r\ : AND3FTT
      port map(A => \I1.N_349_Rd1__net_1\, B => \I1.N_355\, C => 
        \I1.sstate_ns_i_0_a4_0_1l0r_adt_net_107171_\, Y => 
        \I1.sstate_ns_i_0_a4_0_1l0r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I198_Y\ : XOR2FT
      port map(A => \I2.N411_adt_net_4092__net_1\, B => 
        \I2.SUB_21x21_fast_I198_Y_0\, Y => \I2.SUB8_2l2r\);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_1_sqmuxa_0_a4_i_o2_48_tz\ : MUX2L
      port map(A => LEAD_FLAGl1r, B => LEAD_FLAGl0r, S => 
        \I2.PIPE4_DTl21r_net_1\, Y => \I2.N_2330_tz\);
    
    \I2.PIPE8_DT_16l16r\ : AND2
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855164__net_1\, B => 
        \I2.N_582\, Y => \I2.PIPE8_DT_16l16r_net_1\);
    
    \I1.REG_74_0_ivl401r\ : AO21
      port map(A => \REGl401r\, B => \I1.N_273\, C => 
        \I1.REG_74l401r_adt_net_110014_\, Y => \I1.REG_74l401r\);
    
    \I3.VDBOFFA_31_IV_0L5R_2532\ : AND2
      port map(A => \REGl274r\, B => \I3.REGMAPl31r_net_1\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163660_\);
    
    \I2.STATE1l9r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3208_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1l9r_net_1\);
    
    \I2.NWPIPE5_927\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE4_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE5_305\);
    
    \I3.RAMAD_VME_25\ : MUX2H
      port map(A => RAMAD_VMEl1r, B => \I3.VASl2r_net_1\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_25_net_1\);
    
    \I2.FID_7_0_ivl18r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl18r_net_1\, 
        C => \I2.FID_7l18r_adt_net_17619_\, Y => \I2.FID_7l18r\);
    
    TDCDB_padl0r : IB33
      port map(PAD => TDCDB(0), Y => TDCDB_cl0r);
    
    \I2.I_1341_ca_0_and2\ : AND2FT
      port map(A => \I2.OFFSETL6R_672\, B => \I2.SUB8l9r_net_1\, 
        Y => \I2.N_3545_i_i\);
    
    \I2.ADEl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l12r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl12r);
    
    \I2.PIPE8_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_537_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl9r_net_1\);
    
    \I2.BNCID_VECT_tile_DOUTl1r\ : MUX2L
      port map(A => \I2.DIN_REG1_0l1r\, B => \I2.DOUT_TMP_0l1r\, 
        S => \I2.N_13\, Y => \I2.BNCID_VECTrxl1r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I65_Y\ : AND2
      port map(A => \I2.N302\, B => \I2.N298\, Y => \I2.N333\);
    
    \I2.MIC_ERR_REGSl37r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_366_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl37r_net_1\);
    
    \I2.DTE_21_1_IV_0L12R_1292\ : AO21FTT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_290\, B => 
        \I2.DT_SRAMl12r_net_1\, C => 
        \I2.DTE_21_1l12r_adt_net_38296_\, Y => 
        \I2.DTE_21_1l12r_adt_net_38297_\);
    
    \I2.FID_7_0_IVL18R_956\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl66r, C => 
        \I2.FID_7l18r_adt_net_17611_\, Y => 
        \I2.FID_7l18r_adt_net_17619_\);
    
    \I3.un106_reg_ads_0_a2_0_a2\ : NAND2FT
      port map(A => \I3.N_562\, B => \I3.N_548\, Y => \I3.N_580\);
    
    \I2.PIPE8_DT_540\ : MUX2L
      port map(A => \I2.PIPE8_DTl12r_net_1\, B => 
        \I2.PIPE8_DT_21l12r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_540_net_1\);
    
    \I2.FID_422\ : MUX2H
      port map(A => FID_cl6r, B => \I2.FID_7l6r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        Y => \I2.FID_422_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL9R_1469\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl41r_net_1\, C => 
        \I2.PIPE1_DT_42l9r_adt_net_50179_\, Y => 
        \I2.PIPE1_DT_42l9r_adt_net_50197_\);
    
    \I2.DTO_1_881\ : MUX2L
      port map(A => \I2.DTO_1l7r_Rd1__net_1\, B => 
        \I2.DTO_16_1l7r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834776_Rd1__net_1\, Y
         => \I2.DTO_1l7r\);
    
    \I2.un28_sram_empty_3_0\ : MUX2L
      port map(A => \I2.N_621\, B => \I2.N_620\, S => 
        \I2.RPAGEL14R_612\, Y => \I2.N_622\);
    
    \I2.PIPE9_DT_296\ : MUX2L
      port map(A => \I2.PIPE9_DTl27r_net_1\, B => 
        \I2.PIPE8_DTl27r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_296_net_1\);
    
    \I2.PIPE3_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl15r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl15r_net_1\);
    
    \I1.N_1169_adt_net_854812_\ : BFR
      port map(A => \I1.N_1169_168\, Y => 
        \I1.N_1169_adt_net_854812__net_1\);
    
    \I3.PIPEB_108\ : MUX2H
      port map(A => \I3.PIPEBl29r_net_1\, B => 
        \I3.PIPEB_4l29r_net_1\, S => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_108_net_1\);
    
    \I3.un1_REGMAP_34_0_a2_0_a2\ : NOR2FT
      port map(A => \I3.un1_REGMAP_30\, B => 
        \I3.N_178_ADT_NET_1360__125\, Y => \I3.un1_REGMAP_34\);
    
    \I2.ADEl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl2r);
    
    \I1.N_321_adt_net_855540_\ : BFR
      port map(A => \I1.N_321\, Y => 
        \I1.N_321_adt_net_855540__net_1\);
    
    \I3.VDBi_57l2r_adt_net_145218_\ : NOR3FFT
      port map(A => REGl2r, B => \I3.REGMAPl1r_net_1\, C => 
        \I3.N_2031\, Y => \I3.VDBi_57l2r_adt_net_145218__net_1\);
    
    \I3.PIPEA1_12l25r\ : AND2
      port map(A => DPR_cl25r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854488__net_1\, Y => 
        \I3.PIPEA1_12l25r_net_1\);
    
    \I2.RAMAD1_12l11r\ : MUX2L
      port map(A => \I2.TDCDASl22r_net_1\, B => 
        \I2.TDCDBSl22r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855180__net_1\, Y => 
        \I2.RAMAD1_12l11r_net_1\);
    
    \I1.REG_74_12_220_m9_i\ : OR3FTT
      port map(A => \I1.REG_74_12_300_N_15\, B => 
        \I1.N_145_12_adt_net_123179_\, C => 
        \I1.REG_74_12_220_m9_i_adt_net_127882_\, Y => 
        \I1.REG_74_12_220_m9_i_net_1\);
    
    \I2.TDCDASl9r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl9r, Q => 
        \I2.TDCDASl9r_net_1\);
    
    \I3.REG_1_167\ : MUX2L
      port map(A => VDB_inl18r, B => REGl66r, S => 
        \I3.N_1935_adt_net_855324__net_1\, Y => \I3.REG_1_167_0\);
    
    \I3.N_178_adt_net_1360_\ : OR2FT
      port map(A => \I3.N_2083\, B => 
        \I3.N_178_adt_net_134608__net_1\, Y => 
        \I3.N_178_adt_net_1360__net_1\);
    
    REGl253r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_154_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl253r\);
    
    \I2.RESYN_0_I2_TRGCNT_C3_I_942\ : AOI21TTF
      port map(A => \I2.TRGCNT_i_0_il3r\, B => 
        \I2.un9_tdctrgi_i_0\, C => \I2.N_3763\, Y => 
        \I2.N_3764_adt_net_16233_\);
    
    \I5.sstate2l1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate2se_2_i_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.sstate2l1r_net_1\);
    
    \I2.SUB8l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_510_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l7r_net_1\);
    
    \I2.DTE_0_sqmuxa_i_o2_m6_i_a5_2_i_adt_net_2404_\ : OAI21
      port map(A => \I2.REG_0L3R_ADT_NET_19771_RD1__887\, B => 
        \I2.REG_0L3R_ADT_NET_19773_RD1__888\, C => 
        \I2.END_EVNT10_891\, Y => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_a5_2_i_adt_net_2404__net_1\);
    
    \I3.REG3_0_sqmuxa_adt_net_855628_\ : BFR
      port map(A => \I3.REG3_0_sqmuxa\, Y => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\);
    
    \I2.RAMDT4L5R_3057\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_811\);
    
    \I2.G_EVNT_NUM_n8_i_o2_1288\ : AND2
      port map(A => \I2.N_201\, B => \I2.G_EVNT_NUMl8r_net_1\, Y
         => \I2.N_207_550\);
    
    \I2.N_4293_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I2.N_4293\, SET => 
        CLEAR_STAT_i_0, Q => \I2.N_4293_Rd1__net_1\);
    
    REGl216r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_117_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl216r\);
    
    \I3.VDBml8r\ : MUX2L
      port map(A => \I3.VDBil8r_net_1\, B => \I3.N_150\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml8r_net_1\);
    
    \I3.VDBoffbl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_55_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl3r_net_1\);
    
    \I3.VADm_0_a3l18r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl18r_net_1\, Y => \I3.VADml18r\);
    
    \I2.PIPE1_DTl16r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_743_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl16r_net_1\);
    
    \I2.DTESl21r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl21r, Q => 
        \I2.DTESl21r_net_1\);
    
    \I1.REG_74_12_348_M9_I_1853\ : OAI21FTF
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854400__net_1\, 
        B => \I1.REG_74_1_380_N_16\, C => 
        \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, Y => 
        \I1.REG_74_12_348_m9_i_adt_net_115329_\);
    
    \I2.OFFSET_37_5l2r\ : MUX2L
      port map(A => \REGl399r\, B => \REGl335r\, S => 
        \I2.PIPE7_DTL27R_82\, Y => \I2.N_669\);
    
    \I2.L2SERVl2r_1505\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_920_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL14R_612\);
    
    \I2.PIPE9_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_272_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl3r_net_1\);
    
    \I3.PIPEA_253\ : MUX2L
      port map(A => \I3.PIPEAl22r_net_1\, B => 
        \I3.PIPEA_8l22r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854660__net_1\, Y
         => \I3.PIPEA_253_net_1\);
    
    \I1.REG_74_0_ivl267r\ : AO21
      port map(A => \REGl267r\, B => 
        \I1.N_137_adt_net_854760__net_1\, C => 
        \I1.REG_74l267r_adt_net_124113_\, Y => \I1.REG_74l267r\);
    
    \I2.PIPE5_DT_699\ : MUX2H
      port map(A => \I2.PIPE4_DTl23r_net_1\, B => 
        \I2.PIPE5_DTl23r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_699_net_1\);
    
    \I1.REG_0_SQMUXA_I_0_O2_0_1749\ : NOR2
      port map(A => \I1.BYTECNT_309_net_1\, B => 
        \I1.BYTECNT_310_net_1\, Y => 
        \I1.N_304_adt_net_105325_Ra1_\);
    
    \I3.VDBi_356\ : MUX2L
      port map(A => \I3.VDBil16r_net_1\, B => \I3.VDBi_57l16r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_356_net_1\);
    
    \I3.un1_EVREAD_DS_1_sqmuxa_1\ : OR2FT
      port map(A => \I3.N_1896\, B => 
        \I3.un1_EVREAD_DS_1_sqmuxa_1_adt_net_158292_\, Y => 
        \I3.un1_EVREAD_DS_1_sqmuxa_1_net_1\);
    
    \I2.G_EVNT_NUM_n8_i_a2\ : NOR2
      port map(A => \I2.N_201_adt_net_855048__net_1\, B => 
        \I2.G_EVNT_NUMl8r_net_1\, Y => \I2.N_282\);
    
    \I4.un4_bcnt_I_9\ : XOR2
      port map(A => \I4.bcnt_i_0_il2r_net_1\, B => \I4.N_7\, Y
         => \I4.I_9\);
    
    \I2.FID_420\ : MUX2H
      port map(A => FID_cl4r, B => \I2.FID_7l4r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        Y => \I2.FID_420_net_1\);
    
    \I2.PIPE8_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_552_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl24r_net_1\);
    
    \I5.REG_1_33\ : MUX2L
      port map(A => \I5.TEMPDATAl0r_net_1\, B => REGl420r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_33_net_1\);
    
    FID_P_pad : OB33PH
      port map(PAD => FID_P, A => \GND\);
    
    \I2.FID_7_0_ivl7r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl7r_net_1\, 
        C => \I2.FID_7l7r_adt_net_92841_\, Y => \I2.FID_7l7r\);
    
    \I2.WOFFSETl0r_adt_net_854640_\ : BFR
      port map(A => \I2.WOFFSETl0r_adt_net_854644__net_1\, Y => 
        \I2.WOFFSETl0r_adt_net_854640__net_1\);
    
    \I3.PULSE_46_0_IV_0_0L5R_2292\ : NOR2FT
      port map(A => \I3.REGMAPl10r_net_1\, B => \I3.N_303\, Y => 
        \I3.PULSE_46l5r_adt_net_147097_\);
    
    \I3.VDBi_16_m_i_o3l3r_887\ : OR2
      port map(A => \I3.REGMAPL8R_739\, B => \I3.REGMAPL9R_785\, 
        Y => \I3.N_1907_265\);
    
    \I2.resyn_0_I2_FID_441\ : MUX2H
      port map(A => FID_cl25r, B => \I2.FID_7l25r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\, 
        Y => \I2.FID_441\);
    
    \I2.MIC_REG2L3R_ADT_NET_834020_RD1__2846\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.MIC_REG2_312_adt_net_855644__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2L3R_ADT_NET_834020_RD1__215\);
    
    \I3.VDBi_347\ : MUX2L
      port map(A => \I3.VDBil7r_net_1\, B => \I3.VDBi_57l7r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_347_net_1\);
    
    \I2.PIPE1_DT_737\ : MUX2L
      port map(A => \I2.PIPE1_DTl10r_net_1\, B => 
        \I2.PIPE1_DT_42l10r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854580__net_1\, 
        Y => \I2.PIPE1_DT_737_net_1\);
    
    \I2.TEMPF_1131\ : DFFC
      port map(CLK => CLK_c, D => \I2.TEMPF_760_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TEMPF_393\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I30_Y_1645\ : OR2
      port map(A => \I2.SUB8l12r_net_1\, B => \I2.SUB8l13r_net_1\, 
        Y => \I2.N295_adt_net_68996_\);
    
    \I1.BITCNTL1R_2864\ : DFFC
      port map(CLK => CLK_c, D => \I1.BITCNT_316_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BITCNTL1R_260\);
    
    \I1.REG_74_0_IVL192R_2042\ : AND2
      port map(A => \FBOUTl3r\, B => \I1.REG_4_sqmuxa\, Y => 
        \I1.REG_74l192r_adt_net_131269_\);
    
    \I1.REG_74_0_IVL242R_1984\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_10_sqmuxa_adt_net_854716__net_1\, Y => 
        \I1.REG_74l242r_adt_net_126555_\);
    
    \I3.VDBm_0l27r\ : MUX2L
      port map(A => \I3.PIPEAl27r_net_1\, B => 
        \I3.PIPEBl27r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_169\);
    
    \I1.REG_1_91\ : MUX2H
      port map(A => \REGl190r\, B => \I1.REG_74l190r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, Y => 
        \I1.REG_1_91_net_1\);
    
    \I1.BYTECNTlde_i_a2_i_o2\ : NOR3FFT
      port map(A => \I1.BYTECNT_314_net_1\, B => \I1.N_304_Ra1_\, 
        C => \I1.N_333_Ra1_\, Y => \I1.N_341_Ra1_\);
    
    \I2.EVNT_NUM_c3\ : AND2
      port map(A => \I2.EVNT_NUML3R_597\, B => 
        \I2.EVNT_NUM_c2_net_1\, Y => \I2.EVNT_NUM_c3_net_1\);
    
    \I3.VDBi_40_1l10r\ : MUX2L
      port map(A => REGl127r, B => \I3.VDBi_31l10r_net_1\, S => 
        \I3.REGMAPl16r_net_1\, Y => \I3.N_348\);
    
    \I3.TCNT3_i_0_il6r\ : DFFC
      port map(CLK => CLK_c, D => TCNT3_373, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT3_i_0_il6r_net_1\);
    
    \I2.PIPE1_DT_30l6r\ : MUX2L
      port map(A => \I2.TDCDBSl6r_net_1\, B => 
        \I2.TDCDBSl4r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, Y
         => \I2.PIPE1_DT_30l6r_net_1\);
    
    \I3.RAMDTSl6r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl6r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl6r_net_1\);
    
    \I2.RAMDT4L12R_3043\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_797\);
    
    \I2.MIC_ERR_REGS_367\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl39r_net_1\, B => 
        \I2.MIC_ERR_REGSl38r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_367_net_1\);
    
    \I1.REG_74_0_IV_I_A2_IL206R_2028\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, Y => 
        \I1.N_282_adt_net_130017_\);
    
    \I1.REG_74_0_IVL351R_1862\ : NOR2FT
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_24_sqmuxa_adt_net_854780__net_1\, Y => 
        \I1.REG_74l351r_adt_net_116031_\);
    
    \I1.REG_24_sqmuxa_0_a2\ : OR2
      port map(A => \I1.N_253\, B => \I1.N_240\, Y => 
        \I1.REG_24_sqmuxa\);
    
    \I2.PIPE7_DTL27R_2786\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_79\);
    
    \I2.L2AF3\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2AF2_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L2AF3_net_1\);
    
    \I2.PIPE1_DT_12l17r\ : MUX2L
      port map(A => \I2.TDCDASl17r_net_1\, B => 
        \I2.TDCDASl15r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, Y
         => \I2.PIPE1_DT_12l17r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I76_Y\ : AOI21
      port map(A => \I2.N310\, B => \I2.N313_0\, C => \I2.N309\, 
        Y => \I2.N344\);
    
    TDCDA_padl3r : IB33
      port map(PAD => TDCDA(3), Y => TDCDA_cl3r);
    
    \I3.REG_1_221\ : MUX2L
      port map(A => VDB_inl8r, B => REGl414r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_221_0\);
    
    \I2.un1_STATE1_39\ : AOI21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, B => 
        \I2.N_3887_adt_net_855068__net_1\, C => 
        \I2.un1_STATE1_39_6_i\, Y => \I2.un1_STATE1_39_i_0\);
    
    \I3.REG1l3r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG1_136_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l3r_net_1\);
    
    \I2.TDCDBSl26r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl26r, Q => 
        \I2.TDCDBSl26r_net_1\);
    
    \I2.DT_TEMP_7l31r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854232__net_1\, B => 
        \I2.DT_SRAMl31r_net_1\, Y => \I2.DT_TEMP_7l31r_net_1\);
    
    \I1.REG_10_sqmuxa_adt_net_854720_\ : BFR
      port map(A => \I1.REG_10_sqmuxa\, Y => 
        \I1.REG_10_sqmuxa_adt_net_854720__net_1\);
    
    \I3.VDBi_57_0_iv_0_0_a2l13r_743\ : NAND2FT
      port map(A => \I3.REGMAPl16r_net_1\, B => \I3.N_354_0_129\, 
        Y => \I3.N_2014_121\);
    
    \I2.PIPE5_DT_6l11r\ : MUX2L
      port map(A => \I2.PIPE4_DTl11r_net_1\, B => \I2.N_1080\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\, Y
         => \I2.PIPE5_DT_6l11r_net_1\);
    
    \I2.BITCNT_n1_i\ : NOR3
      port map(A => \I2.ERR_WORDS_RDY_0_sqmuxa\, B => \I2.N_4334\, 
        C => \I2.N_4327\, Y => \I2.N_4322\);
    
    \I1.REG_1_190\ : MUX2H
      port map(A => \REGl289r\, B => \I1.REG_74l289r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\, Y => 
        \I1.REG_1_190_net_1\);
    
    \I2.TDCDBSl4r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl4r, Q => 
        \I2.TDCDBSl4r_net_1\);
    
    \I1.REG_74_0_ivl166r\ : AO21
      port map(A => \REGl166r\, B => \I1.N_41\, C => 
        \I1.REG_74l166r_adt_net_133579_\, Y => \I1.REG_74l166r\);
    
    \I2.MIC_REG1_308\ : MUX2H
      port map(A => \I2.MIC_REG1l7r_net_1\, B => 
        \I2.MTDIAS_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768__net_1\, Y => 
        \I2.MIC_REG1_308_net_1\);
    
    \I2.TOKOUTAS_1247\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKOUTAS_3_i_net_1\, 
        Q => \I2.TOKOUTAS_509\);
    
    \I2.DTE_21_1_IV_0L26R_1241\ : AO21
      port map(A => \I2.DT_SRAMl26r_net_1\, B => 
        \I2.N_199_0_ADT_NET_1054__37\, C => 
        \I2.DTE_21_1l26r_adt_net_36951_\, Y => 
        \I2.DTE_21_1l26r_adt_net_36962_\);
    
    \I2.SUB9_577\ : MUX2H
      port map(A => \I2.SUB9_i_0_il9r\, B => \I2.SUB9_1l9r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_577_net_1\);
    
    \I2.TDCDBSl28r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl28r, Q => 
        \I2.TDCDBSl28r_net_1\);
    
    \I1.REG_74_0_IVL383R_1810\ : AND2
      port map(A => \FBOUTl2r\, B => \I1.REG_28_sqmuxa\, Y => 
        \I1.REG_74l383r_adt_net_111749_\);
    
    \I3.VDBi_360\ : MUX2L
      port map(A => \I3.VDBil20r_net_1\, B => \I3.VDBi_57l20r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_360_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_2671\ : OAI21TTF
      port map(A => \I2.N_72_0\, B => \I2.N_95_0\, C => 
        \I2.N_107_0_adt_net_320362_\, Y => 
        \I2.N525_0_adt_net_318487_\);
    
    \I3.PIPEA_8_0l27r\ : MUX2L
      port map(A => DPR_cl27r, B => \I3.PIPEA1l27r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855356__net_1\, Y => \I3.N_236\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2279\ : NOR3FFT
      port map(A => REGl117r, B => \I3.N_354_0\, C => 
        \I3.REGMAPL55R_782\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146446_\);
    
    RAMAD_padl8r : OB33PH
      port map(PAD => RAMAD(8), A => RAMAD_cl8r);
    
    \I5.REG_1_sqmuxa_0\ : AND2FT
      port map(A => \I5.AIR_CHAIN_net_1\, B => 
        \I5.sstate2_5_sqmuxa\, Y => \I5.REG_1_sqmuxa_0_net_1\);
    
    \I1.REG_74_4l404r\ : AND3FTT
      port map(A => \I1.N_1169_adt_net_854820__net_1\, B => 
        \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Rd1__net_1\, C
         => \I1.REG_74_11_a0l404r_net_1\, Y => \I1.N_273_11_i\);
    
    \I2.N_118_i_1_adt_net_24217_\ : OR3
      port map(A => \I2.SRAM_FULL_593\, B => 
        \I2.sram_empty_0_i_0_i\, C => \I2.sram_empty_2_i_0_i\, Y
         => \I2.N_118_i_1_adt_net_24217__net_1\);
    
    \I2.PIPE7_DTl9r_1589\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL9R_696\);
    
    \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775_\ : OR3FFT
      port map(A => \I2.N_2870\, B => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854628__net_1\, 
        C => \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35789__net_1\, Y
         => \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\);
    
    \I2.resyn_0_I2_FID_439\ : MUX2H
      port map(A => FID_cl23r, B => \I2.FID_7l23r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        Y => \I2.FID_439\);
    
    \I1.NCS0_1_sqmuxa_1_i_0_a4\ : NAND2
      port map(A => \I1.SSTATEL10R_882\, B => \I1.N_328_I_0_498\, 
        Y => \I1.N_436_i_i\);
    
    \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__2754\ : OAI21TTF
      port map(A => \I2.N_176_i_adt_net_855708__net_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, C => 
        \I2.N_4667_1_ADT_NET_1046__34\, Y => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\);
    
    \I3.STATE1_ILLEGAL_2132\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => \I3.N_1180\, C
         => \I3.N_1193_ip_adt_net_136554_\, Y => 
        \I3.N_1193_ip_adt_net_136555_\);
    
    \I3.un141_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_639\, B => \I3.N_551\, Y => 
        \I3.un141_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.FID_7_0_ivl10r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl10r_net_1\, 
        C => \I2.FID_7l10r_adt_net_18371_\, Y => \I2.FID_7l10r\);
    
    \I3.VDBi_57l2r_adt_net_145226_\ : OAI21TTF
      port map(A => GA_cl2r, B => \I3.N_2042\, C => 
        \I3.VDBi_57l2r_adt_net_145225__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145226__net_1\);
    
    \I2.OFFSET_37_22l4r\ : MUX2L
      port map(A => \REGl241r\, B => \REGl177r\, S => 
        \I2.PIPE7_DTL27R_80\, Y => \I2.N_807\);
    
    FCS_pad : OB33PH
      port map(PAD => FCS, A => FCS_c);
    
    \I3.TCNT_383\ : MUX2H
      port map(A => \I3.TCNTl1r_net_1\, B => \I3.TCNT_n1\, S => 
        \I3.TCNTe\, Y => \I3.TCNT_383_net_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I27_Y_1644\ : NOR2
      port map(A => \I2.N_3558_i_net_1\, B => \I2.SUB8l15r_net_1\, 
        Y => \I2.N292_adt_net_68955_\);
    
    \I2.DTE_21_1l20r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l20r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l20r_Rd1__net_1\);
    
    \I2.CRC32_12_il14r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_4026_i_0\, Y => 
        \I2.N_3931\);
    
    \I2.PIPE4_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl19r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl19r_net_1\);
    
    \I1.REG_74_0_IVL389R_1801\ : NOR2FT
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, Y => 
        \I1.REG_74l389r_adt_net_111128_\);
    
    \I2.L2TYPE_4_0l15r\ : AO21
      port map(A => \I2.L2TYPEl15r_net_1\, B => \I2.N_4468\, C
         => \I2.L2TYPE_4l15r_adt_net_66837_\, Y => 
        \I2.L2TYPE_4l15r\);
    
    \I3.VDBi_57l6r_adt_net_143243_\ : NOR2FT
      port map(A => REGl38r, B => \I3.N_2033\, Y => 
        \I3.VDBi_57l6r_adt_net_143243__net_1\);
    
    \I1.REG_6_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_243\, B => \I1.N_259\, Y => 
        \I1.REG_6_sqmuxa\);
    
    \I2.PIPE1_DT_42_0_0l27r_964\ : NOR3
      port map(A => \I2.PIPE1_DT_42_0l27r_net_1\, B => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\, C => \I2.N_12169_i\, Y => 
        \I2.PIPE1_DT_42_3_0L28R_342\);
    
    \I2.WOFFSET_831\ : MUX2L
      port map(A => \I2.WOFFSETl4r_Rd1__net_1\, B => 
        \I2.N_4247_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835312_Rd1__net_1\, Y
         => \I2.WOFFSETl4r\);
    
    \I2.DTO_16_1l16r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l16r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l16r_Rd1__net_1\);
    
    \I2.un1_STATE1_8_i_a3_0_a3\ : NOR3
      port map(A => \I2.STATE1l18r_net_1\, B => 
        \I2.STATE1l5r_net_1\, C => \I2.STATE1l8r_net_1\, Y => 
        \I2.N_3302\);
    
    \I2.LSRAM_INl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_390_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl6r_net_1\);
    
    \I2.EVNT_NUM_955\ : MUX2L
      port map(A => \I2.EVNT_NUMl8r_net_1\, B => 
        \I2.EVNT_NUM_n8_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_955_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A4_0_1563\ : AND2
      port map(A => \I2.RAMDT4L12R_797\, B => 
        \I2.PIPE4_DTl18r_net_1\, Y => \I2.N_41_0_adt_net_55921_\);
    
    \I2.DTE_21_1_IV_0L9R_1308\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.DTE_2_1l9r_net_1\, C
         => \I2.DTE_21_1l9r_adt_net_38625_\, Y => 
        \I2.DTE_21_1l9r_adt_net_38636_\);
    
    \I2.PIPE9_DT_292\ : MUX2L
      port map(A => \I2.PIPE9_DTl23r_net_1\, B => 
        \I2.PIPE8_DTl23r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_292_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL21R_1386\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_340\, B => 
        \I2.EVNT_NUMl5r_net_1\, Y => 
        \I2.PIPE1_DT_42l21r_adt_net_46861_\);
    
    \I2.ENDF_1140_1730\ : DFFC
      port map(CLK => CLK_c, D => \I2.ENDF_712_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ENDF_837\);
    
    \I3.VDBOFFB_30_IV_0L4R_2411\ : AO21
      port map(A => \REGl385r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l4r_adt_net_162322_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162360_\);
    
    \I3.REG_1_184\ : MUX2L
      port map(A => VDB_inl3r, B => \I3.REGl136r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, Y => 
        \I3.REG_1_184_0\);
    
    \I2.INT_ERRAF1_494_1706\ : AND2
      port map(A => \I2.N_3877_adt_net_855268__net_1\, B => 
        \I2.INT_ERRAF1_net_1\, Y => 
        \I2.INT_ERRAF1_494_adt_net_90420_\);
    
    \I1.PAGECNTLDE_0_O4_1758\ : AO21FTT
      port map(A => \I1.SSTATEL4R_418\, B => 
        \I1.N_606_Rd1__net_1\, C => \I1.N_370_adt_net_106310_\, Y
         => \I1.N_370_adt_net_106316_\);
    
    \I0.EV_RESi_1461\ : DFFC
      port map(CLK => CLK_c, D => \I0.EV_RESi_1_net_1\, CLR => 
        \I0.un4_hwresi_i\, Q => EV_RES_C_568);
    
    \I2.SUB9_1_ADD_18x18_fast_I72_Y\ : AO21
      port map(A => \I2.N309\, B => \I2.N306\, C => \I2.N305\, Y
         => \I2.N340\);
    
    \I3.N_178_ADT_NET_1360__2805\ : OR2FT
      port map(A => \I3.N_2083\, B => 
        \I3.N_178_adt_net_134608__net_1\, Y => 
        \I3.N_178_ADT_NET_1360__125\);
    
    \I3.VDBI_57_0_IVL11R_2211\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => 
        \I3.VDBi_55l11r_net_1\, C => 
        \I3.VDBi_57l11r_adt_net_141440_\, Y => 
        \I3.VDBi_57l11r_adt_net_141441_\);
    
    \I2.PIPE10_DT_17_i_0l14r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855596__net_1\, B => 
        \I2.PIPE9_DTl14r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l14r_net_1\);
    
    \I2.DTO_16_1_iv_0_0_1l0r\ : AO21FTT
      port map(A => \I2.DTO_1l0r_net_1\, B => \I2.N_196_53\, C
         => \I2.DTO_16_1_iv_0_0_1l0r_adt_net_35388_\, Y => 
        \I2.DTO_16_1_iv_0_0_1l0r_net_1\);
    
    \I2.DT_SRAM_0l29r\ : MUX2L
      port map(A => \I2.PIPE10_DTl29r_net_1\, B => 
        \I2.PIPE5_DTl29r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, Y => 
        \I2.N_897\);
    
    \I2.EVNT_NUM_n3\ : NOR2
      port map(A => EV_RES_C_569, B => \I2.EVNT_NUM_n3_tz_i\, Y
         => \I2.EVNT_NUM_n3_net_1\);
    
    \I2.DT_TEMPl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_770_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl9r_net_1\);
    
    \I2.CHAINB_EN244_c_0_adt_net_855244_\ : BFR
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\, 
        Y => \I2.CHAINB_EN244_c_0_adt_net_855244__net_1\);
    
    DPR_padl13r : IB33
      port map(PAD => DPR(13), Y => DPR_cl13r);
    
    \I2.INC_EVNT_NUM\ : DFFC
      port map(CLK => CLK_c, D => \I2.INC_EVNT_NUM_759_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.INC_EVNT_NUM_net_1\);
    
    \I2.WPAGEl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_949_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEl14r_net_1\);
    
    \I3.PIPEA_8l9r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854480__net_1\, B => 
        \I3.N_218\, Y => \I3.PIPEA_8l9r_net_1\);
    
    \I2.PIPE1_DT_731\ : MUX2L
      port map(A => \I2.PIPE1_DTl4r_net_1\, B => 
        \I2.PIPE1_DT_42l4r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854584__net_1\, 
        Y => \I2.PIPE1_DT_731_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I8_P0N_i_a2\ : NOR2
      port map(A => \I2.RAMDT4L12R_140\, B => 
        \I2.PIPE4_DTl8r_net_1\, Y => \I2.N_95_0\);
    
    \I3.VDBoffal4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_48_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal4r_net_1\);
    
    \I1.PAGECNTL8R_2940\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_319_adt_net_854860__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL8R_457\);
    
    \I1.REG_1_257\ : MUX2H
      port map(A => \REGl356r\, B => \I1.REG_74l356r_net_1\, S
         => \I1.N_50_0_ADT_NET_1409__20\, Y => 
        \I1.REG_1_257_net_1\);
    
    \I2.TDCDASl22r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl22r, Q => 
        \I2.TDCDASl22r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2538\ : AO21
      port map(A => \REGl210r\, B => 
        \I3.REGMAPl23r_adt_net_855012__net_1\, C => 
        \I3.VDBoffa_31l5r_adt_net_163656_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163691_\);
    
    \I3.REG_1_272\ : MUX2H
      port map(A => VDB_inl0r, B => \I3.REGl91r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_272_0\);
    
    \I2.DTO_16_1_IV_0L13R_1155\ : AO21
      port map(A => \I2.N_197_153\, B => \I2.N_4048\, C => 
        \I2.DTO_16_1l13r_adt_net_32386_\, Y => 
        \I2.DTO_16_1l13r_adt_net_32396_\);
    
    \I2.N_4531_adt_net_1150_\ : AO21FTT
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_215\, C
         => LEAD_FLAGl4r, Y => \I2.N_4531_adt_net_1150__net_1\);
    
    \I2.STATE3_ns_i_o7l11r\ : OR2FT
      port map(A => \I2.STATE3L3R_415\, B => \I2.STOP_RDSRAM_595\, 
        Y => \I2.N_3019\);
    
    \I2.PIPE7_DTl7r_1591\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL7R_698\);
    
    \I2.PIPE6_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_455_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl1r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2468\ : AO21
      port map(A => \REGl326r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l1r_adt_net_162904_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162933_\);
    
    \I3.REG_1l152r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_200_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl152r\);
    
    \I3.VDBi_57l7r_adt_net_143023_\ : AND2
      port map(A => REGl55r, B => \I3.N_2044\, Y => 
        \I3.VDBi_57l7r_adt_net_143023__net_1\);
    
    \I3.un17_reg_ads_0_a2_3_a2\ : NAND3FFT
      port map(A => \I3.VASl4r_net_1\, B => \I3.VASl2r_net_1\, C
         => \I3.N_552\, Y => \I3.N_581\);
    
    \I2.PIPE8_DT_21_i_1l28r\ : AO21
      port map(A => \I2.PIPE8_DT_21_i_1l28r_adt_net_1233__net_1\, 
        B => \I2.PIPE8_DT_21_i_1l28r_adt_net_82784_\, C => 
        \I2.PIPE8_DT_21_i_1l28r_adt_net_82871_\, Y => 
        \I2.PIPE8_DT_21_i_1l28r_net_1\);
    
    \I3.REG_1l156r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_204_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl156r\);
    
    \I2.CRC32_12_i_x2l16r\ : XOR2FT
      port map(A => \I2.CRC32l16r_net_1\, B => \I2.N_3961_i_i\, Y
         => \I2.N_112_i_i_0\);
    
    \I5.REG_1_29\ : MUX2H
      port map(A => \I5.SENS_ADDRl2r_net_1\, B => REGl446r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_29_net_1\);
    
    REGl180r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_81_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl180r\);
    
    \I1.REG_74_9_0_o4_a0l372r\ : OR2FT
      port map(A => \I1.REG_74_9_0_o4_a0_2l372r\, B => 
        \I1.N_1367_i_adt_net_112072_\, Y => \I1.N_347\);
    
    \I2.RAMDT4L10R_2925\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl10r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L10R_442\);
    
    \I2.DTO_16_1_ivl11r\ : OR2
      port map(A => \I2.DTO_16_1l11r_adt_net_32879_\, B => 
        \I2.DTO_16_1l11r_adt_net_32880_\, Y => \I2.DTO_16_1l11r\);
    
    \I2.PIPE1_DT_42_1_IVL20R_1394\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, B => 
        \I2.PIPE1_DT_30l20r_net_1\, C => 
        \I2.PIPE1_DT_42l20r_adt_net_47053_\, Y => 
        \I2.PIPE1_DT_42l20r_adt_net_47068_\);
    
    \I2.PIPE1_DT_42_1_IVL11R_1454\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl27r_net_1\, Y => 
        \I2.PIPE1_DT_42l11r_adt_net_49685_\);
    
    \I2.INT_ERRBF1\ : DFFC
      port map(CLK => CLK_c, D => \I2.INT_ERRBF1_495_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.INT_ERRBF1_net_1\);
    
    \I2.ADEl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl0r);
    
    \I2.PIPE6_DT_0_SQMUXA_I_O4_1597\ : AO21
      port map(A => \I2.N_4543\, B => \I2.N_4673\, C => 
        \I2.N_4551_adt_net_63757_\, Y => 
        \I2.N_4551_adt_net_63759_\);
    
    \I1.REG_1_198\ : MUX2H
      port map(A => \REGl297r\, B => \I1.REG_74l297r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\, Y => 
        \I1.REG_1_198_net_1\);
    
    \I1.PAGECNTl5r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_322_adt_net_854384__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTl5r_net_1\);
    
    \I2.DTESl26r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl26r, Q => 
        \I2.DTESl26r_net_1\);
    
    \I3.VDBi_29l4r\ : AO21
      port map(A => \I3.REGMAPL14R_735\, B => \I3.REGl95r\, C => 
        \I3.VDBi_29l4r_adt_net_144161_\, Y => 
        \I3.VDBi_29l4r_net_1\);
    
    \I2.DTO_16_1_iv_0l2r\ : OA21FTF
      port map(A => \I2.N_182_ADT_NET_1007__386\, B => 
        \I2.N_4193\, C => \I2.DTO_16_1_iv_0_1l2r_net_1\, Y => 
        \I2.DTO_16_1_ivl2r\);
    
    N_1_I3_TCNT2_n7 : XOR2FT
      port map(A => \I3.TCNT2l7r_net_1\, B => \N_1.I3.TCNT2_c6\, 
        Y => \N_1.I3.TCNT2_n7\);
    
    \I2.LSRAM_IN_384\ : MUX2L
      port map(A => \I2.PIPE5_DTl0r_net_1\, B => 
        \I2.LSRAM_INl0r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_384_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL6R_1487\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl38r_net_1\, C => 
        \I2.PIPE1_DT_42l6r_adt_net_50920_\, Y => 
        \I2.PIPE1_DT_42l6r_adt_net_50938_\);
    
    \I3.REG3_126\ : MUX2L
      port map(A => VDB_inl1r, B => \I3.REG3l1r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855624__net_1\, Y => 
        \I3.REG3_126_net_1\);
    
    \I2.PIPE7_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl1r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I177_Y\ : AND2
      port map(A => \I2.N285\, B => \I2.N282\, Y => 
        \I2.N477_adt_net_371248_\);
    
    \I2.STATE3l10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3l11r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE3_i_il10r\);
    
    FID_padl23r : OB33PH
      port map(PAD => FID(23), A => FID_cl23r);
    
    \I2.ROFFSETl0r_1243\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_918_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETL0R_505\);
    
    \I2.TDCDBSl12r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl12r, Q => 
        \I2.TDCDBSl12r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L7R_2357\ : AO21
      port map(A => \REGl388r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l7r_adt_net_161752_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161790_\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854488_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854492__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854488__net_1\);
    
    \I1.REG_0_sqmuxa_i_0_o2\ : NOR3FFT
      port map(A => \I1.PAGECNT_319_adt_net_854864__net_1\, B => 
        \I1.PAGECNT_320_adt_net_854868__net_1\, C => 
        \I1.N_299_Ra1_\, Y => \I1.N_311_i_i_Ra1_\);
    
    \I3.N_1168_adt_net_1509_\ : OR2
      port map(A => \I3.STATE1L10R_728\, B => 
        \I3.STATE1_IPL8R_426\, Y => 
        \I3.N_1168_adt_net_1509__net_1\);
    
    \I3.VDBml18r\ : MUX2L
      port map(A => \I3.VDBil18r_net_1\, B => \I3.N_160\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml18r_net_1\);
    
    \I2.DTE_21_1_IV_0L16R_1271\ : AO21
      port map(A => \I2.DT_SRAMl16r_net_1\, B => 
        \I2.N_199_0_adt_net_1054__net_1\, C => 
        \I2.DTE_21_1l16r_adt_net_37819_\, Y => 
        \I2.DTE_21_1l16r_adt_net_37833_\);
    
    \I2.PIPE1_DT_42_1_IVL1R_1514\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl17r_net_1\, Y => 
        \I2.PIPE1_DT_42l1r_adt_net_52027_\);
    
    \I2.DTO_16_1_iv_0l4r\ : OR2
      port map(A => \I2.DTO_16_1l4r_adt_net_34385_\, B => 
        \I2.DTO_16_1l4r_adt_net_34386_\, Y => \I2.DTO_16_1l4r\);
    
    \I1.RAMDT_SPI_e_0\ : DFFC
      port map(CLK => CLK_c, D => \I1.LOAD_RES_i_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.RAMDT_SPI_E_0\);
    
    \I2.N_4671_adt_net_854600_\ : BFR
      port map(A => \I2.N_4671\, Y => 
        \I2.N_4671_adt_net_854600__net_1\);
    
    REGl308r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_209_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl308r\);
    
    \I3.REGMAPL37R_2932\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un166_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL37R_449\);
    
    \I2.DTE_1l29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_867_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l29r_net_1\);
    
    REGl257r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_158_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl257r\);
    
    \I2.PIPE1_DT_42_1_IVL16R_1412\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_342\, B => 
        \I2.EVNT_NUMl0r_net_1\, Y => 
        \I2.PIPE1_DT_42l16r_adt_net_47837_\);
    
    \I2.N_4535_adt_net_1178_\ : AO21FTT
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_217\, C
         => LEAD_FLAGl0r, Y => \I2.N_4535_adt_net_1178__net_1\);
    
    \I2.DT_TEMP_7l21r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854240__net_1\, B => 
        \I2.DT_SRAMl21r_net_1\, Y => \I2.DT_TEMP_7l21r_net_1\);
    
    VAD_padl16r : OTB33PH
      port map(PAD => VAD(16), A => \I3.VADml16r\, EN => 
        NOEAD_c_i_0);
    
    \I1.REG_74_0_ivl380r\ : AO21
      port map(A => \REGl380r\, B => \I1.N_249\, C => 
        \I1.REG_74l380r_adt_net_112485_\, Y => 
        \I1.REG_74l380r_net_1\);
    
    \I5.un1_sstate1_12_i_a2_1_i_o2\ : AND2
      port map(A => \I5.sstate1l0r_net_1\, B => 
        \I5.COMMANDl2r_net_1\, Y => \I5.N_74\);
    
    \I2.PIPE7_DTl3r_1594\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL3R_701\);
    
    \I2.PIPE1_DT_42_1_ivl28r\ : OR3FTT
      port map(A => \I2.PIPE1_DT_42_3_0l28r\, B => 
        \I2.PIPE1_DT_42l28r_adt_net_45929_\, C => 
        \I2.PIPE1_DT_42l28r_adt_net_45931_\, Y => 
        \I2.PIPE1_DT_42l28r\);
    
    \I3.TCNT2l3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT2_393_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT2l3r_net_1\);
    
    \I2.SRAM_EVNT_c1_i_a2_0\ : NAND3FFT
      port map(A => \I2.SRAM_EVNTl0r_net_1\, B => 
        \I2.SRAM_EVNTl1r_net_1\, C => \I2.N_132\, Y => \I2.N_135\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_2_757\ : AO21
      port map(A => \I2.N_128_adt_net_54290_\, B => 
        \I2.N_128_adt_net_54291_\, C => 
        \I2.N_107_ADT_NET_256840__384\, Y => \I2.N_128_135\);
    
    \I2.SUB9_1_ADD_18x18_fast_I31_Y\ : AO21
      port map(A => \I2.SUB8l12r_net_1\, B => \I2.SUB8l13r_net_1\, 
        C => \I2.N296_adt_net_69573_\, Y => \I2.N296\);
    
    \I2.PIPE8_DT_16l20r\ : MUX2H
      port map(A => \I2.PIPE8_DTl20r_net_1\, B => 
        \I2.PIPE7_DTl20r_net_1\, S => \I2.N_4681_i\, Y => 
        \I2.PIPE8_DT_16l20r_net_1\);
    
    \I2.ADOl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l12r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl12r);
    
    \I2.G_EVNT_NUM_n8_i_o2\ : AND2
      port map(A => \I2.N_201_adt_net_855048__net_1\, B => 
        \I2.G_EVNT_NUMl8r_net_1\, Y => \I2.N_207\);
    
    \I3.un6_asb_1_0_x2\ : XOR2FT
      port map(A => VAD_inl29r, B => GA_cl1r, Y => \I3.N_261_i_0\);
    
    \I2.DT_SRAMl19r\ : MUX2L
      port map(A => \I2.N_887\, B => \I2.PIPE2_DTl19r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.DT_SRAMl19r_net_1\);
    
    \I2.L2AF2\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2AF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L2AF2_net_1\);
    
    SP1_pad : OB33PH
      port map(PAD => SP1, A => \GND\);
    
    \I2.REG_0l3r_adt_net_19773_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.REG_0l3r_adt_net_19773_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.REG_0l3r_adt_net_19773_Rd1__net_1\);
    
    \I2.DTE_1l19r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l19r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l19r_Rd1__net_1\);
    
    \I2.STATE2l1r_adt_net_855124_\ : BFR
      port map(A => \I2.STATE2l1r_adt_net_855132__net_1\, Y => 
        \I2.STATE2l1r_adt_net_855124__net_1\);
    
    \I1.PAGECNTL6R_2855\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_321_adt_net_854880__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL6R_249\);
    
    \I2.RAMDT4L5R_3058\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_812\);
    
    \I2.un21_sram_empty_2\ : XOR2
      port map(A => \I2.RPAGEL14R_616\, B => \I2.L2ARRL2R_604\, Y
         => \I2.un21_sram_empty_2_net_1\);
    
    \I2.REG_1_c0_i\ : OA21FTF
      port map(A => \I2.un8_evread_1_adt_net_855780__net_1\, B
         => \I2.N_119\, C => REGl32r, Y => \I2.N_3829\);
    
    \I1.REG_74_0_ivl286r\ : AO21
      port map(A => \REGl286r\, B => \I1.N_161\, C => 
        \I1.REG_74l286r_adt_net_122205_\, Y => \I1.REG_74l286r\);
    
    \I2.PIPE1_DTl18r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_745_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl18r_net_1\);
    
    DTO_padl6r : IOB33PH
      port map(PAD => DTO(6), A => \I2.DTO_1l6r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl6r);
    
    \I3.UN1_STATE1_13_1_ADT_NET_1351__2804\ : OR3
      port map(A => \I3.un1_STATE1_13_1_adt_net_137890__net_1\, B
         => \I3.un1_STATE1_13_1_adt_net_137896__net_1\, C => 
        \I3.un1_STATE1_13_1_adt_net_137902__net_1\, Y => 
        \I3.UN1_STATE1_13_1_ADT_NET_1351__116\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_3_1556\ : 
        OAI21
      port map(A => \I2.PIPE4_DTL13R_642\, B => 
        \I2.PIPE4_DTL14R_639\, C => \I2.RAMDT4L12R_828\, Y => 
        \I2.N_163_0_adt_net_55087_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I120_Y_0_o2_0\ : NAND2
      port map(A => \I2.N_64_0\, B => \I2.N_89_0_109\, Y => 
        \I2.N_72_0\);
    
    \I2.LSRAM_IN_386\ : MUX2L
      port map(A => \I2.PIPE5_DTl2r_net_1\, B => 
        \I2.LSRAM_INl2r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_386_net_1\);
    
    \I3.PIPEA1_12l20r\ : AND2
      port map(A => DPR_cl20r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854496__net_1\, Y => 
        \I3.PIPEA1_12l20r_net_1\);
    
    \I2.UN1_SRAM_EVNT12_I_1709\ : NOR3
      port map(A => \I2.N_3860\, B => \I2.SRAM_EVNTl4r_net_1\, C
         => \I2.N_128_1\, Y => \I2.N_3823_adt_net_90689_\);
    
    \I2.PIPE3_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl18r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl18r_net_1\);
    
    \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35702_\ : MUX2H
      port map(A => NOESRAME_C_834, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_4146__net_1\, S => 
        \I2.WOFFSETl0r_adt_net_854640__net_1\, Y => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35702__net_1\);
    
    \I2.resyn_0_I2_BITCNT_936\ : MUX2H
      port map(A => \I2.BITCNT_i_0_il4r\, B => \I2.N_4325\, S => 
        \I2.BITCNTe\, Y => \I2.BITCNT_936\);
    
    \I3.VDBml14r\ : MUX2L
      port map(A => \I3.VDBil14r_net_1\, B => \I3.N_156\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml14r_net_1\);
    
    \I2.PIPE1_DTl9r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_736_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl9r_net_1\);
    
    \I1.REG_74_0_IVL286R_1933\ : NOR2FT
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l286r_adt_net_122205_\);
    
    \I2.PIPE6_DT_477\ : MUX2H
      port map(A => \I2.PIPE5_DTl23r_net_1\, B => 
        \I2.PIPE6_DTl23r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_477_net_1\);
    
    \I1.REG_74_0_IVL305R_1913\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l305r_adt_net_120438_\);
    
    \I1.N_311_i_i_Rd1__adt_net_854920_\ : BFR
      port map(A => \I1.N_311_i_i_Rd1__net_1\, Y => 
        \I1.N_311_i_i_Rd1__adt_net_854920__net_1\);
    
    \I2.N_40_adt_net_589803_\ : OAI21
      port map(A => \I2.PIPE4_DTL11R_410\, B => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_2_i_adt_net_271662_\, C
         => \I2.RAMDT4L5R_818\, Y => 
        \I2.N_40_adt_net_589803__net_1\);
    
    \I2.RAMAD1_12l0r\ : MUX2L
      port map(A => \I2.TDCDASl19r_net_1\, B => 
        \I2.TDCDBSl19r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855176__net_1\, Y => 
        \I2.RAMAD1_12l0r_net_1\);
    
    \I1.REG_1_96\ : MUX2H
      port map(A => \REGl195r\, B => \I1.REG_74l195r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\, Y => 
        \I1.REG_1_96_net_1\);
    
    \I5.SCLB_i_a2\ : NAND2FT
      port map(A => \I5.SCL_net_1\, B => \I5.CHAIN_SELECT_net_1\, 
        Y => \I5.N_106\);
    
    \I3.VDBi_57l6r_adt_net_143328_\ : AO21FTT
      port map(A => \I3.N_2017\, B => 
        \I3.VDBi_57l6r_adt_net_3761__net_1\, C => 
        \I3.VDBi_57l6r_adt_net_143314__net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143328__net_1\);
    
    \I3.PIPEA_256\ : MUX2L
      port map(A => \I3.PIPEAl25r_net_1\, B => 
        \I3.PIPEA_8l25r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854656__net_1\, Y
         => \I3.PIPEA_256_net_1\);
    
    DTO_padl30r : IOB33PH
      port map(PAD => DTO(30), A => \I2.DTO_1l30r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl30r);
    
    \I2.STATE1_ns_i_0l13r\ : OAI21FTF
      port map(A => \I2.N_3351\, B => \I2.N_3347_1\, C => 
        \I2.N_3214_i_0_adt_net_22011_\, Y => \I2.N_3214_i_0\);
    
    DTE_padl13r : IOB33PH
      port map(PAD => DTE(13), A => \I2.DTE_1l13r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl13r);
    
    DTE_padl0r : IOB33PH
      port map(PAD => DTE(0), A => \I2.DTE_1l0r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl0r);
    
    \I2.ROFFSET_908\ : MUX2H
      port map(A => \I2.ROFFSETl10r_net_1\, B => 
        \I2.ROFFSET_n10_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_908_net_1\);
    
    \I3.PIPEB_98\ : AO21
      port map(A => DPR_cl19r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855276__net_1\, 
        C => \I3.PIPEB_98_adt_net_159915_\, Y => 
        \I3.PIPEB_98_net_1\);
    
    \I3.PIPEA1_314\ : MUX2L
      port map(A => \I3.PIPEA1l16r_net_1\, B => 
        \I3.PIPEA1_12l16r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__252\, Y => 
        \I3.PIPEA1_314_net_1\);
    
    \I2.resyn_0_I2_TRGCNT_n3_0\ : XOR2
      port map(A => \I2.TRGCNT_i_0_il3r\, B => 
        \I2.un9_tdctrgi_i_0\, Y => \I2.TRGCNT_n3_0\);
    
    \I2.G_EVNT_NUM_n2_i_0_o2\ : NAND3
      port map(A => \I2.G_EVNT_NUM_I_0_IL0R_312\, B => 
        \I2.G_EVNT_NUML1R_306\, C => \I2.G_EVNT_NUML2R_333\, Y
         => \I2.N_187\);
    
    \I3.VDBml27r\ : MUX2L
      port map(A => \I3.VDBil27r_net_1\, B => \I3.N_169\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml27r_net_1\);
    
    \I2.SUB9_584\ : MUX2H
      port map(A => \I2.SUB9l16r_net_1\, B => \I2.SUB9_1l16r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_584_net_1\);
    
    \I1.REG_74_3l404r\ : OR2
      port map(A => \I1.N_273_10_adt_net_114360_\, B => 
        \I1.N_273_10_adt_net_114361_\, Y => \I1.N_273_10\);
    
    \I2.DTE_1_846\ : MUX2L
      port map(A => \I2.DTE_1l6r_Rd1__net_1\, B => 
        \I2.DTE_21_1l6r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836004_Rd1__net_1\, Y => 
        \I2.DTE_1l6r\);
    
    \I2.MIC_ERR_REGS_368\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl40r_net_1\, B => 
        \I2.MIC_ERR_REGSl39r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_368_net_1\);
    
    \I0.CLEARF1_i\ : INV
      port map(A => \I0.CLEARF1_net_1\, Y => \I0.CLEARF1_i_net_1\);
    
    \I3.PIPEA_260\ : MUX2L
      port map(A => \I3.PIPEAl29r_net_1\, B => 
        \I3.PIPEA_8l29r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854652__net_1\, Y
         => \I3.PIPEA_260_net_1\);
    
    \I1.REG_74_0_IVL234R_1992\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_9_sqmuxa_adt_net_854724__net_1\, Y => 
        \I1.REG_74l234r_adt_net_127280_\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855500_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__294\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I138_Y_0\ : AND2FT
      port map(A => \I2.N_100\, B => \I2.N513_i_adt_net_58503_\, 
        Y => \I2.N513_i\);
    
    \I2.DTE_21_1_IV_0_0L4R_1330\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855124__net_1\, B => 
        \I2.EVNT_WORDl0r_net_1\, Y => 
        \I2.DTE_21_1l4r_adt_net_39195_\);
    
    \I2.LSRAM_WADDR_382\ : MUX2L
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => 
        \I2.LSRAM_WADDRl1r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_WADDR_382_net_1\);
    
    \I3.VDBI_57_0_IV_0L21R_2164\ : AND2
      port map(A => \I3.PIPEAl21r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l21r_adt_net_139183_\);
    
    \I2.N_4283_i_0_a2_m1_e_0_857\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__46\, B => 
        \I2.TEMPF_net_1\, Y => \I2.N_4283_I_0_235\);
    
    \I2.CRC32_807\ : MUX2L
      port map(A => \I2.CRC32l12r_net_1\, B => \I2.N_3929\, S => 
        \I2.N_2826_1_ADT_NET_794__331\, Y => \I2.CRC32_807_net_1\);
    
    \I2.EVNT_WORDl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_714_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl1r_net_1\);
    
    \I3.VDBi_57_iv_0_0l7r\ : OR3
      port map(A => \I3.VDBi_57l7r_adt_net_143103_\, B => 
        \I3.VDBi_57l7r_adt_net_143111_\, C => 
        \I3.VDBi_57l7r_adt_net_143112_\, Y => \I3.VDBi_57l7r\);
    
    \I2.NWEN_450\ : MUX2L
      port map(A => NWEN_c, B => \I2.un1_STATE3_8\, S => 
        \I2.N_2989\, Y => \I2.NWEN_450_net_1\);
    
    \I1.REG_1_145\ : MUX2H
      port map(A => \REGl244r\, B => \I1.REG_74l244r_net_1\, S
         => \I1.N_50_0_ADT_NET_1409__293\, Y => 
        \I1.REG_1_145_net_1\);
    
    \I2.PIPE3_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl20r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl20r_net_1\);
    
    \I2.CRC32_12_0_0_x2l28r\ : XOR2FT
      port map(A => \I2.CRC32l28r_net_1\, B => \I2.N_4156_i_i\, Y
         => \I2.N_19_i_0_i_0\);
    
    \I1.REG_74l316r\ : OR2
      port map(A => \I1.REG_20_sqmuxa\, B => 
        \I1.N_193_adt_net_1425__net_1\, Y => \I1.N_185\);
    
    \I2.PIPE1_DTl13r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_740_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl13r_net_1\);
    
    \I2.DTO_1l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_875_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l1r_net_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I124_Y_1651\ : AO21
      port map(A => \I2.N288\, B => \I2.N434_adt_net_3677__net_1\, 
        C => \I2.N287\, Y => \I2.N434_adt_net_69748_\);
    
    \I2.PIPE1_DT_732\ : MUX2L
      port map(A => \I2.PIPE1_DTl5r_net_1\, B => 
        \I2.PIPE1_DT_42l5r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854584__net_1\, 
        Y => \I2.PIPE1_DT_732_net_1\);
    
    \I1.REG_1_147\ : MUX2H
      port map(A => \REGl246r\, B => \I1.REG_74l246r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_147_net_1\);
    
    \I2.PIPE3_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl22r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl22r_net_1\);
    
    \I2.PIPE7_DTl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl18r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl18r_net_1\);
    
    \I3.VDBm_0l14r\ : MUX2L
      port map(A => \I3.PIPEAl14r_net_1\, B => 
        \I3.PIPEBl14r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_156\);
    
    \I3.TCNT4_385\ : MUX2H
      port map(A => \I3.TCNT4l3r_net_1\, B => \I3.TCNT4_n3_net_1\, 
        S => \I3.TICKl2r_net_1\, Y => \I3.TCNT4_385_net_1\);
    
    \I2.BITCNTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.BITCNT_936\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.BITCNT_i_0_il4r\);
    
    \I2.WPAGE_n3\ : XOR2FT
      port map(A => \I2.WPAGEl15r_net_1\, B => 
        \I2.WPAGE_c2_net_1\, Y => \I2.WPAGE_n3_net_1\);
    
    \I2.TOKOUTBS_785\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKOUTBS_3_i_net_1\, 
        Q => \I2.TOKOUTBS_163\);
    
    \I2.SUB8_520_2726\ : AO21
      port map(A => \I2.N298_0\, B => 
        \I2.SUB8_520_adt_net_531295_\, C => 
        \I2.SUB8_520_adt_net_635605_\, Y => 
        \I2.SUB8_520_adt_net_635612_\);
    
    \I1.REG_74_13_388_m8_i\ : OR2
      port map(A => \I1.N_1169_adt_net_854824__net_1\, B => 
        \I1.REG_74_13_388_N_11_adt_net_109571_\, Y => 
        \I1.REG_74_13_388_N_11\);
    
    \I1.REG_1_130\ : MUX2H
      port map(A => \REGl229r\, B => \I1.REG_74l229r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\, Y => 
        \I1.REG_1_130_net_1\);
    
    \I5.sstate1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el8r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l5r_net_1\);
    
    \I2.RAMAD1l5r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_659_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l5r_net_1\);
    
    \I2.MIC_REG2_309\ : MUX2L
      port map(A => \I2.MIC_REG2l1r_net_1\, B => 
        \I2.MIC_REG2l0r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG2_309_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I92_Y_1280\ : NOR2
      port map(A => \I2.N303_0_543\, B => \I2.N307_2\, Y => 
        \I2.N346_0_542\);
    
    \I3.VDBOFFA_48_2564\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal4r_net_1\, Y => 
        \I3.VDBoffa_48_adt_net_163928_\);
    
    \I4.resyn_0_I4_LSRAM_FL_RADDR_10\ : MUX2L
      port map(A => \I4.bcntl1r_net_1\, B => \LSRAM_FL_RADDRl1r\, 
        S => \I4.LSRAM_FL_RADDR_0_sqmuxa_1\, Y => 
        \I4.LSRAM_FL_RADDR_10\);
    
    \I2.L2SERVl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEl15r\);
    
    \I3.PULSE_333\ : MUX2L
      port map(A => PULSEl3r, B => \I3.N_49\, S => 
        \I3.N_1409_adt_net_854744__net_1\, Y => 
        \I3.PULSE_333_net_1\);
    
    \I2.TRGSERVL0R_2948\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.DWACT_ADD_CI_0_partial_sum_1l0r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGSERVL0R_465\);
    
    \I2.resyn_0_I2_FID_445\ : MUX2H
      port map(A => FID_cl29r, B => \I2.FID_7l29r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\, 
        Y => \I2.FID_445\);
    
    \I2.PIPE5_DTl23r_1517\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_699_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL23R_624\);
    
    \I3.VDBi_348\ : MUX2L
      port map(A => \I3.VDBil8r_net_1\, B => \I3.VDBi_57l8r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_348_net_1\);
    
    \I1.REG_74_1l300r\ : AND2
      port map(A => \I1.REG_74_i_o2_i_0l364r_net_1\, B => 
        \I1.REG_74_1l308r_adt_net_120140_\, Y => 
        \I1.REG_74_1l308r\);
    
    \I2.LSRAM_INl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_402_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl18r_net_1\);
    
    \I3.UN12_TCNT3_2643\ : AND3FFT
      port map(A => \I3.TCNT3_i_0_il4r_net_1\, B => 
        \I3.TCNT3l3r_net_1\, C => \I3.un12_tcnt3_adt_net_165618_\, 
        Y => \I3.un12_tcnt3_adt_net_165621_\);
    
    \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768_\ : BFR
      port map(A => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768__net_1\);
    
    \I2.DTO_9_IVL15R_1139\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl15r_net_1\, C => 
        \I2.DTO_9l15r_adt_net_31888_\, Y => 
        \I2.DTO_9l15r_adt_net_31896_\);
    
    \I2.OFFSET_37_19l1r\ : MUX2L
      port map(A => \REGl278r\, B => \REGl214r\, S => 
        \I2.PIPE7_DTL27R_91\, Y => \I2.N_780\);
    
    \I3.REGMAPL57R_3053\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un231_reg_ads_0_a2_4_a3_net_1\, Q => 
        \I3.REGMAPL57R_807\);
    
    \I2.RAMADl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l12r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl12r);
    
    DPR_padl10r : IB33
      port map(PAD => DPR(10), Y => DPR_cl10r);
    
    \I2.MIC_ERR_REGS_331\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl3r_net_1\, B => 
        \I2.MIC_ERR_REGSl2r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_331_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl0r\ : OR2
      port map(A => \I2.PIPE1_DT_42l0r_adt_net_52248_\, B => 
        \I2.PIPE1_DT_42l0r_adt_net_52249_\, Y => 
        \I2.PIPE1_DT_42l0r\);
    
    \I2.MIC_ERR_REGS_339\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl11r_net_1\, B => 
        \I2.MIC_ERR_REGSl10r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\, Y => 
        \I2.MIC_ERR_REGS_339_net_1\);
    
    \I2.TDCDBSl24r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl24r, Q => 
        \I2.TDCDBSl24r_net_1\);
    
    \I2.RESYN_0_I2_LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_948\ : AND2
      port map(A => \I2.PIPE4_DTl22r_net_1\, B => \I2.N_2327_tz\, 
        Y => \I2.N_4524_adt_net_16740_\);
    
    \I3.VDBOFFB_30_IV_0L6R_2368\ : AND2
      port map(A => \REGl307r\, B => \I3.REGMAPl35r_net_1\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161942_\);
    
    \I3.VDBm_i_m2_i_m2l5r\ : MUX2L
      port map(A => \I3.PIPEAl5r_net_1\, B => \I3.PIPEBl5r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_284\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I140_Y_0_1562\ : AND2
      port map(A => \I2.N_2358_tz_tz_adt_net_854956__net_1\, B
         => \I2.N_59_0\, Y => \I2.N519_0_adt_net_55614_\);
    
    \I3.N_1180_adt_net_1502_\ : OR2
      port map(A => \I3.STATE1_ipl4r\, B => \I3.N_1174\, Y => 
        \I3.N_1180_adt_net_1502__net_1\);
    
    \I2.RAMAD_4_0l8r\ : MUX2H
      port map(A => \I2.RAMAD1l8r_net_1\, B => RAMAD_VMEl8r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_535\);
    
    \I2.LEAD_FLAG6_0_sqmuxa_0_a2\ : NAND3FFT
      port map(A => \I2.NWPIPE5_net_1\, B => 
        \I2.PIPE5_DTL30R_621\, C => \I2.PIPE5_DTL31R_620\, Y => 
        \I2.LEAD_FLAG6_0_sqmuxa\);
    
    EV_RESIN_pad : IB33
      port map(PAD => EV_RESIN, Y => EV_RESIN_c);
    
    \I3.REG_1l112r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_293_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl112r);
    
    \I3.REG3_127\ : MUX2L
      port map(A => VDB_inl2r, B => \I3.REG3l2r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855624__net_1\, Y => 
        \I3.REG3_127_net_1\);
    
    \I2.RAMAD_4l6r\ : MUX2L
      port map(A => \I2.N_533\, B => \I1.BYTECNTl6r_net_1\, S => 
        LOAD_RES, Y => \I2.RAMAD_4l6r_net_1\);
    
    \I3.REG3_132\ : MUX2L
      port map(A => VDB_inl7r, B => \I3.REG3l7r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG3_132_net_1\);
    
    \I2.DT_SRAMl30r_adt_net_854200_\ : BFR
      port map(A => \I2.DT_SRAMl30r_net_1\, Y => 
        \I2.DT_SRAMl30r_adt_net_854200__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I46_Y\ : AO21
      port map(A => \I2.N282\, B => \I2.N296_0_adt_net_86403_\, C
         => \I2.N296_0_adt_net_86398_\, Y => \I2.N296_0\);
    
    \I3.TCNT1_i_0_il3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT1_n3_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT1_i_0_il3r_net_1\);
    
    N_1_I3_TCNT2_c2 : AND2
      port map(A => \I3.TCNT2_i_0_il2r_net_1\, B => \I3.TCNT2_c1\, 
        Y => \I3.TCNT2_c2\);
    
    \I3.REG_1l116r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_297_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl116r);
    
    \I1.REG_74_0_iv_0l366r\ : AO21
      port map(A => \REGl366r\, B => \I1.N_660\, C => 
        \I1.REG_74l366r_adt_net_113826_\, Y => \I1.REG_74l366r\);
    
    \I2.ROFFSET_0_sqmuxa_1_0_a7\ : NOR2FT
      port map(A => \I2.STATE3L2R_412\, B => \I2.N_3016\, Y => 
        \I2.ROFFSET_0_sqmuxa_1\);
    
    \I1.REG_74_0_ivl347r\ : AO21
      port map(A => \REGl347r\, B => \I1.N_217\, C => 
        \I1.REG_74l347r_adt_net_116412_\, Y => \I1.REG_74l347r\);
    
    \I1.PAGECNT_n7_i_i_x2\ : XOR2FT
      port map(A => \I1.PAGECNTl7r_net_1\, B => \I1.N_345\, Y => 
        \I1.N_403_i_i_0_i\);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854256_\ : BFR
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854260__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\);
    
    \I2.BNCID_VECTra12_1\ : NOR2
      port map(A => \I2.TRGSERVL0R_467\, B => \I2.TRGSERVL1R_470\, 
        Y => \I2.BNCID_VECTra12_1_net_1\);
    
    \I3.NRDMEBi_230\ : AO21
      port map(A => NRDMEB_c, B => \I3.N_12180_i\, C => 
        \I3.un1_NRDMEBi_2_sqmuxa_3_net_1\, Y => 
        \I3.NRDMEBi_230_net_1\);
    
    \I2.FIRST_TDC_675\ : OR3
      port map(A => \I2.STATE1l9r_net_1\, B => 
        \I2.STATE1l4r_net_1\, C => 
        \I2.FIRST_TDC_675_adt_net_61236_\, Y => 
        \I2.FIRST_TDC_675_net_1\);
    
    \I1.REG_74_0_IVL282R_1937\ : NOR2FT
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l282r_adt_net_122549_\);
    
    \I4.END_FLUSH_1452\ : DFFC
      port map(CLK => CLK_c, D => \I4.END_FLUSH_2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => END_FLUSH_559);
    
    \I2.DT_TEMP_783\ : MUX2H
      port map(A => \I2.DT_TEMPl22r_net_1\, B => 
        \I2.DT_TEMP_7l22r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_783_net_1\);
    
    \I2.N_4530_adt_net_1143_\ : AO21FTT
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_219\, C
         => LEAD_FLAGl5r, Y => \I2.N_4530_adt_net_1143__net_1\);
    
    \I2.L2TYPE_4_IL3R_1636\ : AND2FT
      port map(A => \I2.L2AS_adt_net_855720__net_1\, B => 
        \I2.N_4465\, Y => \I2.N_4449_adt_net_68340_\);
    
    \I2.G_EVNT_NUMl4r_1499\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_930_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUML4R_606\);
    
    \I2.DTO_16_1_IVL10R_1172\ : AO21
      port map(A => \I2.N_197_154\, B => \I2.DT_SRAMl10r_net_1\, 
        C => \I2.DTO_16_1l10r_adt_net_33054_\, Y => 
        \I2.DTO_16_1l10r_adt_net_33066_\);
    
    \I1.REG_1_143\ : MUX2H
      port map(A => \REGl242r\, B => \I1.REG_74l242r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_143_net_1\);
    
    \I1.REG_74_0_IV_0_0L252R_1974\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l252r_adt_net_125605_\);
    
    \I1.REG_74_0_IVL307R_1911\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l307r_adt_net_120266_\);
    
    \I3.PIPEA1_326\ : MUX2L
      port map(A => \I3.PIPEA1l28r_net_1\, B => 
        \I3.PIPEA1_12l28r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, Y => 
        \I3.PIPEA1_326_net_1\);
    
    \I2.PIPE6_DT_457\ : MUX2H
      port map(A => \I2.PIPE5_DTl3r_net_1\, B => 
        \I2.PIPE6_DTl3r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_457_net_1\);
    
    \I3.VDBoff_4_i_il0r\ : MUX2L
      port map(A => \I3.VDBoffbl0r_net_1\, B => 
        \I3.VDBoffal0r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_2064\);
    
    \I2.PIPE1_DT_42_1_IV_0L24R_1374\ : NOR2
      port map(A => \I2.TDCDASl24r_net_1\, B => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        Y => \I2.PIPE1_DT_42_1_iv_0_il24r_adt_net_46513_\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854560_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854560__net_1\);
    
    \I2.RESYN_0_I2_UN1_TRGCNT14_I_938\ : AND3FTT
      port map(A => \I2.N_3794\, B => \I2.TRGCNTl0r_net_1\, C => 
        \I2.N_3760_adt_net_15916_\, Y => 
        \I2.N_3760_adt_net_15910_\);
    
    \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834776_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_0_sqmuxa_i_0_N_3_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834776_Rd1__net_1\);
    
    \I3.un3_noe32wi_0_a2_i_o2_881\ : OR2
      port map(A => \I3.MBLTCYC_422\, B => 
        \I3.N_264_0_ADT_NET_1653_RD1__147\, Y => \I3.N_268_259\);
    
    \I3.PIPEA1_313\ : MUX2L
      port map(A => \I3.PIPEA1l15r_net_1\, B => 
        \I3.PIPEA1_12l15r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__252\, Y => 
        \I3.PIPEA1_313_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I36_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl15r\, B => 
        \I2.PIPE7_DTL15R_690\, Y => \I2.N276\);
    
    \I2.LSRAM_IN_400\ : MUX2L
      port map(A => \I2.PIPE5_DTl16r_net_1\, B => 
        \I2.LSRAM_INl16r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_400_net_1\);
    
    VDB_padl8r : IOB33PH
      port map(PAD => VDB(8), A => \I3.VDBml8r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl8r);
    
    \I2.un7_bnc_id_1_I_66\ : XOR2
      port map(A => \I2.BNC_IDl11r_net_1\, B => \I2.N_4_0\, Y => 
        \I2.I_66_0\);
    
    \I1.REG_74_0_ivl230r\ : AO21
      port map(A => \REGl230r\, B => \I1.N_105\, C => 
        \I1.REG_74l230r_adt_net_127624_\, Y => \I1.REG_74l230r\);
    
    \I3.REG1_135\ : MUX2L
      port map(A => VDB_inl2r, B => \I3.REG1l2r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG1_135_net_1\);
    
    \I3.PIPEA_8l31r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854456__net_1\, B => 
        \I3.N_240\, Y => \I3.PIPEA_8l31r_net_1\);
    
    \I2.un1_NWPIPE7_2_920\ : OR2FT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855156__net_1\, B
         => \I2.un1_NWPIPE7_2_adt_net_73606_\, Y => 
        \I2.UN1_NWPIPE7_2_298\);
    
    \I2.PIPE8_DT_16l17r\ : AND2
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855164__net_1\, B => 
        \I2.N_583\, Y => \I2.PIPE8_DT_16l17r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L0R_2489\ : OR2
      port map(A => \I3.VDBoffb_30l0r_adt_net_163121_\, B => 
        \I3.VDBoffb_30l0r_adt_net_163122_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163127_\);
    
    \I3.VDBoffbl5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_57_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl5r_net_1\);
    
    \I2.RAMAD_4l17r\ : MUX2L
      port map(A => \I2.N_544\, B => 
        \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, S => 
        LOAD_RES_1, Y => \I2.RAMAD_4l17r_net_1\);
    
    TDCGDA_pad : OB33PH
      port map(PAD => TDCGDA, A => TDCGDA_c);
    
    REGl388r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_289_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl388r\);
    
    \I2.DTE_21_1_IV_0_0_18_M7_1218\ : AO21
      port map(A => \I2.DTO_16_1l18r_adt_net_756__net_1\, B => 
        \I2.N_199_0_adt_net_1054__net_1\, C => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35897_\, Y => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35904_\);
    
    \I3.PIPEA1_298\ : MUX2L
      port map(A => \I3.PIPEA1l0r_net_1\, B => 
        \I3.PIPEA1_12l0r_net_1\, S => 
        \I3.un1_STATE2_15_1_adt_net_1342__net_1\, Y => 
        \I3.PIPEA1_298_net_1\);
    
    \I1.PAGECNT_327_825\ : MUX2H
      port map(A => \I1.PAGECNTl0r_adt_net_833884_Rd1__net_1\, B
         => \I1.PAGECNT_n0\, S => 
        \I1.PAGECNTe_adt_net_854900__net_1\, Y => 
        \I1.PAGECNT_327_203\);
    
    \I3.VDBOFFB_30_IV_0L6R_2369\ : AND2
      port map(A => \REGl291r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161946_\);
    
    \I1.REG_74_0_ivl377r\ : AO21
      port map(A => \REGl377r\, B => \I1.N_249\, C => 
        \I1.REG_74l377r_adt_net_112743_\, Y => \I1.REG_74l377r\);
    
    \I3.VDBOFFA_31_IV_0L4R_2562\ : OR3
      port map(A => \I3.VDBoffa_31l4r_adt_net_163885_\, B => 
        \I3.VDBoffa_31l4r_adt_net_163879_\, C => 
        \I3.VDBoffa_31l4r_adt_net_163880_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163889_\);
    
    \I5.REG_1_23\ : MUX2H
      port map(A => \I5.TEMPDATAl4r_net_1\, B => REGl440r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_23_net_1\);
    
    \I3.VDBI_40_0_A3_0L5R_2242\ : OAI21FTF
      port map(A => \I3.REGMAPl17r_adt_net_854292__net_1\, B => 
        \I3.REGl138r\, C => \I3.N_2014\, Y => 
        \I3.N_1772_adt_net_143704_\);
    
    \I2.TOKOUT_FL_674\ : AND2FT
      port map(A => \I2.N_3902\, B => 
        \I2.TOKOUT_FL_674_adt_net_61319_\, Y => 
        \I2.TOKOUT_FL_674_net_1\);
    
    \I2.DT_TEMP_785\ : MUX2H
      port map(A => \I2.DT_TEMPl24r_net_1\, B => 
        \I2.DT_TEMP_7l24r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_785_net_1\);
    
    \I2.G_EVNT_NUMl3r_1137\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_931_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUML3R_399\);
    
    \I3.VDBOFFA_31_IV_0L7R_2499\ : AO21
      port map(A => \REGl188r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.VDBoffa_31l7r_adt_net_163264_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163308_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I15_P0N\ : NAND2FT
      port map(A => \I2.N_3562_i\, B => \I2.SUB8l19r_net_1\, Y
         => \I2.N271\);
    
    \I3.VDBi_57_0_iv_0_0l13r\ : OR2
      port map(A => \I3.VDBi_57l13r_adt_net_140596_\, B => 
        \I3.VDBi_57l13r_adt_net_140597_\, Y => \I3.VDBi_57l13r\);
    
    \I2.PIPE2_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl26r_net_1\);
    
    \I2.DTOSl13r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl13r, Q => 
        \I2.DTOSl13r_net_1\);
    
    \I3.REGMAP_i_0_il24r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un101_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il24r_net_1\);
    
    \I2.DTO_16_1_IV_0_0L18R_1128\ : AO21
      port map(A => \I2.G_EVNT_NUMl2r_net_1\, B => \I2.N_457\, C
         => \I2.DTO_16_1l18r_adt_net_31339_\, Y => 
        \I2.DTO_16_1l18r_adt_net_31345_\);
    
    \I2.CRC32l13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_808_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l13r_net_1\);
    
    \I2.SUB9_570\ : MUX2H
      port map(A => \I2.SUB9l2r_net_1\, B => \I2.SUB9_1l2r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_570_net_1\);
    
    \I1.SBYTE_8_0_a2_il1r\ : AND2
      port map(A => \I1.N_371_i\, B => \I1.N_406\, Y => 
        \I1.N_188\);
    
    \I3.PIPEA_8_0l10r\ : MUX2L
      port map(A => DPR_cl10r, B => \I3.PIPEA1l10r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855352__net_1\, Y => \I3.N_219\);
    
    \I1.REG_1_138\ : MUX2H
      port map(A => \REGl237r\, B => \I1.REG_74l237r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\, Y => 
        \I1.REG_1_138_net_1\);
    
    \I2.N_3836_i_0_adt_net_2390_\ : NAND2FT
      port map(A => \I2.un8_evread_1_adt_net_855780__net_1\, B
         => \I2.N_3849\, Y => \I2.N_3836_i_0_adt_net_2390__net_1\);
    
    \I1.REG_23_sqmuxa_0_a2_m2_e_2\ : AND2FT
      port map(A => \I1.REG_74_1_380_m8_i_0_Rd1__net_1\, B => 
        \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Rd1__net_1\, Y
         => \I1.REG_74_9_0_o4_a0_2l372r\);
    
    \I2.PIPE1_DT_12l13r\ : MUX2L
      port map(A => \I2.TDCDASl13r_net_1\, B => 
        \I2.TDCDASl11r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, Y
         => \I2.PIPE1_DT_12l13r_net_1\);
    
    \I2.CRC32_12_il12r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_116_i_i_0\, Y => 
        \I2.N_3929\);
    
    \I1.REG_1_146\ : MUX2H
      port map(A => \REGl245r\, B => \I1.REG_74l245r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_146_net_1\);
    
    \I2.CRC32_817\ : MUX2L
      port map(A => \I2.CRC32l22r_net_1\, B => \I2.N_3939\, S => 
        \I2.N_2826_1_ADT_NET_794__330\, Y => \I2.CRC32_817_net_1\);
    
    \I2.TOKENTOA_RES_648\ : AO21TTF
      port map(A => \I2.TOKENTOA_RES_net_1\, B => \I2.N_3306\, C
         => \I2.un1_STATE1_28\, Y => \I2.TOKENTOA_RES_648_net_1\);
    
    \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146205_\ : OAI21FTF
      port map(A => \FBOUTl0r\, B => \I3.N_2047\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146197__net_1\, Y
         => \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146205__net_1\);
    
    \I2.TDCDBSl27r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl27r, Q => 
        \I2.TDCDBSl27r_net_1\);
    
    ADO_padl9r : OB33PH
      port map(PAD => ADO(9), A => ADO_cl9r);
    
    REGl183r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_84_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl183r\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l1r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl1r_net_1\, Q => 
        \I2.DIN_REG1_0l1r\);
    
    \I2.MIC_ERR_REGSl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_352_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl23r_net_1\);
    
    \I3.un47_reg_ads_0_a2_0_a2_992\ : OR2FT
      port map(A => \I3.WRITES_8\, B => \I3.N_546_373\, Y => 
        \I3.N_547_370\);
    
    \I2.PIPE1_DT_42_1_ivl3r\ : OR2
      port map(A => \I2.PIPE1_DT_42l3r_adt_net_51636_\, B => 
        \I2.PIPE1_DT_42l3r_adt_net_51637_\, Y => 
        \I2.PIPE1_DT_42l3r\);
    
    \I2.DTO_16_1_IV_0L9R_1174\ : AND2
      port map(A => \I2.DTO_1l9r\, B => \I2.N_196_52\, Y => 
        \I2.DTO_16_1l9r_adt_net_33242_\);
    
    \I2.CHAINA_ERRF1_492\ : MUX2H
      port map(A => CHAINA_ERR_c, B => \I2.CHAINA_ERRF1_net_1\, S
         => \I2.N_3877_adt_net_855268__net_1\, Y => 
        \I2.CHAINA_ERRF1_492_net_1\);
    
    REGl345r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_246_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl345r\);
    
    \I3.N_1906_i_0_0_adt_net_855640_\ : BFR
      port map(A => \I3.N_1906_i_0_0\, Y => 
        \I3.N_1906_i_0_0_adt_net_855640__net_1\);
    
    \I2.PIPE4_DTL10R_3038\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL10R_792\);
    
    \I1.REG_74_0_ivl314r\ : AO21
      port map(A => \REGl314r\, B => \I1.N_185\, C => 
        \I1.REG_74l314r_adt_net_119561_\, Y => \I1.REG_74l314r\);
    
    \I1.BYTECNTL0R_2919\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_314_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTL0R_436\);
    
    \I2.STATE3l7r_1129\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl6r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3L7R_391\);
    
    \I2.OFFSET_37_14l4r\ : MUX2L
      port map(A => \I2.N_735\, B => \I2.N_687\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_743\);
    
    \I2.STATE2_NS_4_0L2R_1050\ : OAI21FTT
      port map(A => \I2.STATE2l0r_net_1\, B => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, C => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854612__net_1\, 
        Y => \I2.STATE2_nsl2r_adt_net_24916_\);
    
    \I3.PIPEBl30r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEB_109_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl30r_net_1\);
    
    \I2.SUB8_520_2723\ : AND3
      port map(A => \I2.N299_0\, B => \I2.N481_adt_net_88982_\, C
         => \I2.SUB8_520_adt_net_531295_\, Y => 
        \I2.SUB8_520_adt_net_635603_\);
    
    \I5.N_64_adt_net_855868_\ : BFR
      port map(A => \I5.N_64\, Y => 
        \I5.N_64_adt_net_855868__net_1\);
    
    \I2.SUB9l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_575_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l7r_net_1\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855420_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__321\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\);
    
    DTE_padl4r : IOB33PH
      port map(PAD => DTE(4), A => \I2.DTE_1l4r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl4r);
    
    \I2.DTO_1l25r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l25r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l25r_Rd1__net_1\);
    
    \I3.PIPEBl18r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_97_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl18r_net_1\);
    
    \I3.PIPEB_79_2344\ : NOR2FT
      port map(A => \I3.PIPEBl0r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_79_adt_net_160713_\);
    
    \I2.RAMDT4L12R_3046\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_800\);
    
    \I2.MIC_ERR_REGS_377\ : MUX2H
      port map(A => \I2.MIC_ERR_REGSl48r_net_1\, B => 
        \I2.MTDIAS_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_377_net_1\);
    
    \I2.OFFSET_37_13l6r\ : MUX2L
      port map(A => \I2.N_729\, B => \I2.N_713\, S => 
        \I2.PIPE7_DTL25R_684\, Y => \I2.N_737\);
    
    \I2.PIPE1_DT_42_1_iv_1l29r\ : NOR2
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.STATE1l3r_net_1\, Y => \I2.PIPE1_DT_42_1l29r\);
    
    \I2.MIC_ERR_REGS_363\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl35r_net_1\, B => 
        \I2.MIC_ERR_REGSl34r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_363_net_1\);
    
    \I3.REG_1_222\ : MUX2L
      port map(A => VDB_inl9r, B => REGl415r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_222_0\);
    
    \I3.REG2_143\ : MUX2L
      port map(A => VDB_inl2r, B => \I3.REG2l2r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG2_143_net_1\);
    
    DTE_pad_i_1l31r : AND2
      port map(A => \I2.DTE_cl_32l31r\, B => \I2.DTE_cll31r\, Y
         => \I2.N_4178_i_0_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2714\ : OR2
      port map(A => \I2.N_152_i_0_adt_net_502546_\, B => 
        \I2.N_152_i_0_adt_net_55873_\, Y => 
        \I2.N_152_i_0_adt_net_610542_\);
    
    \I1.REG_1_270\ : MUX2H
      port map(A => \REGl369r\, B => \I1.REG_74l369r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_270_net_1\);
    
    \I2.CHAINA_EN244_i_0_a2\ : OR2
      port map(A => REGl26r, B => \I2.N_3877\, Y => 
        \I2.CHAINA_EN244_i\);
    
    \I1.SSTATE_NS_1_IV_0_I_A4_2L8R_1765\ : NAND3FFT
      port map(A => \I1.sstatel6r_net_1\, B => 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r_adt_net_107356_\, C => 
        \I1.N_368\, Y => 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r_adt_net_107364_\);
    
    \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__2913\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__382\);
    
    \I1.REG_74_0_ivl244r\ : AO21
      port map(A => \REGl244r\, B => \I1.N_113\, C => 
        \I1.REG_74l244r_adt_net_126383_\, Y => 
        \I1.REG_74l244r_net_1\);
    
    \I1.SBYTE_59\ : MUX2L
      port map(A => \FBOUTl1r\, B => \I1.N_188\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_59_net_1\);
    
    \I3.VDBOFFA_31_IV_0L7R_2508\ : OR3
      port map(A => \I3.VDBoffa_31l7r_adt_net_163315_\, B => 
        \I3.VDBoffa_31l7r_adt_net_163309_\, C => 
        \I3.VDBoffa_31l7r_adt_net_163310_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163319_\);
    
    \I2.un1_STATE2_3_sqmuxa_1_adt_net_839_\ : OAI21TTF
      port map(A => \I2.N_176_i_adt_net_855708__net_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, C => 
        \I2.N_4667_1_ADT_NET_1046__31\, Y => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\);
    
    \I2.resyn_0_I2_TRGCNT_n2\ : XOR2FT
      port map(A => \I2.N_3762\, B => \I2.TRGCNT_n2_0\, Y => 
        \I2.TRGCNT_n2\);
    
    \I1.NCS0_56\ : OR3
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.N_420_i_adt_net_107486_\, C => 
        \I1.NCS0_56_adt_net_133847_\, Y => \I1.NCS0_56_net_1\);
    
    RAMAD_padl10r : OB33PH
      port map(PAD => RAMAD(10), A => RAMAD_cl10r);
    
    \I2.FCNT_947\ : MUX2L
      port map(A => \I2.FCNT_c0\, B => \I2.N_1236\, S => 
        \I2.N_3267\, Y => \I2.FCNT_947_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I188_Y\ : XOR2FT
      port map(A => \I2.N_2\, B => \I2.ADD_21x21_fast_I188_Y_0\, 
        Y => \I2.un27_pipe5_dt0l18r\);
    
    \I1.REG_74_0_ivl389r\ : AO21
      port map(A => \REGl389r\, B => \I1.N_265\, C => 
        \I1.REG_74l389r_adt_net_111128_\, Y => \I1.REG_74l389r\);
    
    \I3.VDBi_16_i_m2l10r\ : MUX2H
      port map(A => REGl26r, B => REG_i_0_il42r, S => 
        \I3.REGMAPl7r_net_1\, Y => \I3.N_2261\);
    
    \I3.VDBm_0l13r\ : MUX2L
      port map(A => \I3.PIPEAl13r_net_1\, B => 
        \I3.PIPEBl13r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_155\);
    
    \I2.LEAD_FLAG6l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_640_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl3r);
    
    \I3.un216_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.N_558\, B => \I3.N_584\, Y => 
        \I3.un216_reg_ads_0_a2_1_a3_net_1\);
    
    \I2.OFFSET_37_29l1r\ : MUX2L
      port map(A => \I2.N_852\, B => \I2.N_740\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l1r\);
    
    \I3.VDBi_31l16r\ : MUX2L
      port map(A => \I3.REGl149r\, B => \I3.VDBi_20l16r\, S => 
        \I3.REGMAPl17r_adt_net_854280__net_1\, Y => 
        \I3.VDBi_31l16r_net_1\);
    
    \I1.REG_74_0_iv_0l362r\ : AO21
      port map(A => \REGl362r\, B => \I1.N_661\, C => 
        \I1.REG_74l362r_adt_net_114697_\, Y => \I1.REG_74l362r\);
    
    \I3.TCNT4_n1\ : XOR2
      port map(A => \I3.TCNT4_i_0_il0r_net_1\, B => 
        \I3.TCNT4l1r_net_1\, Y => \I3.TCNT4_n1_net_1\);
    
    \I2.DTE_1_872\ : MUX2L
      port map(A => \I2.DTE_1l17r_Rd1__net_1\, B => 
        \I2.DTE_21_1l17r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835988_Rd1__net_1\, Y => 
        \I2.DTE_1l17r\);
    
    \I3.VDBml16r\ : MUX2L
      port map(A => \I3.VDBil16r_net_1\, B => \I3.N_158\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml16r_net_1\);
    
    \I3.VDBi_352\ : MUX2L
      port map(A => \I3.VDBil12r_net_1\, B => \I3.VDBi_57l12r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_352_net_1\);
    
    \I1.REG_16_sqmuxa_0_a2_0_719\ : OR2FT
      port map(A => \I1.PAGECNT_0l9r_adt_net_835132_Rd1__net_1\, 
        B => \I1.REG_74_1_A0_0L228R_101\, Y => \I1.N_253_97\);
    
    \I2.CRC32l12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_807_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l12r_net_1\);
    
    GA_padl0r : IB33
      port map(PAD => GA(0), Y => GA_cl0r);
    
    \I2.SUB8_507\ : MUX2H
      port map(A => \I2.SUB8l4r_net_1\, B => \I2.SUB8_2l4r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855148__net_1\, Y => 
        \I2.SUB8_507_net_1\);
    
    \I2.DTESl17r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl17r, Q => 
        \I2.DTESl17r_net_1\);
    
    \I1.REG_74_0_IVL356R_1857\ : NOR2FT
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_24_sqmuxa_adt_net_854776__net_1\, Y => 
        \I1.REG_74l356r_adt_net_115601_\);
    
    \I2.DT_SRAM_0l22r\ : MUX2L
      port map(A => \I2.PIPE10_DTl22r_net_1\, B => 
        \I2.PIPE5_DTL22R_666\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\, Y => 
        \I2.N_890\);
    
    \I2.OFFSET_37_12l7r\ : MUX2L
      port map(A => \REGl348r\, B => \I2.N_722\, S => 
        \I2.PIPE7_DTL26R_355\, Y => \I2.N_730\);
    
    \I3.N_311_adt_net_854748_\ : BFR
      port map(A => \I3.N_311_adt_net_854752__net_1\, Y => 
        \I3.N_311_adt_net_854748__net_1\);
    
    \I3.STATE1_tr24_i_0_o2_1_0\ : AO21
      port map(A => \I3.N_68\, B => 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135385_\, C => 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135386_\, Y => 
        \I3.STATE1_tr24_i_0_o2_1_i\);
    
    \I1.REG_1_273\ : MUX2H
      port map(A => \REGl372r\, B => \I1.REG_74l372r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_273_net_1\);
    
    \I2.PIPE1_DT_728\ : MUX2L
      port map(A => \I2.PIPE1_DTl1r_net_1\, B => 
        \I2.PIPE1_DT_42l1r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854588__net_1\, 
        Y => \I2.PIPE1_DT_728_net_1\);
    
    DTO_padl21r : IOB33PH
      port map(PAD => DTO(21), A => \I2.DTO_1l21r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl21r);
    
    \I1.REG_74L220R_2011\ : AO21
      port map(A => \I1.N_232_1\, B => \I1.N_89_adt_net_128731_\, 
        C => \I1.N_89_adt_net_128717_\, Y => 
        \I1.N_89_adt_net_128732_\);
    
    \I3.N_1935_adt_net_855324_\ : BFR
      port map(A => \I3.N_1935\, Y => 
        \I3.N_1935_adt_net_855324__net_1\);
    
    \I2.G_EVNT_NUMl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_927_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl7r_net_1\);
    
    \I2.DTO_16_1_IV_0L21R_1111\ : AND2
      port map(A => \I2.N_4671_adt_net_854592__net_1\, B => 
        \I2.DT_TEMPl21r_net_1\, Y => 
        \I2.DTO_16_1l21r_adt_net_30536_\);
    
    \I1.REG_74_0_ivl274r\ : AO21
      port map(A => \REGl274r\, B => 
        \I1.N_145_adt_net_854768__net_1\, C => 
        \I1.REG_74l274r_adt_net_123474_\, Y => \I1.REG_74l274r\);
    
    \I3.PIPEAl12r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_243_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl12r_net_1\);
    
    \I2.N_2826_1_adt_net_794_\ : OAI21FTF
      port map(A => \I2.N_4261_304\, B => \I2.N_4282\, C => 
        \I2.N_2826_1_adt_net_40744__net_1\, Y => 
        \I2.N_2826_1_adt_net_794__net_1\);
    
    \I2.EVNT_WORDl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_725_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl12r_net_1\);
    
    \I2.DTE_21_1_iv_0l10r\ : OR3
      port map(A => \I2.DTE_21_1l10r_adt_net_38517_\, B => 
        \I2.DTE_21_1l10r_adt_net_38525_\, C => 
        \I2.DTE_21_1l10r_adt_net_38526_\, Y => \I2.DTE_21_1l10r\);
    
    \I2.BNCID_VECTrff_14_251_0_a2_0\ : AND3
      port map(A => TDCTRG_c, B => \I2.TRGARRl2r_net_1\, C => 
        \I2.TRGARRl3r_net_1\, Y => 
        \I2.BNCID_VECTrff_12_253_0_a2_0\);
    
    \I3.REGMAP_I_0_A2L52R_2095\ : AND3
      port map(A => \I3.N_638_adt_net_134645_\, B => 
        \I3.N_638_adt_net_134643_\, C => 
        \I3.N_638_adt_net_134644_\, Y => 
        \I3.N_638_adt_net_134647_\);
    
    \I2.resyn_0_I2_TRGCNT_n1\ : XOR2FT
      port map(A => \I2.N_3761\, B => \I2.TRGCNT_n1_0\, Y => 
        \I2.TRGCNT_n1\);
    
    \I2.REG_1l39r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n7_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl39r);
    
    REGl243r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_144_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl243r\);
    
    \I3.RAMAD_VME_27\ : MUX2H
      port map(A => RAMAD_VMEl3r, B => \I3.VASl4r_net_1\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_27_net_1\);
    
    \I2.L2TYPE_4_il0r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4452_adt_net_68713_\, C => 
        \I2.N_4452_adt_net_68756_\, Y => \I2.N_4452\);
    
    \I3.PIPEA1_12l16r\ : AND2
      port map(A => DPR_cl16r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854500__net_1\, Y => 
        \I3.PIPEA1_12l16r_net_1\);
    
    \I3.un6_asb_2_0_x2_0_x2\ : XOR2FT
      port map(A => VAD_inl30r, B => GA_cl2r, Y => \I3.N_186_i_0\);
    
    \I1.REG_74_12_300_N_13_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.REG_74_12_300_N_13_Ra1_\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.REG_74_12_300_N_13_Rd1__net_1\);
    
    \I1.COMMAND\ : DFFS
      port map(CLK => CLK_c, D => \I1.COMMAND_52_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.COMMAND_net_1\);
    
    REGl365r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_266_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl365r\);
    
    \I3.REGMAP_I_0_IL30R_3018\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un131_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL30R_772\);
    
    REGl403r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_304_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl403r\);
    
    \I2.DT_TEMPl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_780_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl19r_net_1\);
    
    \I1.REG_74_0_ivl242r\ : AO21
      port map(A => \REGl242r\, B => \I1.N_113\, C => 
        \I1.REG_74l242r_adt_net_126555_\, Y => \I1.REG_74l242r\);
    
    \I1.REG_27_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_240\, B => \I1.N_127_i\, Y => 
        \I1.REG_27_sqmuxa\);
    
    \I3.VDBOFFB_30_IV_0L2R_2444\ : AND2
      port map(A => \REGl343r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        Y => \I3.VDBoffb_30l2r_adt_net_162718_\);
    
    \I2.un28_sram_empty_7_0\ : MUX2L
      port map(A => \I2.N_625\, B => \I2.N_622\, S => 
        \I2.RPAGEL13R_609\, Y => \I2.N_626\);
    
    \I1.REG_74_0_IV_0_0L246R_1980\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.N_592_adt_net_854756__net_1\, Y => 
        \I1.REG_74l246r_adt_net_126121_\);
    
    \I1.REG_74_0_ivl327r\ : AO21
      port map(A => \REGl327r\, B => \I1.N_201\, C => 
        \I1.REG_74l327r_adt_net_118346_\, Y => \I1.REG_74l327r\);
    
    \I3.REG1l2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG1_135_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l2r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I60_Y\ : AO21
      port map(A => \I2.N261_0\, B => \I2.N312_0_adt_net_86445_\, 
        C => \I2.N308_0_adt_net_86497_\, Y => \I2.N310_0\);
    
    \I3.un101_reg_ads_0_a2_0_a2\ : NAND3FTT
      port map(A => \I3.VASl1r_net_1\, B => \I3.N_550\, C => 
        \I3.N_548\, Y => \I3.N_582\);
    
    \I2.DTE_1l9r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l9r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l9r_Rd1__net_1\);
    
    \I2.CRC32_826\ : MUX2L
      port map(A => \I2.CRC32l31r_net_1\, B => \I2.N_3948\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_826_net_1\);
    
    \I2.PIPE8_DT_550\ : MUX2L
      port map(A => \I2.PIPE8_DTl22r_net_1\, B => 
        \I2.PIPE8_DT_21l22r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_550_net_1\);
    
    \I2.PIPE7_DTl15r_1583\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl15r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL15R_690\);
    
    \I2.PIPE6_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_454_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl0r_net_1\);
    
    \I3.TCNT4_c2\ : NAND2
      port map(A => \I3.TCNT4_i_0_il2r_net_1\, B => 
        \I3.TCNT4_c1_net_1\, Y => \I3.TCNT4_c2_net_1\);
    
    \I1.REG_74_0_ivl235r\ : AO21
      port map(A => \REGl235r\, B => \I1.N_105\, C => 
        \I1.REG_74l235r_adt_net_127194_\, Y => \I1.REG_74l235r\);
    
    \I5.un1_SENS_ADDR_1_I_14\ : XOR2
      port map(A => \I5.DWACT_ADD_CI_0_g_array_1l0r\, B => 
        \I5.SENS_ADDRl2r_net_1\, Y => \I5.I_14\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I26_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl5r\, B => \I2.PIPE7_DTL5R_700\, 
        Y => \I2.N246_0\);
    
    \I2.L2TYPE_4_IL7R_1629\ : AND2FT
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4466\, Y => \I2.N_4445_adt_net_67839_\);
    
    \I1.REG_74_7_0l188r\ : NAND3FTT
      port map(A => \I1.REG_30_sqmuxa\, B => 
        \I1.REG_29_SQMUXA_219\, C => 
        \I1.N_1367_i_adt_net_854516__net_1\, Y => \I1.N_97_6\);
    
    \I2.ADO_3l5r\ : MUX2L
      port map(A => \I2.WOFFSETl6r\, B => \I2.ROFFSETl6r_net_1\, 
        S => NOESRAME_C_243, Y => \I2.ADO_3l5r_net_1\);
    
    DPR_padl14r : IB33
      port map(PAD => DPR(14), Y => DPR_cl14r);
    
    \I1.REG_74_5_404_m1_e_0_902\ : NOR2FT
      port map(A => \I1.PAGECNT_0l8r_adt_net_834720_Rd1__net_1\, 
        B => \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__361\, Y => 
        \I1.REG_74_5_404_M1_E_0_280\);
    
    \I2.CRC32_12_i_0_m2l6r\ : MUX2L
      port map(A => \I2.DT_TEMPl6r_net_1\, B => 
        \I2.DT_SRAMl6r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854440__net_1\, Y => 
        \I2.N_225_i_i\);
    
    \I1.REG_74_0_IVL289R_1930\ : NOR2FT
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l289r_adt_net_121947_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I5_P0N_i_a4\ : OR2
      port map(A => \I2.RAMDT4L12R_146\, B => 
        \I2.PIPE4_DTl5r_adt_net_854412__net_1\, Y => \I2.N_89_0\);
    
    \I2.PIPE5_DT_695\ : MUX2L
      port map(A => \I2.PIPE5_DTl19r_net_1\, B => 
        \I2.PIPE5_DT_6l19r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_695_net_1\);
    
    \I1.REG_74_0_ivl396r\ : AO21
      port map(A => \REGl396r\, B => \I1.N_265\, C => 
        \I1.REG_74l396r_adt_net_110526_\, Y => 
        \I1.REG_74l396r_net_1\);
    
    \I2.DTE_21_1_IV_2L2R_1339\ : OAI21TTF
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855208__net_1\, 
        B => \I2.DT_TEMPl2r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il2r_adt_net_39443_\, Y => 
        \I2.DTE_21_1_iv_2_il2r_adt_net_39452_\);
    
    \I2.DTE_21_1_IV_0_0L22R_1252\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855196__net_1\, 
        B => \I2.DT_TEMPl22r_net_1\, C => 
        \I2.DTO_16_1l22r_adt_net_30352_\, Y => 
        \I2.DTE_21_1l22r_adt_net_37393_\);
    
    \I2.REG_0l3r_adt_net_848__adt_net_854208_\ : BFR
      port map(A => \I2.REG_0l3r_adt_net_848__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__adt_net_854208__net_1\);
    
    \I2.PIPE8_DT_16_0l12r\ : MUX2H
      port map(A => \I2.PIPE8_DTl12r_net_1\, B => 
        \I2.PIPE7_DTl12r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_578\);
    
    \I4.FLUSH_3_932\ : AND2
      port map(A => \I4.un1_FLUSH_1_sqmuxa_1_net_1\, B => FLUSH, 
        Y => \I4.FLUSH_3_adt_net_15593_\);
    
    \I2.RAMADl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l4r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl4r);
    
    \I3.VDBi_31l4r\ : MUX2L
      port map(A => \I3.REGl137r\, B => \I3.VDBi_29l4r_net_1\, S
         => \I3.REGMAPl17r_adt_net_854292__net_1\, Y => 
        \I3.VDBi_31l4r_net_1\);
    
    \I2.REG_0L3R_ADT_NET_19773_RD1__2883\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.REG_0l3r_adt_net_19773_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.REG_0L3R_ADT_NET_19773_RD1__315\);
    
    \I3.VDBOFFA_31_IV_0L2R_2591\ : AO21
      port map(A => \REGl223r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.VDBoffa_31l2r_adt_net_164222_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164260_\);
    
    \I2.majority_reg_il5r\ : OAI21TTF
      port map(A => \I2.MIC_REG2_i_0_il5r_net_1\, B => 
        \I2.MIC_REG1l5r_net_1\, C => \I2.N_4431_adt_net_22416_\, 
        Y => \I2.N_4431\);
    
    \I2.END_TDC6_268\ : MUX2L
      port map(A => END_TDC, B => \I2.END_TDC5_net_1\, S => 
        END_FLUSH_560, Y => \I2.END_TDC6_268_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I57_Y_0_o2\ : AO21
      port map(A => \I2.N_85\, B => \I2.N357_adt_net_54497_\, C
         => \I2.N357_adt_net_54538_\, Y => \I2.N357\);
    
    \I2.STATE3l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl13r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE3l0r_net_1\);
    
    \I2.STATE2l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl1r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2l4r_net_1\);
    
    \I2.G_EVNT_NUMl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_933_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl1r_net_1\);
    
    \I2.L2TYPE_4_il10r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855716__net_1\, B => 
        \I2.N_4442_adt_net_67433_\, C => 
        \I2.N_4442_adt_net_67476_\, Y => \I2.N_4442\);
    
    REGl318r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_219_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl318r\);
    
    \I3.REGMAPL44R_2934\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un201_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL44R_451\);
    
    \I2.PIPE7_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl0r_net_1\);
    
    \I2.PIPE1_DT_743\ : MUX2L
      port map(A => \I2.PIPE1_DTl16r_net_1\, B => 
        \I2.PIPE1_DT_42l16r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854572__net_1\, 
        Y => \I2.PIPE1_DT_743_net_1\);
    
    \I2.ADO_3l6r\ : MUX2L
      port map(A => \I2.WOFFSETl7r\, B => \I2.ROFFSETl7r_net_1\, 
        S => NOESRAME_C_243, Y => \I2.ADO_3l6r_net_1\);
    
    \I3.PIPEA_8l17r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854468__net_1\, B => 
        \I3.N_226\, Y => \I3.PIPEA_8l17r_net_1\);
    
    \I2.ROFFSETe_0_adt_net_27187_\ : OR3
      port map(A => \I2.ROFFSET_0_sqmuxa_1\, B => 
        \I2.ROFFSETe_0_adt_net_27175__net_1\, C => 
        \I2.ROFFSETe_0_adt_net_27185__net_1\, Y => 
        \I2.ROFFSETe_0_adt_net_27187__net_1\);
    
    \I2.LSRAM_INl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_397_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl13r_net_1\);
    
    \I1.REG_74_1L300R_1909\ : NOR3FTT
      port map(A => \I1.N_347_adt_net_854788__net_1\, B => 
        \I1.N_97_2\, C => \I1.REG_74_12_300_N_11\, Y => 
        \I1.REG_74_1l308r_adt_net_120140_\);
    
    \I2.TDCDBSl9r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl9r, Q => 
        \I2.TDCDBSl9r_net_1\);
    
    \I1.REG_74_0_ivl272r\ : AO21
      port map(A => \REGl272r\, B => 
        \I1.N_145_adt_net_854768__net_1\, C => 
        \I1.REG_74l272r_adt_net_123646_\, Y => \I1.REG_74l272r\);
    
    \I2.DT_SRAMl21r\ : MUX2L
      port map(A => \I2.N_889\, B => \I2.PIPE2_DTl21r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl21r_net_1\);
    
    \I1.REG_74_0_IV_0L269R_1954\ : AND2
      port map(A => \REGl269r\, B => 
        \I1.N_145_adt_net_854772__net_1\, Y => 
        \I1.REG_74l269r_adt_net_123904_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I175_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L5R_139\, B => 
        \I2.PIPE4_DTl5r_adt_net_854412__adt_net_855600__net_1\, Y
         => \I2.ADD_21x21_fast_I175_Y_0\);
    
    \I1.REG_74_0_iv_0_0l258r\ : AO21
      port map(A => \REGl258r\, B => \I1.N_658\, C => 
        \I1.REG_74l258r_adt_net_124970_\, Y => \I1.REG_74l258r\);
    
    \I3.REG_1l85r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_266_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl85r);
    
    \I2.OFFSET_37_24l4r\ : MUX2L
      port map(A => \I2.N_815\, B => \I2.N_807\, S => 
        \I2.PIPE7_DTL26R_358\, Y => \I2.N_823\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I121_Y_i_o2\ : AND3
      port map(A => \I2.N_28\, B => \I2.N_64\, C => \I2.N_158_0\, 
        Y => \I2.N_29_i\);
    
    \I2.PIPE4_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl8r_net_1\);
    
    \I2.DTE_1_840\ : MUX2L
      port map(A => \I2.DTE_1l0r_net_1\, B => 
        \I2.DTE_21_1_iv_i_0l0r\, S => \I2.N_2868_1\, Y => 
        \I2.DTE_1_840_net_1\);
    
    \I2.CHB_DATA8_503\ : MUX2L
      port map(A => \I2.CHB_DATA8_net_1\, B => \I2.N_4397\, S => 
        \I2.NWPIPE7_net_1\, Y => \I2.CHB_DATA8_503_net_1\);
    
    \I2.DTO_16_1_IV_0_1L2R_1206\ : NOR2
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620__net_1\, 
        B => \I2.DT_TEMPl2r_net_1\, Y => 
        \I2.DTO_16_1_iv_0_1l2r_adt_net_34862_\);
    
    \I2.DTE_21_1_IV_0_0L7R_1319\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l7r\, C
         => \I2.DTE_21_1l7r_adt_net_38872_\, Y => 
        \I2.DTE_21_1l7r_adt_net_38873_\);
    
    \I2.ROFFSET_247\ : NAND3FTT
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855704__net_1\, B => 
        \I2.ROFFSETl11r_net_1\, C => \I2.ROFFSET_c10_net_1\, Y
         => \I2.N_1378\);
    
    \I2.REG_0l3r_adt_net_19771_Ra1_\ : AND2
      port map(A => \I3.REG1_136_net_1\, B => \I3.REG2_144_net_1\, 
        Y => \I2.REG_0l3r_adt_net_19771_Ra1__net_1\);
    
    \I5.REG_1_19\ : MUX2H
      port map(A => \I5.TEMPDATAl0r_net_1\, B => REGl436r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\, Y
         => \I5.REG_1_19_net_1\);
    
    \I3.DSSF1\ : DFFS
      port map(CLK => CLK_c, D => \I3.DSSF1_42_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.DSSF1_net_1\);
    
    \I3.REG_44_i_a2_0l84r\ : NOR2
      port map(A => VDB_inl1r, B => \I3.N_98\, Y => \I3.N_1663\);
    
    \I3.STATE1l6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl4r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl6r\);
    
    \I3.PIPEBl6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_85_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl6r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I178_Y\ : XOR2FT
      port map(A => \I2.N_3_0\, B => 
        \I2.ADD_21x21_fast_I178_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l8r\);
    
    \I2.WPAGE_948\ : MUX2H
      port map(A => \I2.WPAGEl15r_net_1\, B => 
        \I2.WPAGE_n3_net_1\, S => 
        \I2.WPAGEe_adt_net_855056__net_1\, Y => 
        \I2.WPAGE_948_net_1\);
    
    \I2.RAMDT4L12R_3042\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_796\);
    
    \I1.REG_74_0_ivl300r\ : AO21
      port map(A => \REGl300r\, B => \I1.N_169\, C => 
        \I1.REG_74l300r_adt_net_120868_\, Y => 
        \I1.REG_74l300r_net_1\);
    
    \I2.REG_1_c10_i_a2_0\ : AND3FFT
      port map(A => REG_i_0_il42r, B => REGl41r, C => \I2.N_129\, 
        Y => \I2.N_131\);
    
    \I2.DTE_1l10r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l10r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l10r_Rd1__net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I154_Y_0_2692\ : AND2FT
      port map(A => \I2.ADD_21x21_fast_I136_Y_0_o2_m4_1_i\, B => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_4_adt_net_56769_\, Y
         => \I2.N502_i_0_adt_net_490398_\);
    
    \I5.DATA_12l8r\ : MUX2L
      port map(A => REGl125r, B => \I5.SBYTEl0r_net_1\, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l8r_net_1\);
    
    \I2.PIPE4_DTl8r_adt_net_854556_\ : BFR
      port map(A => \I2.PIPE4_DTl8r_net_1\, Y => 
        \I2.PIPE4_DTl8r_adt_net_854556__net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_1575\ : AND3
      port map(A => \I2.N_107_0\, B => 
        \I2.N_2358_tz_tz_adt_net_854952__net_1\, C => 
        \I2.N525_0_adt_net_58018_\, Y => 
        \I2.N525_0_adt_net_58015_\);
    
    \I2.OFFSET_37_11l6r\ : MUX2L
      port map(A => \REGl379r\, B => \REGl315r\, S => 
        \I2.PIPE7_DTL27R_77\, Y => \I2.N_721\);
    
    \I2.L2TYPEl15r_1557\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_604_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL15R_664\);
    
    \I2.DTE_1_852\ : MUX2L
      port map(A => \I2.DTE_1l12r_Rd1__net_1\, B => 
        \I2.DTE_21_1l12r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, Y => 
        \I2.DTE_1l12r\);
    
    \I2.OFFSET_37_23l6r\ : MUX2L
      port map(A => \REGl275r\, B => \REGl211r\, S => 
        \I2.PIPE7_DTL27R_87\, Y => \I2.N_817\);
    
    \I2.DTE_21_1_IV_0_0L17R_1221\ : AND2
      port map(A => \I2.N_188\, B => 
        \I2.N_199_0_ADT_NET_1054__36\, Y => 
        \I2.DTE_21_1l17r_adt_net_36140_\);
    
    \I1.REG_74_0_IVL402R_1787\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_30_sqmuxa_adt_net_854376__net_1\, Y => 
        \I1.REG_74l402r_adt_net_109928_\);
    
    \I1.un1_pulse_1_i_a2_0_a4\ : NAND2FT
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.N_380\, Y => \I1.N_1207\);
    
    \I2.PIPE8_DT_529\ : MUX2L
      port map(A => \I2.PIPE8_DTl1r_net_1\, B => 
        \I2.PIPE8_DT_21l1r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_529_net_1\);
    
    \I2.DTE_1l26r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l26r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l26r_Rd1__net_1\);
    
    \I2.TRAIL_MIS6\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRAIL_MIS6_491\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRAIL_MIS6_net_1\);
    
    \I2.DT_TEMPl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_779_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl18r_net_1\);
    
    REGl263r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_164_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl263r\);
    
    \I1.REG_74_0_IVL313R_1903\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l313r_adt_net_119647_\);
    
    \I3.REG_1_ml74r\ : AND2
      port map(A => REGl74r, B => 
        \I3.REGMAPl9r_adt_net_854304__net_1\, Y => 
        \I3.VDBi_20l26r\);
    
    \I2.BNC_IDl3r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_13_2\, CLR => 
        \I2.N_4624_i_0\, SET => \I2.N_4613_i_0\, Q => 
        \I2.BNC_IDl3r_net_1\);
    
    \I2.BNCID_VECTROR_1422\ : OR2
      port map(A => \I2.BNCID_VECTror_adt_net_48365_\, B => 
        \I2.BNCID_VECTror_adt_net_48367_\, Y => 
        \I2.BNCID_VECTror_adt_net_48326_\);
    
    \I3.STATE1_ipl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl7r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl3r_net_1\);
    
    \I3.un1_STATE2_15_1_adt_net_147701_\ : AND3FTT
      port map(A => \I3.EVREAD_DS_net_1\, B => 
        \I3.STATE2l0r_net_1\, C => \I3.END_PK_net_1\, Y => 
        \I3.un1_STATE2_15_1_adt_net_147701__net_1\);
    
    \I2.DTE_21_1_IV_0L12R_1293\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.N_93_i_0\, C => 
        \I2.DTE_21_1l12r_adt_net_38279_\, Y => 
        \I2.DTE_21_1l12r_adt_net_38298_\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2525\ : OR2
      port map(A => \I3.N_2070_adt_net_163501_\, B => 
        \I3.N_2070_adt_net_163502_\, Y => 
        \I3.N_2070_adt_net_163507_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I177_Y\ : XOR2
      port map(A => \I2.N531\, B => \I2.ADD_21x21_fast_I177_Y_0\, 
        Y => \I2.un27_pipe5_dt0l7r\);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_1_sqmuxa_0_a4_i\ : OR2
      port map(A => END_FLUSH_560, B => \I2.N_4524\, Y => 
        \I2.N_4642\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_A2_2_1558\ : 
        AND3FFT
      port map(A => \I2.N_140_0\, B => \I2.N_139_0\, C => 
        \I2.N_72_0_108\, Y => \I2.N_128_0_adt_net_55238_\);
    
    \I2.BITCNTlde_0_a5\ : AND2
      port map(A => \I2.STATE5l0r_net_1\, B => 
        \I2.W_ERR_WORDS_net_1\, Y => \I2.ERR_WORDS_RDY_0_sqmuxa\);
    
    \I1.REG_74_0_ivl315r\ : AO21
      port map(A => \REGl315r\, B => \I1.N_185\, C => 
        \I1.REG_74l315r_adt_net_119475_\, Y => \I1.REG_74l315r\);
    
    \I2.G_EVNT_NUM_N4_I_0_1054\ : OA21TTF
      port map(A => \I2.N_189\, B => \I2.G_EVNT_NUMl4r_net_1\, C
         => EV_RES_C_568, Y => \I2.N_4344_adt_net_26298_\);
    
    \I2.DTE_21_1_iv_0l21r\ : AO21
      port map(A => \I2.DTE_1l21r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.DTE_21_1l21r_adt_net_37497_\, Y => \I2.DTE_21_1l21r\);
    
    \I2.un1_STATE3_10_0_i\ : INV
      port map(A => \I2.STATE3l9r_net_1\, Y => \I2.STATE3_il9r\);
    
    \I2.DTO_1_901\ : MUX2L
      port map(A => \I2.DTO_1l27r_Rd1__net_1\, B => 
        \I2.DTO_16_1l27r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834756_Rd1__net_1\, Y
         => \I2.DTO_1l27r\);
    
    \I2.MIC_ERR_REGS_362\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl34r_net_1\, B => 
        \I2.MIC_ERR_REGSl33r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_362_net_1\);
    
    TDCDB_padl7r : IB33
      port map(PAD => TDCDB(7), Y => TDCDB_cl7r);
    
    \I2.PIPE4_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl5r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl5r_net_1\);
    
    \I2.OFFSET_37_12l2r\ : MUX2L
      port map(A => \REGl343r\, B => \I2.N_717\, S => 
        \I2.PIPE7_DTL26R_359\, Y => \I2.N_725\);
    
    \I3.VDBOFFB_30_IV_0L0R_2483\ : AO21
      port map(A => \REGl381r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l0r_adt_net_163082_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163120_\);
    
    \I2.un1_STATE1_40_1_adt_net_45405_\ : OR3
      port map(A => \I2.STATE1L17R_574\, B => 
        \I2.STATE1_i_0_il15r\, C => \I2.N_3890\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45405__net_1\);
    
    \I2.REG_1_c8_i_o2\ : OR3FFT
      port map(A => REGl39r, B => REGl40r, C => \I2.N_3849\, Y
         => \I2.N_3852\);
    
    REGl251r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_152_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl251r\);
    
    \I3.REGMAPl41r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un186_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPl41r_net_1\);
    
    \I2.DTE_cl_65_il31r\ : AOI21FTF
      port map(A => \I2.DTE_cll31r\, B => 
        \I2.un1_DTO_cl_1_sqmuxa_2\, C => \I2.N_4182\, Y => 
        \I2.N_4180_i_0\);
    
    DPR_padl16r : IB33
      port map(PAD => DPR(16), Y => DPR_cl16r);
    
    \I2.PIPE1_DT_756\ : MUX2L
      port map(A => \I2.PIPE1_DTl29r_net_1\, B => 
        \I2.PIPE1_DT_42l29r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854560__net_1\, 
        Y => \I2.PIPE1_DT_756_net_1\);
    
    \I1.REG_74_0_ivl224r\ : AO21
      port map(A => \REGl224r\, B => \I1.N_97\, C => 
        \I1.REG_74l224r_adt_net_128308_\, Y => \I1.REG_74l224r\);
    
    \I2.MIC_ERR_REGS_357\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl29r_net_1\, B => 
        \I2.MIC_ERR_REGSl28r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_357_net_1\);
    
    \I2.OFFSET_37_22l7r\ : MUX2L
      port map(A => \REGl244r\, B => \REGl180r\, S => 
        \I2.PIPE7_DTL27R_76\, Y => \I2.N_810\);
    
    \I2.N_2358_tz_tz_adt_net_854952_\ : BFR
      port map(A => \I2.N_2358_tz_tz\, Y => 
        \I2.N_2358_tz_tz_adt_net_854952__net_1\);
    
    \I2.BNC_IDl0r\ : DFFB
      port map(CLK => CLK_c, D => \I2.BNC_ID_i_0l0r\, CLR => 
        \I2.N_4621_i_0\, SET => \I2.N_4605_i_0\, Q => 
        \I2.BNC_IDl0r_net_1\);
    
    FID_padl31r : OB33PH
      port map(PAD => FID(31), A => FID_cl31r);
    
    \I2.PIPE5_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_688_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl12r_net_1\);
    
    \I3.VAS_64\ : MUX2L
      port map(A => VAD_inl2r, B => \I3.VASl2r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_64_net_1\);
    
    \I2.PIPE3_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl21r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl21r_net_1\);
    
    \I2.EVNT_NUMl1r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_962_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl1r_net_1\);
    
    \I1.sstatel9r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl1r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel9r_net_1\);
    
    \I5.SCL\ : DFFS
      port map(CLK => CLK_c, D => \I5.SCL_63_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SCL_net_1\);
    
    \I3.VADm_0_a3l6r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl6r_net_1\, Y => \I3.VADml6r\);
    
    \I3.PIPEB_86_2337\ : NOR2FT
      port map(A => \I3.PIPEBl7r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_86_adt_net_160419_\);
    
    \I2.BNCID_VECTROR_9_TZ_1418\ : AND2
      port map(A => \I2.BNCID_VECTra15_1_net_1\, B => 
        \I2.BNCID_VECTro_15\, Y => 
        \I2.BNCID_VECTror_9_tz_adt_net_48091_\);
    
    \I3.REG_1_157\ : MUX2L
      port map(A => VDB_inl8r, B => REGl56r, S => 
        \I3.N_1935_adt_net_855328__net_1\, Y => \I3.REG_1_157_0\);
    
    \I2.PIPE6_DT_468\ : MUX2H
      port map(A => \I2.PIPE5_DTl14r_net_1\, B => 
        \I2.PIPE6_DTl14r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_468_net_1\);
    
    \I1.REG_1_84\ : MUX2H
      port map(A => \REGl183r\, B => \I1.REG_74l183r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\, Y => 
        \I1.REG_1_84_net_1\);
    
    \I3.VDBi_57_iv_0_0_a2_10l7r_741\ : OR2FT
      port map(A => \I3.N_2016\, B => \I3.REGMAPL14R_732\, Y => 
        \I3.N_2017_119\);
    
    \I3.PIPEA1_310\ : MUX2L
      port map(A => \I3.PIPEA1l12r_net_1\, B => 
        \I3.PIPEA1_12l12r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__253\, Y => 
        \I3.PIPEA1_310_net_1\);
    
    \I2.TOKENB_CNT_3_0_a3l1r\ : AND2
      port map(A => \I2.N_177\, B => \I2.I_10\, Y => 
        \I2.TOKENB_CNT_3l1r\);
    
    \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_1038_\ : OAI21TTF
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096__net_1\, B
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        C => \I2.FIRST_TDC_1_sqmuxa_net_1\, Y => 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_1038__net_1\);
    
    \I2.N_3887_adt_net_855068_\ : BFR
      port map(A => \I2.N_3887\, Y => 
        \I2.N_3887_adt_net_855068__net_1\);
    
    \I2.LSRAM_INl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_412_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl28r_net_1\);
    
    \I2.RAMADl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l10r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl10r);
    
    \I3.VDBOFFA_31_IV_0L2R_2588\ : AND2
      port map(A => \REGl263r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        Y => \I3.VDBoffa_31l2r_adt_net_164238_\);
    
    \I2.PIPE5_DT_687\ : MUX2L
      port map(A => \I2.PIPE5_DTl11r_net_1\, B => 
        \I2.PIPE5_DT_6l11r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_687_net_1\);
    
    \I2.PIPE1_DT_754\ : MUX2L
      port map(A => \I2.PIPE1_DTl27r_net_1\, B => 
        \I2.PIPE1_DT_42_1_iv_i_0l27r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854564__net_1\, 
        Y => \I2.PIPE1_DT_754_net_1\);
    
    \I2.START_GIRO\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.START_GIRO_451_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.START_GIRO_net_1\);
    
    \I1.REG_74_0_IVL335R_1881\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l335r_adt_net_117658_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I173_Y\ : XOR2
      port map(A => \I2.N_2360_tz_tz\, B => 
        \I2.ADD_21x21_fast_I173_Y_0\, Y => \I2.un27_pipe5_dt0l3r\);
    
    \I1.REG_74_0_IVL233R_1993\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_9_sqmuxa_adt_net_854724__net_1\, Y => 
        \I1.REG_74l233r_adt_net_127366_\);
    
    \I2.STATE3_NSL6R_1047\ : NOR2FT
      port map(A => \I2.STATE3l7r_net_1\, B => PULSEl3r, Y => 
        \I2.STATE3_nsl6r_adt_net_24857_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I164_Y\ : OA21FTF
      port map(A => \I2.I180_un1_Y_adt_net_240115_\, B => 
        \I2.N495_i_adt_net_207682_\, C => \I2.N308_0\, Y => 
        \I2.N495_i\);
    
    \I2.RAMDT4L5R_2810\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_138\);
    
    \I3.REG_1l162r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_210_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl162r\);
    
    \I2.PIPE8_DT_21l6r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl6r\, B => \I2.N_572\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l6r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL13R_1446\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855224__net_1\, B => 
        \I2.MIC_ERR_REGSl13r_net_1\, C => 
        \I2.PIPE1_DT_42l13r_adt_net_49209_\, Y => 
        \I2.PIPE1_DT_42l13r_adt_net_49210_\);
    
    \I3.STATE1l8r_1164\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl2r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL8R_426\);
    
    \I2.RAMDT4l6r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl6r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l6r_net_1\);
    
    \I3.VDBI_57_0_IVL30R_2141\ : AND2
      port map(A => \I3.PIPEAl30r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l30r_adt_net_138033_\);
    
    \I3.VDBI_57_0_IV_0L27R_2148\ : AND2
      port map(A => \I3.PIPEAl27r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l27r_adt_net_138433_\);
    
    \I2.OFFSETl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_562_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl2r_net_1\);
    
    \I3.VDBi_57_iv_0_0_a2_11l7r\ : AND2FT
      port map(A => \I3.N_2017_317\, B => 
        \I3.REGMAPl9r_adt_net_854328__net_1\, Y => \I3.N_2044\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I179_Y_2686\ : AND3
      port map(A => \I2.N516\, B => \I2.N504_adt_net_88887_\, C
         => \I2.N481_adt_net_423940_\, Y => 
        \I2.N481_adt_net_424217_\);
    
    \I3.VDBI_57_0_IV_0L18R_2176\ : AND2
      port map(A => \I3.PIPEAl18r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l18r_adt_net_139489_\);
    
    \I2.REG_1_n7\ : XOR2FT
      port map(A => \I2.N_3835_i_0\, B => \I2.REG_1_n7_0_net_1\, 
        Y => \I2.REG_1_n7_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL1R_1517\ : OAI21TTF
      port map(A => GA_cl1r, B => \I2.N_3238\, C => 
        \I2.PIPE1_DT_42l1r_adt_net_52043_\, Y => 
        \I2.PIPE1_DT_42l1r_adt_net_52044_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I143_Y\ : XOR2
      port map(A => \I2.N346_adt_net_4075__net_1\, B => 
        \I2.ADD_18x18_fast_I143_Y_0\, Y => \I2.SUB9_1l6r\);
    
    \I3.REG_1_296\ : MUX2L
      port map(A => VDB_inl14r, B => REGl115r, S => 
        \I3.N_318_adt_net_855884__net_1\, Y => \I3.REG_1_296_0\);
    
    REGl169r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_70_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl169r\);
    
    \I5.SENS_ADDR_6l2r\ : AND2
      port map(A => \I5.SENS_ADDR_1_sqmuxa_net_1\, B => \I5.I_14\, 
        Y => \I5.SENS_ADDR_6l2r_net_1\);
    
    \I2.FID_425\ : MUX2H
      port map(A => FID_cl9r, B => \I2.FID_7l9r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        Y => \I2.FID_425_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_2\ : AO21
      port map(A => \I2.N_128_adt_net_54290_\, B => 
        \I2.N_128_adt_net_54291_\, C => 
        \I2.N_107_ADT_NET_256840__384\, Y => \I2.N_128\);
    
    \I2.PIPE4_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl23r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl23r_net_1\);
    
    \I2.WPAGE_951\ : XOR2
      port map(A => \I2.WPAGEl12r_net_1\, B => 
        \I2.WPAGEe_adt_net_855060__net_1\, Y => 
        \I2.WPAGE_951_net_1\);
    
    \I3.RAMAD_VMEl17r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_41_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl17r);
    
    \I2.WPAGEe_adt_net_855056_\ : BFR
      port map(A => \I2.WPAGEe_adt_net_855060__net_1\, Y => 
        \I2.WPAGEe_adt_net_855056__net_1\);
    
    \I2.PIPE4_DT_I_IL1R_3085\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DT_I_IL1R_849\);
    
    \I2.PIPE1_DT_42_1_ivl16r\ : OR3
      port map(A => \I2.PIPE1_DT_42l16r_adt_net_47837_\, B => 
        \I2.PIPE1_DT_42l16r_adt_net_47851_\, C => 
        \I2.PIPE1_DT_42l16r_adt_net_47852_\, Y => 
        \I2.PIPE1_DT_42l16r\);
    
    \I1.REG_74_0_ivl222r\ : AO21
      port map(A => \REGl222r\, B => \I1.N_97\, C => 
        \I1.REG_74l222r_adt_net_128480_\, Y => \I1.REG_74l222r\);
    
    \I2.un21_pipe5_dt_0_0\ : XOR2
      port map(A => \I2.RAMDT4L5R_815\, B => 
        \I2.un21_pipe5_dt_4_net_1\, Y => \I2.dataout_0\);
    
    REGl325r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_226_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl325r\);
    
    \I2.PIPE4_DTl8r_adt_net_854556__adt_net_855024_\ : BFR
      port map(A => \I2.PIPE4_DTl8r_adt_net_854556__net_1\, Y => 
        \I2.PIPE4_DTl8r_adt_net_854556__adt_net_855024__net_1\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044_\ : BFR
      port map(A => \I2.PIPE1_DT_2_SQMUXA_ADT_NET_803__299\, Y
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044__net_1\);
    
    \I2.DTE_21_1_ivl14r\ : AO21
      port map(A => \I2.DTE_1l14r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.DTE_21_1l14r_adt_net_38071_\, Y => \I2.DTE_21_1l14r\);
    
    \I2.DTO_16_1_iv_0l17r\ : OR2
      port map(A => \I2.DTO_16_1l17r_adt_net_31531_\, B => 
        \I2.DTO_16_1l17r_adt_net_31532_\, Y => \I2.DTO_16_1l17r\);
    
    \I2.BITCNT_n3_i_a5\ : NOR2
      port map(A => \I2.N_4328\, B => \I2.BITCNTl3r_net_1\, Y => 
        \I2.N_4336\);
    
    FID_padl19r : OB33PH
      port map(PAD => FID(19), A => FID_cl19r);
    
    \I2.PIPE8_DT_16_0l4r\ : MUX2H
      port map(A => \I2.PIPE8_DTl4r_net_1\, B => 
        \I2.PIPE7_DTl4r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_570\);
    
    \I2.EVNT_NUM_101\ : NAND3FTT
      port map(A => EV_RES_c, B => \I2.EVNT_NUMl10r_net_1\, C => 
        \I2.EVNT_NUM_c9_net_1\, Y => \I2.N_1232\);
    
    \I1.REG_74_0_ivl172r\ : AO21
      port map(A => \REGl172r\, B => \I1.N_41\, C => 
        \I1.REG_74l172r_adt_net_133063_\, Y => 
        \I1.REG_74l172r_net_1\);
    
    \I2.DTOSl2r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl2r, Q => 
        \I2.DTOSl2r_net_1\);
    
    \I2.REG_1_n12_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => REGl44r, Y => \I2.REG_1_n12_0_net_1\);
    
    \I2.DTO_cl_63_871\ : MUX2L
      port map(A => \I2.DTO_cl_32l31r\, B => \I2.N_2836\, S => 
        \I2.un1_DTO_cl_0_sqmuxa\, Y => \I2.DTO_cl_63_871_net_1\);
    
    \I3.VDBI_29L4R_2721\ : OA21
      port map(A => \I3.VDBi_13l4r_adt_net_284333_\, B => 
        \I3.VDBi_13l4r_adt_net_284335_\, C => 
        \I3.VDBi_29l4r_adt_net_621825_\, Y => 
        \I3.VDBi_29l4r_adt_net_621921_\);
    
    \I3.STATE1l4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl6r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl4r\);
    
    REGl247r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_148_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl247r\);
    
    \I3.MAJORITY_0_REG_5_I_IL0R_1540\ : OA21
      port map(A => \I3.REG2l0r_net_1\, B => \I3.REG3L0R_745\, C
         => \I3.REG1l0r_net_1\, Y => \REGl0r_adt_net_53773_\);
    
    \I1.REG_74_0_IV_0_0L253R_1972\ : AND2
      port map(A => \FBOUTl0r\, B => \I1.N_596\, Y => 
        \I1.REG_74l253r_adt_net_125400_\);
    
    \I1.REG_1_90\ : MUX2H
      port map(A => \REGl189r\, B => \I1.REG_74l189r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, Y => 
        \I1.REG_1_90_net_1\);
    
    \I3.REGMAPl29r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un126_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPl29r_net_1\);
    
    \I2.PIPE6_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_468_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl14r_net_1\);
    
    \I2.N_4667_1_ADT_NET_1046__2756\ : OAI21FTF
      port map(A => \I2.N_4261\, B => \I2.N_4283_I_0_42\, C => 
        \I2.STATE2L2R_589\, Y => \I2.N_4667_1_ADT_NET_1046__32\);
    
    \I3.VDBI_57_0_IV_0_0L8R_2225\ : AO21
      port map(A => \I3.N_2034_adt_net_854684__net_1\, B => 
        \I3.RAMDTSl8r_net_1\, C => 
        \I3.VDBi_57l8r_adt_net_142780_\, Y => 
        \I3.VDBi_57l8r_adt_net_142792_\);
    
    \I2.PIPE7_DTl25r_1576\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL25R_683\);
    
    \I2.PIPE3_DTl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl26r_net_1\);
    
    \I2.L2SERVl3r_1258\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_520\);
    
    \I2.DTO_1_905\ : MUX2L
      port map(A => \I2.DTO_1l31r_net_1\, B => \I2.DTO_16_1l31r\, 
        S => \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => 
        \I2.DTO_1_905_net_1\);
    
    \I3.REG_1l59r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_160_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl59r);
    
    \I2.STATE5L2R_3009\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE5_ns_il1r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.STATE5L2R_763\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_2_756\ : AO21
      port map(A => \I2.N_128_adt_net_54290_\, B => 
        \I2.N_128_adt_net_54291__adt_net_854408__net_1\, C => 
        \I2.N_107_adt_net_256840_\, Y => \I2.N_128_134\);
    
    \I2.DTO_1l15r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l15r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l15r_Rd1__net_1\);
    
    \I2.CRC32l31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_826_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l31r_net_1\);
    
    \I3.REG_1l61r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_162_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl61r);
    
    \I2.OFFSET_37_21l6r\ : MUX2L
      port map(A => \I2.N_793\, B => \I2.N_769\, S => 
        \I2.PIPE7_DTL25R_684\, Y => \I2.N_801\);
    
    \I2.un28_sram_empty_12_0\ : MUX2L
      port map(A => \I2.L2TYPEL15R_664\, B => \I2.L2TYPEL7R_663\, 
        S => \I2.RPAGEL15R_521\, Y => \I2.N_631\);
    
    \I3.VDBi_57_0_iv_0_0_a2l8r\ : NOR2
      port map(A => \I3.N_2015_120\, B => \I3.REGMAPL55R_781\, Y
         => \I3.N_2016\);
    
    \I3.REG3_125\ : MUX2L
      port map(A => VDB_inl0r, B => \I3.REG3l0r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855624__net_1\, Y => 
        \I3.REG3_125_net_1\);
    
    \I1.REG_74_0_IVL403R_1786\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_30_sqmuxa_adt_net_854372__net_1\, Y => 
        \I1.REG_74l403r_adt_net_109842_\);
    
    \I2.REG_1_c9_i_o2\ : NOR2FT
      port map(A => REGl41r, B => \I2.N_3852\, Y => \I2.N_3853\);
    
    \I1.un1_sbyte13_1_i_1_adt_net_106369__adt_net_854528_\ : BFR
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_106369_\, Y => 
        \I1.un1_sbyte13_1_i_1_adt_net_106369__adt_net_854528__net_1\);
    
    \I3.VDBI_57_IV_0L5R_2247\ : AO21
      port map(A => \I3.PIPEAl5r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l5r_adt_net_143850_\, Y => 
        \I3.VDBi_57l5r_adt_net_143861_\);
    
    \I3.UN1_REGMAP_30_0_A2_2084\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_134453_\, B => 
        \I3.N_58_i_0\, Y => \I3.un1_REGMAP_30_adt_net_134454_\);
    
    \I2.PIPE5_DT_6l15r\ : MUX2L
      port map(A => \I2.PIPE4_DTl15r_net_1\, B => \I2.N_1084\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\, Y
         => \I2.PIPE5_DT_6l15r_net_1\);
    
    \I3.TCNT4_n3\ : XOR2FT
      port map(A => \I3.TCNT4l3r_net_1\, B => \I3.TCNT4_c2_net_1\, 
        Y => \I3.TCNT4_n3_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I46_Y\ : OA21
      port map(A => \I2.N_3537_i_i\, B => 
        \I2.N311_adt_net_69399_\, C => \I2.G_1_3\, Y => \I2.N311\);
    
    \I2.PIPE9_DT_275\ : MUX2L
      port map(A => \I2.PIPE9_DTl6r_net_1\, B => 
        \I2.PIPE8_DTl6r_net_1\, S => \I2.NWPIPE8_i_0_i_0_0\, Y
         => \I2.PIPE9_DT_275_net_1\);
    
    FID_padl1r : OB33PH
      port map(PAD => FID(1), A => FID_cl1r);
    
    \I2.un9_clear_stat\ : OR2FT
      port map(A => CLEAR_STAT_12, B => \I2.CHAINA_ERRS_net_1\, Y
         => \I2.un9_clear_stat_i\);
    
    \I2.MIC_ERR_REGSl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_338_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl9r_net_1\);
    
    \I1.REG_74_0_IV_0_0_A2L253R_1963\ : NOR3FTT
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        B => \I1.PAGECNTl7r_net_1\, C => 
        \I1.N_268_Rd1__adt_net_854800__net_1\, Y => 
        \I1.N_596_adt_net_124704_\);
    
    \I3.VDBOFFB_30_IV_0L1R_2463\ : AO21
      port map(A => \REGl398r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l1r_adt_net_162884_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162928_\);
    
    \I2.PIPE4_DT_i_il1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DT_i_il1r_net_1\);
    
    \I3.VDBI_57_0_IVL23R_2160\ : AO21
      port map(A => \I3.VDBil23r_net_1\, B => 
        \I3.N_1910_0_adt_net_854344__net_1\, C => 
        \I3.VDBi_57l23r_adt_net_138945_\, Y => 
        \I3.VDBi_57l23r_adt_net_138951_\);
    
    \I2.PIPE8_DT_16l13r\ : AND2
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\, B => 
        \I2.N_579\, Y => \I2.PIPE8_DT_16l13r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL8R_1477\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\, B => 
        \I2.PIPE1_DT_30l8r_net_1\, C => 
        \I2.PIPE1_DT_42l8r_adt_net_50430_\, Y => 
        \I2.PIPE1_DT_42l8r_adt_net_50446_\);
    
    \I2.FID_7_0_ivl0r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl0r_net_1\, 
        C => \I2.FID_7l0r_adt_net_93577_\, Y => \I2.FID_7l0r\);
    
    \I2.L2TYPE_4_IL4R_1634\ : NAND2
      port map(A => \I2.N_4458\, B => \I2.N_4460\, Y => 
        \I2.N_4448_adt_net_68212_\);
    
    \I3.VDBOFFB_30_IV_0L1R_2457\ : AND2
      port map(A => \REGl350r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162888_\);
    
    \I2.PIPE8_DT_16_0l10r\ : MUX2H
      port map(A => \I2.PIPE8_DTl10r_net_1\, B => 
        \I2.PIPE7_DTl10r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_576\);
    
    \I2.DTE_21_1_IV_0L20R_1262\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l20r\, C
         => \I2.DTE_21_1l20r_adt_net_37614_\, Y => 
        \I2.DTE_21_1l20r_adt_net_37615_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I153_Y_i\ : NAND3
      port map(A => \I2.N_20_i_0\, B => \I2.N_33_0\, C => 
        \I2.N_86_i_0\, Y => \I2.N_2_0\);
    
    \I3.VASl9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_71_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl9r_net_1\);
    
    \I2.N507_adt_net_258084_\ : AND3FFT
      port map(A => \I2.N_74_i_0_i_adt_net_54331_\, B => 
        \I2.N_80\, C => \I2.N507_adt_net_56251__net_1\, Y => 
        \I2.N507_adt_net_258084__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I183_Y\ : XOR2FT
      port map(A => \I2.N513_i_0\, B => 
        \I2.ADD_21x21_fast_I183_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l13r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I139_Y_i\ : NAND2
      port map(A => \I2.N_91\, B => \I2.N_96\, Y => \I2.N_42_0\);
    
    DPR_padl27r : IB33
      port map(PAD => DPR(27), Y => DPR_cl27r);
    
    \I1.RAMDT_SPI_1l3r\ : DFFC
      port map(CLK => CLK_c, D => \FBOUTl3r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.RAMDT_SPI_1l3r_net_1\);
    
    \I1.sstate_ns_i_0l0r\ : AOI21TTF
      port map(A => \I1.N_628\, B => \I1.sstate_ns_i_0_a4_0_1l0r\, 
        C => \I1.N_292\, Y => \I1.N_43_i_0\);
    
    \I2.OFFSET_37_22l2r\ : MUX2L
      port map(A => \REGl239r\, B => \REGl175r\, S => 
        \I2.PIPE7_DTL27R_83\, Y => \I2.N_805\);
    
    \I3.STATE1_TR24_I_0_O2_1_0_2110\ : AND3FFT
      port map(A => \I3.REGMAPl47r_net_1\, B => 
        \I3.REGMAP_i_il46r_net_1\, C => 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135383_\, Y => 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135385_\);
    
    \I3.PIPEA_234\ : MUX2L
      port map(A => \I3.PIPEAl3r_net_1\, B => 
        \I3.PIPEA_8l3r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854680__net_1\, Y
         => \I3.PIPEA_234_net_1\);
    
    \I2.DTO_16_1_iv_0_o2_0l6r\ : OAI21FTT
      port map(A => \I2.STATE2l4r_net_1\, B => 
        \I2.N_4283_I_0_234\, C => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\, Y => 
        \I2.N_4671\);
    
    \I1.REG_1_220\ : MUX2H
      port map(A => \REGl319r\, B => \I1.REG_74l319r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_220_net_1\);
    
    \I2.ROFFSETl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_906_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl12r_net_1\);
    
    \I1.REG_74_0_iv_0l371r\ : AO21
      port map(A => \REGl371r\, B => \I1.N_660\, C => 
        \I1.REG_74l371r_adt_net_113396_\, Y => \I1.REG_74l371r\);
    
    DPR_padl5r : IB33
      port map(PAD => DPR(5), Y => DPR_cl5r);
    
    \I3.TCNT2l7r\ : DFFC
      port map(CLK => CLK_c, D => TCNT2_389, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT2l7r_net_1\);
    
    \I1.REG_74_0_IVL175R_2059\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, Y => 
        \I1.REG_74l175r_adt_net_132768_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I180_Y\ : XOR2FT
      port map(A => \I2.N522\, B => \I2.ADD_21x21_fast_I180_Y_0\, 
        Y => \I2.un27_pipe5_dt0l10r\);
    
    \I1.REG_74_0_ivl175r\ : AO21
      port map(A => \REGl175r\, B => \I1.N_49\, C => 
        \I1.REG_74l175r_adt_net_132768_\, Y => \I1.REG_74l175r\);
    
    \I2.FID_7_0_IVL27R_982\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl75r, C => 
        \I2.FID_7l27r_adt_net_18833_\, Y => 
        \I2.FID_7l27r_adt_net_18841_\);
    
    \I2.SRAM_EVNT_n3_0\ : XOR2FT
      port map(A => \I2.SRAM_EVNTl3r_net_1\, B => \I2.N_128_1\, Y
         => \I2.SRAM_EVNT_n3_0_net_1\);
    
    \I2.DTE_1l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_842_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l2r_net_1\);
    
    \I3.VADm_0_a3l29r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl29r_net_1\, Y => \I3.VADml29r\);
    
    \I3.REGMAPl17r_adt_net_854280_\ : BFR
      port map(A => \I3.REGMAPl17r_adt_net_854288__net_1\, Y => 
        \I3.REGMAPl17r_adt_net_854280__net_1\);
    
    \I3.SINGCYC_115\ : MUX2H
      port map(A => \I3.SINGCYC_881\, B => 
        \I3.un7_cycs_0_a3_0_a3_net_1\, S => \I3.N_1510\, Y => 
        \I3.SINGCYC_115_net_1\);
    
    \I2.un1_TOKENA_CNT_I_10\ : XOR2
      port map(A => \I2.TOKENA_CNTl1r_net_1\, B => 
        \I2.DWACT_ADD_CI_0_TMP_2l0r\, Y => \I2.I_10_0\);
    
    \I2.CRC32_12_i_0_m2l17r\ : MUX2L
      port map(A => \I2.DT_TEMPl17r_net_1\, B => \I2.N_188\, S
         => \I2.N_4667_1_adt_net_1046__adt_net_854196__net_1\, Y
         => \I2.N_224_i_i\);
    
    \I2.PIPE4_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl25r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I185_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_801\, B => 
        \I2.PIPE4_DTl15r_net_1\, Y => 
        \I2.ADD_21x21_fast_I185_Y_0_0\);
    
    \I2.DT_TEMPl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_766_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl5r_net_1\);
    
    \I3.PIPEAl31r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_262_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl31r_net_1\);
    
    \I2.ROFFSET_c4\ : NOR2FT
      port map(A => \I2.ROFFSETL4R_874\, B => 
        \I2.ROFFSET_c3_net_1\, Y => \I2.ROFFSET_c4_net_1\);
    
    REGl166r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_67_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl166r\);
    
    REGl223r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_124_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl223r\);
    
    \I1.REG_74_0_ivl313r\ : AO21
      port map(A => \REGl313r\, B => \I1.N_185\, C => 
        \I1.REG_74l313r_adt_net_119647_\, Y => \I1.REG_74l313r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I5_P0N_i_a4_732\ : OR2
      port map(A => \I2.RAMDT4L12R_141\, B => 
        \I2.PIPE4_DTl5r_adt_net_854416__net_1\, Y => 
        \I2.N_89_0_110\);
    
    \I2.REG_1l46r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n14_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl46r);
    
    \I3.un1_STATE1_8_i\ : AO21FTT
      port map(A => \I3.STATE1_ipl8r\, B => \I3.STATE1_IPL9R_11\, 
        C => \I3.N_1906_i_0_0_adt_net_855640__net_1\, Y => 
        \I3.N_127\);
    
    \I3.PIPEA_8l27r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854456__net_1\, B => 
        \I3.N_236\, Y => \I3.PIPEA_8l27r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I150_Y_0\ : XOR2FT
      port map(A => \I2.SUB8l14r_adt_net_855568__net_1\, B => 
        \I2.SUB8l13r_adt_net_855564__net_1\, Y => 
        \I2.ADD_18x18_fast_I150_Y_0\);
    
    \I2.REG_1_c4_i\ : AND2FT
      port map(A => \I2.N_124\, B => 
        \I2.N_3834_i_0_adt_net_1384__net_1\, Y => \I2.N_3833_i_0\);
    
    \I2.UN1_END_EVNT1_0_SQMUXA_I_0_1007\ : AO21FTF
      port map(A => \I2.N_3877_adt_net_855268__net_1\, B => 
        \I2.STATE1L18R_875\, C => \I2.N_3888\, Y => 
        \I2.N_3234_adt_net_21449_\);
    
    \I2.TRAIL_MIS6_i\ : INV
      port map(A => \I2.TRAIL_MIS6_net_1\, Y => 
        \I2.TRAIL_MIS6_i_net_1\);
    
    \I2.DTO_16_1_IVL14R_1148\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.N_126_i_0\, Y => 
        \I2.DTO_16_1l14r_adt_net_32202_\);
    
    RAMAD_padl1r : OB33PH
      port map(PAD => RAMAD(1), A => RAMAD_cl1r);
    
    \I2.G_EVNT_NUM_n3_i_0\ : NOR3
      port map(A => EV_RES_C_569, B => \I2.N_317\, C => 
        \I2.N_189\, Y => \I2.N_4343\);
    
    \I2.WREi\ : DFFS
      port map(CLK => CLK_c, D => \I2.WREi_794_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.WREi_net_1\);
    
    \I1.REG_74_24_404_m8_i_x2\ : XOR2
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        B => \I1.REG_74_24_404_m3_e_net_1\, Y => 
        \I1.REG_74_24_404_N_6_i_i\);
    
    \I3.VDBml21r\ : MUX2L
      port map(A => \I3.VDBil21r_net_1\, B => \I3.N_163\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml21r_net_1\);
    
    \I2.PIPE7_DTl33r\ : DFFS
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_il33r_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DT_i_0l33r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I42_Y\ : AND2
      port map(A => \I2.G_1_1\, B => \I2.N307_1_adt_net_69278_\, 
        Y => \I2.N307_1\);
    
    \I2.DT_SRAM_i_1_m2l2r_999\ : MUX2L
      port map(A => \I2.N_4191\, B => \I2.PIPE2_DTl2r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.N_4193_377\);
    
    REGl267r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_168_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl267r\);
    
    \I1.REG_1_223\ : MUX2H
      port map(A => \REGl322r\, B => \I1.REG_74l322r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y => 
        \I1.REG_1_223_net_1\);
    
    WMIC_pad : OB33PH
      port map(PAD => WMIC, A => WMIC_c);
    
    \I3.VADm_0_a3l21r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl21r_net_1\, Y => \I3.VADml21r\);
    
    \I2.CRC32_12_0_0_x3l18r\ : XOR2FT
      port map(A => \I2.CRC32l18r_net_1\, B => \I2.N_4096_i_i\, Y
         => \I2.N_52_i_0_i_0\);
    
    \I2.ROFFSETl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_914_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl4r_net_1\);
    
    \I2.RAMAD1_665\ : MUX2L
      port map(A => \I2.RAMAD1_12l11r_net_1\, B => 
        \I2.RAMAD1l11r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__171\, Y => 
        \I2.RAMAD1_665_net_1\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__2768\ : NAND3FFT
      port map(A => \I2.ENDF_618\, B => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149__net_1\, C => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_61\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__57\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I162_Y\ : AND2FT
      port map(A => \I2.I162_un1_Y\, B => 
        \I2.N489_i_adt_net_89351_\, Y => \I2.N489_i\);
    
    \I2.DTE_21_1_IV_0L24R_1246\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855196__net_1\, 
        B => \I2.DT_TEMPl24r_net_1\, C => 
        \I2.DTO_16_1l24r_adt_net_29860_\, Y => 
        \I2.DTE_21_1l24r_adt_net_37173_\);
    
    \I3.PIPEBl20r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_99_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl20r_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_A2_1_1_1542\ : 
        NAND2FT
      port map(A => \I2.N_107_adt_net_276024_\, B => \I2.N_17\, Y
         => \I2.N_108_adt_net_54237_\);
    
    \I3.STATE2l2r_1614\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE2l3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.STATE2L2R_721\);
    
    \I2.TRGARR_3_I_18\ : XOR2
      port map(A => \I2.DWACT_ADD_CI_0_g_array_1l0r\, B => 
        \I2.TRGARRl2r_net_1\, Y => \I2.TRGARR_3l2r\);
    
    \I2.LEAD_FLAG6l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_641_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl4r);
    
    DPR_padl22r : IB33
      port map(PAD => DPR(22), Y => DPR_cl22r);
    
    \I1.N_606_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_606_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_606_Rd1__net_1\);
    
    \I2.PIPE1_DT_30l0r\ : MUX2H
      port map(A => \I2.TDCDBSl19r_net_1\, B => 
        \I2.TDCDBSl0r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, Y
         => \I2.PIPE1_DT_30l0r_net_1\);
    
    \I2.CRC32_12_i_0l19r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_247_i_i_0\, Y => 
        \I2.N_3936\);
    
    \I1.N_50_0_adt_net_109757_\ : NOR3
      port map(A => \I1.BYTECNTl3r_net_1\, B => 
        \I1.BYTECNT_i_0_il1r_net_1\, C => 
        \I1.N_311_i_i_Rd1__adt_net_854920__net_1\, Y => 
        \I1.N_50_0_adt_net_109757__net_1\);
    
    \I1.PAGECNT_0l7r_adt_net_835112_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_320_adt_net_854876__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__net_1\);
    
    \I1.PAGECNT_n6_i_i\ : AO21FTF
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_854524__net_1\, 
        B => \I1.N_1377_adt_net_1517__net_1\, C => \I1.N_473_206\, 
        Y => \I1.N_1377\);
    
    \I2.STATE1l10r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3206_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1l10r_net_1\);
    
    \I1.REG_1_272\ : MUX2H
      port map(A => \REGl371r\, B => \I1.REG_74l371r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_272_net_1\);
    
    \I3.un12_tcnt3\ : AND3FTT
      port map(A => \I3.un10_tcnt2_net_1\, B => 
        \I3.un12_tcnt3_adt_net_165620_\, C => 
        \I3.un12_tcnt3_adt_net_165621_\, Y => 
        \I3.un12_tcnt3_net_1\);
    
    \I2.un1_tdc_res_29_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl408r, Y => 
        \I2.N_4610_i_0\);
    
    \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L3R_2581\ : OR3
      port map(A => \I3.VDBoffa_31l3r_adt_net_164077_\, B => 
        \I3.VDBoffa_31l3r_adt_net_164073_\, C => 
        \I3.VDBoffa_31l3r_adt_net_164074_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164080_\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I120_Y_0_78_TZ_TZ_1548\ : 
        AND2
      port map(A => \I2.RAMDT4L2R_767\, B => \I2.PIPE4_DTL2R_860\, 
        Y => \I2.N_2360_tz_tz_adt_net_54584_\);
    
    \I2.REG_1l47r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n15_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl47r);
    
    \I2.TOKENA_CNT_i_0l1r\ : NAND2
      port map(A => CLEAR_STAT_12, B => \I2.TOKENTOA_RES_net_1\, 
        Y => \I2.un6_clear_stat_i\);
    
    \I2.EVNT_NUM_956\ : MUX2L
      port map(A => \I2.EVNT_NUMl7r_net_1\, B => 
        \I2.EVNT_NUM_n7_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_956_net_1\);
    
    \I3.TCNTl3r_1772\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_381_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTL3R_878\);
    
    \I2.DTO_16_1_IV_0L7R_1187\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854624__net_1\, 
        B => \I2.DT_TEMPl7r_net_1\, C => 
        \I2.DTO_16_1l7r_adt_net_33728_\, Y => 
        \I2.DTO_16_1l7r_adt_net_33734_\);
    
    \I1.BITCNT_n1_i_i_m4\ : AO21TTF
      port map(A => \I1.N_1376_i_0\, B => \I1.N_387_i_0\, C => 
        \I1.N_604\, Y => \I1.N_416\);
    
    \I2.ROFFSET_n8_tz\ : XOR2
      port map(A => \I2.ROFFSETl8r_net_1\, B => 
        \I2.ROFFSET_c7_net_1\, Y => \I2.ROFFSET_n8_tz_i\);
    
    \I2.DTO_1l4r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l4r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l4r_Rd1__net_1\);
    
    \I1.REG_1_274\ : MUX2H
      port map(A => \REGl373r\, B => \I1.REG_74l373r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_274_net_1\);
    
    \I2.DT_SRAMl15r\ : MUX2L
      port map(A => \I2.N_883\, B => \I2.PIPE2_DTl15r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668__net_1\, 
        Y => \I2.DT_SRAMl15r_net_1\);
    
    \I2.G_EVNT_NUM_n4_i_0\ : AND2
      port map(A => \I2.N_4669_adt_net_855052__net_1\, B => 
        \I2.N_4344_adt_net_26298_\, Y => \I2.N_4344\);
    
    \I2.SUB8_523_2743\ : OR3
      port map(A => \I2.SUB8_523_adt_net_670059_\, B => 
        \I2.SUB8_523_adt_net_670064_\, C => 
        \I2.SUB8_523_adt_net_670055_\, Y => \I2.SUB8_523_net_1\);
    
    \I2.N_3279_0_adt_net_855224_\ : BFR
      port map(A => \I2.N_3279_0_adt_net_855236__net_1\, Y => 
        \I2.N_3279_0_adt_net_855224__net_1\);
    
    \I2.L2TYPE_595\ : MUX2L
      port map(A => \I2.L2TYPEl6r_net_1\, B => \I2.N_4446\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_595_net_1\);
    
    \I1.REG_1_295\ : MUX2H
      port map(A => \REGl394r\, B => \I1.REG_74l394r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y => 
        \I1.REG_1_295_net_1\);
    
    \I2.un1_STATE3_3_0\ : OR2
      port map(A => \I2.STATE3l5r_net_1\, B => 
        \I2.STATE3l13r_net_1\, Y => \I2.un1_STATE3_3\);
    
    \I3.PIPEA1l21r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_319_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l21r_net_1\);
    
    \I1.REG_74_0_ivl309r\ : AO21
      port map(A => \REGl309r\, B => \I1.N_185\, C => 
        \I1.REG_74l309r_adt_net_119991_\, Y => \I1.REG_74l309r\);
    
    \I0.COM_SERSi\ : DFFC
      port map(CLK => CLK_c, D => \I0.COM_SERF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => COM_SERS);
    
    \I2.DTE_21_1_iv_0l27r\ : AO21
      port map(A => \I2.DTE_1l27r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.DTE_21_1l27r_adt_net_36861_\, Y => \I2.DTE_21_1l27r\);
    
    \I3.RAMAD_VME_30\ : MUX2H
      port map(A => RAMAD_VMEl6r, B => \I3.VAS_i_0_il7r\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_30_net_1\);
    
    \I2.MIC_ERR_REGS_373\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl45r_net_1\, B => 
        \I2.MIC_ERR_REGSl44r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_373_net_1\);
    
    \I2.MIC_ERR_REGS_358\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl30r_net_1\, B => 
        \I2.MIC_ERR_REGSl29r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_358_net_1\);
    
    \I2.STATEe_ns_a3l2r\ : OA21TTF
      port map(A => \I2.STATEe_ipl1r\, B => 
        \I2.N_3496_adt_net_926__net_1\, C => 
        \I2.CHAIN_ERRS_net_1\, Y => \I2.STATEe_nsl2r\);
    
    \I3.STATE1_ipl0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_ipl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl0r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I103_Y\ : AOI21
      port map(A => \I2.N318\, B => \I2.N315\, C => \I2.N314\, Y
         => \I2.N357_1\);
    
    \I2.CRC32_12_i_0l27r\ : NOR2
      port map(A => \I2.N_2867_1_adt_net_854964__net_1\, B => 
        \I2.N_246_i_i_0\, Y => \I2.N_3944\);
    
    \I2.DT_SRAM_0l6r\ : MUX2L
      port map(A => \I2.PIPE10_DTl6r_net_1\, B => 
        \I2.PIPE5_DTl6r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854224__net_1\, Y => 
        \I2.N_874\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I176_Y\ : XOR2FT
      port map(A => \I2.N_31_0\, B => 
        \I2.ADD_21x21_fast_I176_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l6r\);
    
    \I3.REGMAP_I_IL46R_2930\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un211_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_IL46R_447\);
    
    \I2.TDC_652\ : MUX2H
      port map(A => \I2.TDCl2r_net_1\, B => 
        \I2.RAMAD1_12l15r_net_1\, S => 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_1038__net_1\, Y => 
        \I2.TDC_652_net_1\);
    
    \I5.SSTATE1SE_13_0_900\ : AOI21TTF
      port map(A => TICKL0R_557, B => \I5.PULSE_FL_net_1\, C => 
        \I5.sstate1l13r_net_1\, Y => 
        \I5.sstate1_ns_el0r_adt_net_8036_\);
    
    \I1.REG_74_0_IVL280R_1939\ : NOR2FT
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l280r_adt_net_122721_\);
    
    \I2.CRC32_12_0_0_m2l26r\ : MUX2L
      port map(A => \I2.DT_TEMPl26r_net_1\, B => 
        \I2.DT_SRAMl26r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854192__net_1\, Y => 
        \I2.N_4271_i_i\);
    
    \I2.RAMDT4L12R_3040\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_794\);
    
    \I3.VDBOFFA_31_IV_0L4R_2560\ : AO21
      port map(A => \REGl185r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.VDBoffa_31l4r_adt_net_163878_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163885_\);
    
    \I3.VDBml12r\ : MUX2L
      port map(A => \I3.VDBil12r_net_1\, B => \I3.N_154\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml12r_net_1\);
    
    \I3.TCNT3_374\ : MUX2H
      port map(A => \I3.TCNT3l5r_net_1\, B => \I3.TCNT3_n5_net_1\, 
        S => \TICKl1r\, Y => \I3.TCNT3_374_net_1\);
    
    \I3.VASl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_64_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl2r_net_1\);
    
    \I1.REG_74_0_iv_i_a2l210r\ : AO21
      port map(A => \REGl210r\, B => \I1.N_183_i_0\, C => 
        \I1.N_1349_adt_net_129673_\, Y => \I1.N_1349\);
    
    \I2.DTOSl25r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl25r, Q => 
        \I2.DTOSl25r_net_1\);
    
    \I2.BNC_IDl3r_1478\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_13_2\, CLR => 
        \I2.N_4624_i_0\, SET => \I2.N_4613_i_0\, Q => 
        \I2.BNC_IDL3R_585\);
    
    \I3.PIPEA1_328\ : MUX2L
      port map(A => \I3.PIPEA1l30r_net_1\, B => 
        \I3.PIPEA1_12l30r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, Y => 
        \I3.PIPEA1_328_net_1\);
    
    \I1.REG_74_11_a0l404r\ : NAND2
      port map(A => \I1.N_267\, B => \I1.N_260_222\, Y => 
        \I1.REG_74_11_a0l404r_net_1\);
    
    \I3.REG_1_I_IL2R_1006\ : OA21
      port map(A => \I3.REG3L2R_742\, B => \I3.REG2l2r_net_1\, C
         => \I3.REG1l2r_net_1\, Y => \REGl2r_adt_net_21315_\);
    
    \I3.STATE1_ILLEGAL_2134\ : AO21
      port map(A => \I3.STATE1_ipl1r\, B => \I3.N_1186\, C => 
        \I3.N_1193_ip_adt_net_136556_\, Y => 
        \I3.N_1193_ip_adt_net_136557_\);
    
    \I2.UN1_REG80_I_1698\ : NOR2
      port map(A => REGl37r, B => REGl47r, Y => 
        \I2.N_3824_adt_net_90289_\);
    
    \I3.REG2_141\ : MUX2L
      port map(A => VDB_inl0r, B => \I3.REG2l0r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG2_141_net_1\);
    
    \I2.END_CHAINB1_1487\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.END_CHAINB1_709_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.END_CHAINB1_594\);
    
    \I2.L_LUT_498\ : AO21FTT
      port map(A => \I2.STATE2l0r_net_1\, B => \I2.L_LUT_net_1\, 
        C => \I2.L_LUT_498_adt_net_90208_\, Y => 
        \I2.L_LUT_498_net_1\);
    
    \I2.un1_PIPE1_DT_0_sqmuxa_1_i_a3_i_a3\ : NOR2
      port map(A => \I2.END_CHAINA1_net_1\, B => \I2.N_3288\, Y
         => \I2.N_148\);
    
    \I2.PIPE1_DT_42_1_IVL6R_1484\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl22r_net_1\, Y => 
        \I2.PIPE1_DT_42l6r_adt_net_50920_\);
    
    \I2.PIPE10_DT_627\ : MUX2L
      port map(A => \I2.PIPE10_DTl22r_net_1\, B => 
        \I2.PIPE9_DTl22r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_627_net_1\);
    
    \I2.PIPE1_DT_747\ : MUX2L
      port map(A => \I2.PIPE1_DTl20r_net_1\, B => 
        \I2.PIPE1_DT_42l20r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854568__net_1\, 
        Y => \I2.PIPE1_DT_747_net_1\);
    
    \I2.N411_adt_net_194931_\ : OR2FT
      port map(A => \I2.LSRAM_OUTl0r\, B => 
        \I2.PIPE7_DTl0r_net_1\, Y => 
        \I2.N411_adt_net_194931__net_1\);
    
    \I2.LSRAM_RADDRi_1_sqmuxa_0_a4_i_o2_45_tz\ : AO21FTT
      port map(A => LEAD_FLAGl3r, B => \I2.PIPE4_DTl21r_net_1\, C
         => \I2.N_2327_tz_adt_net_16395_\, Y => \I2.N_2327_tz\);
    
    \I2.FIDl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_435\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl19r);
    
    \I2.PIPE4_DTL10R_2958\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL10R_475\);
    
    \I3.VDBI_57_0_IVL25R_2154\ : AO21
      port map(A => \I3.VDBil25r_net_1\, B => 
        \I3.N_1910_0_adt_net_854344__net_1\, C => 
        \I3.VDBi_57l25r_adt_net_138707_\, Y => 
        \I3.VDBi_57l25r_adt_net_138713_\);
    
    \I2.LSRAM_INl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_407_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl23r_net_1\);
    
    REGl306r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_207_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl306r\);
    
    \I2.RAMAD_4_0l6r\ : MUX2H
      port map(A => \I2.RAMAD1l6r_net_1\, B => RAMAD_VMEl6r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_533\);
    
    \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840_\ : BFR
      port map(A => \I2.MIC_REG1_1_sqmuxa_0\, Y => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\);
    
    \I2.PIPE10_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_627_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl22r_net_1\);
    
    \I2.DT_TEMP_7l1r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, B => 
        \I2.DT_SRAMl1r_net_1\, Y => \I2.DT_TEMP_7l1r_net_1\);
    
    \I3.PULSE_46_0_iv_0_il1r\ : AO21
      port map(A => \I3.REGMAP_i_0_il5r\, B => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        C => PULSEl1r, Y => \I3.N_118_adt_net_147476_\);
    
    \I3.VDBi_57_iv_0_0_a2_10l7r_740\ : OR2FT
      port map(A => \I3.N_2016\, B => \I3.REGMAPl14r_net_1\, Y
         => \I3.N_2017_118\);
    
    \I1.REG_1_95\ : MUX2H
      port map(A => \REGl194r\, B => \I1.REG_74l194r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\, Y => 
        \I1.REG_1_95_net_1\);
    
    \I2.STATE2_NS_0L1R_1052\ : NOR3
      port map(A => NOESRAME_C_243, B => 
        \I2.WOFFSETl0r_adt_net_854636__net_1\, C => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, Y => 
        \I2.STATE2_nsl1r_adt_net_24965_\);
    
    \I3.PIPEA1l24r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_322_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l24r_net_1\);
    
    \I2.DTO_16_1_IV_0_0L16R_1136\ : AO21
      port map(A => \I2.G_EVNT_NUM_i_0_il0r_net_1\, B => 
        \I2.N_457\, C => \I2.DTO_16_1l16r_adt_net_31706_\, Y => 
        \I2.DTO_16_1l16r_adt_net_31717_\);
    
    \I2.DTO_16_1_IVL10R_1169\ : AND2
      port map(A => \I2.DTO_1l10r\, B => \I2.N_196_52\, Y => 
        \I2.DTO_16_1l10r_adt_net_33054_\);
    
    \I1.REG_74_0_iv_0l220r\ : AO21
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.REG_7_sqmuxa\, 
        C => \I1.REG_74l220r_adt_net_128776_\, Y => 
        \I1.REG_74l220r_net_1\);
    
    \I2.STATEe_i_0l0r\ : OR2FT
      port map(A => CLEAR_STAT_12, B => 
        \I2.STATEe_illegalpipe2_net_1\, Y => 
        \I2.STATEe_i_0l0r_net_1\);
    
    \I5.COMMAND_4l0r\ : MUX2L
      port map(A => \I5.AIR_WDATAl0r_net_1\, B => REGl101r, S => 
        REGl7r, Y => \I5.COMMAND_4l0r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I64_Y\ : AO21
      port map(A => \I2.N301_1\, B => \I2.N298\, C => \I2.N297\, 
        Y => \I2.N332\);
    
    \I5.COMMANDl14r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_51_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl14r_net_1\);
    
    \I2.RESYN_0_I2_LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_945\ : AO21
      port map(A => \I2.PIPE4_DTl22r_net_1\, B => \I2.N_2329_tz\, 
        C => \I2.N_4524_adt_net_16635_\, Y => 
        \I2.N_4524_adt_net_16596_\);
    
    \I1.REG_74_0_iv_0_o2_0l253r\ : OAI21TTF
      port map(A => \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, 
        B => 
        \I1.PAGECNT_0l7r_adt_net_835112_Rd1__adt_net_855516__net_1\, 
        C => \PULSE_0L0R_ADT_NET_834380_RD1__831\, Y => 
        \I1.REG_74_0_iv_0_o2_0_il253r\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_2_755\ : AO21
      port map(A => \I2.N_128_adt_net_54290_\, B => 
        \I2.N_128_adt_net_54291__adt_net_854408__net_1\, C => 
        \I2.N_107_adt_net_256840_\, Y => \I2.N_128_133\);
    
    \I3.PIPEA_8_0l18r\ : MUX2L
      port map(A => DPR_cl18r, B => \I3.PIPEA1l18r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855348__net_1\, Y => \I3.N_227\);
    
    \I1.REG_74_8_0_o4_0l380r_813\ : NAND2
      port map(A => \I1.N_1366\, B => \I1.N_1367_i\, Y => 
        \I1.N_396_191\);
    
    \I2.FID_421\ : MUX2H
      port map(A => FID_cl5r, B => \I2.FID_7_0_ivl5r_net_1\, S
         => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        Y => \I2.FID_421_net_1\);
    
    \I2.STATE1_NSL6R_1036\ : NOR2
      port map(A => TDCDRYA_c, B => \I2.STATE1_ns_1l7r\, Y => 
        \I2.STATE1_nsl6r_adt_net_23511_\);
    
    \I2.RAMAD_4_0l10r\ : MUX2H
      port map(A => \I2.RAMAD1l10r_net_1\, B => RAMAD_VMEl10r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_537\);
    
    \I3.un1_STATE1_13_1_adt_net_137896_\ : NOR3
      port map(A => \I3.STATE1_IPL9R_11\, B => \I3.STATE1_ipl7r\, 
        C => \I3.N_1910_0\, Y => 
        \I3.un1_STATE1_13_1_adt_net_137896__net_1\);
    
    \I2.FIDl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_427\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl11r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I180_Y\ : XOR2FT
      port map(A => \I2.N522_0\, B => 
        \I2.ADD_21x21_fast_I180_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l10r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I35_Y\ : AOI21FTF
      port map(A => \I2.SUB8l11r_net_1\, B => \I2.SUB8l12r_net_1\, 
        C => \I2.N247\, Y => \I2.N300\);
    
    \I1.REG_74_0_ivl174r\ : AO21
      port map(A => \REGl174r\, B => \I1.N_49\, C => 
        \I1.REG_74l174r_adt_net_132854_\, Y => \I1.REG_74l174r\);
    
    \I2.N_3_0_adt_net_1070_\ : AOI21
      port map(A => \I2.PIPE4_DTL6R_853\, B => 
        \I2.PIPE4_DTl7r_net_1\, C => \I2.RAMDT4L12R_142\, Y => 
        \I2.N_3_0_adt_net_1070__net_1\);
    
    \I2.PIPE10_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_606_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl1r_net_1\);
    
    \I5.SDANOE_8_0_914\ : NOR2
      port map(A => \I5.sstate1l9r_net_1\, B => 
        \I5.sstate1l11r_net_1\, Y => \I5.SDAnoe_8_adt_net_9736_\);
    
    \I2.N_2864_0_adt_net_854272_\ : BFR
      port map(A => \I2.N_2864_0\, Y => 
        \I2.N_2864_0_adt_net_854272__net_1\);
    
    \I3.VDBm_0l19r\ : MUX2L
      port map(A => \I3.PIPEAl19r_net_1\, B => 
        \I3.PIPEBl19r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_161\);
    
    \I3.CYCS1\ : DFFS
      port map(CLK => CLK_c, D => \I3.un7_cycs_i_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.CYCS1_i_0\);
    
    \I2.L2AS\ : AND2FT
      port map(A => \I2.L2AF3_net_1\, B => \I2.L2AF2_net_1\, Y
         => \I2.L2AS_net_1\);
    
    \I2.L2TYPE_591\ : MUX2L
      port map(A => \I2.L2TYPEl2r_net_1\, B => \I2.N_4450\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_591_net_1\);
    
    \I3.REG_1l75r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_176_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl75r);
    
    \I3.PIPEBl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_80_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl1r_net_1\);
    
    \I2.RAMDT4l4r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl4r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l4r_net_1\);
    
    \I2.OFFSET_37_10l1r\ : MUX2L
      port map(A => \I2.N_700\, B => \I2.N_692\, S => 
        \I2.PIPE7_DTL26R_355\, Y => \I2.N_708\);
    
    \I3.REG_1_163\ : MUX2L
      port map(A => VDB_inl14r, B => REGl62r, S => 
        \I3.N_1935_adt_net_855324__net_1\, Y => \I3.REG_1_163_0\);
    
    DPR_padl28r : IB33
      port map(PAD => DPR(28), Y => DPR_cl28r);
    
    \I2.MIC_REG2L3R_ADT_NET_834020_RD1__2936\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.MIC_REG2_312_adt_net_855644__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2L3R_ADT_NET_834020_RD1__453\);
    
    \I2.UN1_STATE1_31_I_1591\ : NOR2FT
      port map(A => \I2.STATE1l6r_net_1\, B => 
        \I2.STATE1l7r_net_1\, Y => \I2.N_3866_adt_net_61361_\);
    
    \I2.FCNT_n2\ : OR2
      port map(A => \I2.un1_STATE1_22\, B => \I2.FCNT_n2_tz_i\, Y
         => \I2.FCNT_n2_i\);
    
    \I2.resyn_0_I2_un1_trgcnt14_i\ : NAND2FT
      port map(A => \I2.N_3760_adt_net_15910_\, B => 
        \I2.un9_tdctrgi_i_0\, Y => \I2.N_3760\);
    
    \I1.N_304_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_304_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_304_Rd1__net_1\);
    
    \I3.un1_REGMAP_34_0_a2_0_a2_745\ : NOR2FT
      port map(A => \I3.un1_REGMAP_30\, B => 
        \I3.N_178_ADT_NET_1360__126\, Y => \I3.UN1_REGMAP_34_123\);
    
    REGl402r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_303_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl402r\);
    
    \I2.PIPE1_DT_30l7r\ : MUX2L
      port map(A => \I2.TDCDBSl7r_net_1\, B => 
        \I2.TDCDBSl5r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, Y
         => \I2.PIPE1_DT_30l7r_net_1\);
    
    \I3.PIPEA1_322\ : MUX2L
      port map(A => \I3.PIPEA1l24r_net_1\, B => 
        \I3.PIPEA1_12l24r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__251\, Y => 
        \I3.PIPEA1_322_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I57_Y_0_O2_1546\ : OR2
      port map(A => \I2.RAMDT4L1R_769\, B => 
        \I2.PIPE4_DT_I_IL1R_848\, Y => \I2.N357_adt_net_54497_\);
    
    \I2.un1_PIPE1_DT_0_sqmuxa_i_0_o2_0\ : OR2
      port map(A => \I2.N_3272_343\, B => \I2.END_CHAINB1_594\, Y
         => \I2.N_3885\);
    
    \I2.CHA_DATA8_2_I_1694\ : AND2FT
      port map(A => \I2.PIPE7_DTl28r_net_1\, B => \I2.N_4403\, Y
         => \I2.N_4398_adt_net_90118_\);
    
    \I2.BNCID_VECTrff_10_255_0\ : AO21
      port map(A => \I2.BNCID_VECTwa14_1_net_1\, B => 
        \I2.BNCID_VECTrff_8_257_0_a2_0\, C => 
        \I2.BNCID_VECTro_10\, Y => 
        \I2.BNCID_VECTrff_10_255_0_net_1\);
    
    F_SO_pad : IB33
      port map(PAD => F_SO, Y => F_SO_c);
    
    \I2.END_CHAINA1_708_1538\ : AND2
      port map(A => \I2.STATE1l12r_adt_net_855184__net_1\, B => 
        \I2.END_CHAINA1_1_sqmuxa_3\, Y => 
        \I2.END_CHAINA1_708_adt_net_53509_\);
    
    \I2.DTO_16_1_IVL23R_1103\ : AO21
      port map(A => \I2.DTO_1l23r\, B => \I2.N_196_53\, C => 
        \I2.DTO_16_1l23r_adt_net_30100_\, Y => 
        \I2.DTO_16_1l23r_adt_net_30116_\);
    
    \I5.COMMAND_4l2r\ : MUX2L
      port map(A => \I5.AIR_WDATAl2r_net_1\, B => REGl103r, S => 
        REGl7r, Y => \I5.COMMAND_4l2r_net_1\);
    
    \I2.LSRAM_IN_411\ : MUX2L
      port map(A => \I2.PIPE5_DTl27r_net_1\, B => 
        \I2.LSRAM_INl27r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_411_net_1\);
    
    \I3.PIPEB_89_2334\ : NOR2FT
      port map(A => \I3.PIPEBl10r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_89_adt_net_160293_\);
    
    \I2.WOFFSET_833\ : MUX2L
      port map(A => \I2.WOFFSETl6r_Rd1__net_1\, B => 
        \I2.N_4249_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835308_Rd1__net_1\, Y
         => \I2.WOFFSETl6r\);
    
    \I2.N_22_i_0_adt_net_855592_\ : BFR
      port map(A => \I2.N_22_i_0_adt_net_855596__net_1\, Y => 
        \I2.N_22_i_0_adt_net_855592__net_1\);
    
    \I3.VDBi_20_ivl3r\ : AND2
      port map(A => REGl51r, B => 
        \I3.REGMAPl9r_adt_net_854332__net_1\, Y => 
        \I3.VDBi_20l3r_adt_net_144750_\);
    
    \I2.PIPE5_DTl21r_1519_1788\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_697_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL21R_894\);
    
    \I1.REG_74_0_IVL278R_1941\ : NOR2FT
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l278r_adt_net_122893_\);
    
    \I3.PIPEA_255\ : MUX2L
      port map(A => \I3.PIPEAl24r_net_1\, B => 
        \I3.PIPEA_8l24r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854656__net_1\, Y
         => \I3.PIPEA_255_net_1\);
    
    \I2.FIDl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_422_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl6r);
    
    \I1.REG_15_sqmuxa_adt_net_1457__adt_net_854380_\ : BFR
      port map(A => \I1.REG_15_sqmuxa_adt_net_1457__net_1\, Y => 
        \I1.REG_15_sqmuxa_adt_net_1457__adt_net_854380__net_1\);
    
    \I5.AIR_WDATA_9l9r\ : AND2
      port map(A => \I5.SENS_ADDRl0r_net_1\, B => 
        \I5.sstate2l3r_net_1\, Y => \I5.AIR_WDATA_9l9r_net_1\);
    
    \I2.un1_PIPE1_DT_0_sqmuxa_i_0_o2\ : NOR2FT
      port map(A => \I2.STATE1L5R_591\, B => \I2.N_3885\, Y => 
        \I2.N_3891\);
    
    \I2.DTO_16_1_IV_0_0_1L0R_1213\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.DTO_9_ivl0r\, C => 
        \I2.DTO_16_1_iv_0_0_1l0r_adt_net_35382_\, Y => 
        \I2.DTO_16_1_iv_0_0_1l0r_adt_net_35388_\);
    
    \I3.UN1_STATE1_11_I_2345\ : NOR3FTT
      port map(A => \I3.REGMAPl10r_net_1\, B => \I3.N_276\, C => 
        \I3.WRITES_8\, Y => \I3.N_1902_adt_net_160759_\);
    
    \I1.REG_1_189\ : MUX2H
      port map(A => \REGl288r\, B => \I1.REG_74l288r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\, Y => 
        \I1.REG_1_189_net_1\);
    
    \I2.TOKOUT_FL\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKOUT_FL_674_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.TOKOUT_FL_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl20r\ : OR3
      port map(A => \I2.PIPE1_DT_42l20r_adt_net_47055_\, B => 
        \I2.PIPE1_DT_42l20r_adt_net_47067_\, C => 
        \I2.PIPE1_DT_42l20r_adt_net_47068_\, Y => 
        \I2.PIPE1_DT_42l20r\);
    
    TDCDB_padl21r : IB33
      port map(PAD => TDCDB(21), Y => TDCDB_cl21r);
    
    REGl177r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_78_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl177r\);
    
    TDCDB_padl5r : IB33
      port map(PAD => TDCDB(5), Y => TDCDB_cl5r);
    
    N_1_I3_TCNT3_c3 : AND2
      port map(A => \I3.TCNT3l3r_net_1\, B => \I3.TCNT3_c2\, Y
         => \I3.TCNT3_c3\);
    
    \I3.un136_reg_ads_0_a2_2_a2_0_986\ : NAND2FT
      port map(A => \I3.VASl2r_net_1\, B => \I3.N_548_367\, Y => 
        \I3.N_549_364\);
    
    \I2.DTE_cl_0_sqmuxa_2_0_a2_0_a2_0\ : OR2FT
      port map(A => \I2.N_4241_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, Y => 
        \I2.DTE_cl_0_sqmuxa_2_0\);
    
    \I5.TEMPDATAl6r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_80_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl6r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I207_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl11r\, B => 
        \I2.PIPE7_DTl11r_net_1\, Y => 
        \I2.SUB_21x21_fast_I207_Y_0\);
    
    \I1.SSTATEL10R_3096\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_43_i_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL10R_882\);
    
    \I2.PIPE1_DT_12l7r\ : MUX2L
      port map(A => \I2.TDCDASl7r_net_1\, B => 
        \I2.TDCDASl5r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, Y
         => \I2.PIPE1_DT_12l7r_net_1\);
    
    \I2.un1_STATE1_30\ : OR3FTT
      port map(A => \I2.N_3870\, B => 
        \I2.STATE1_nsl6r_adt_net_23511_\, C => 
        \I2.END_CHAINA1_708_adt_net_53509_\, Y => 
        \I2.un1_STATE1_30_net_1\);
    
    \I2.PIPE1_DT_741\ : MUX2L
      port map(A => \I2.PIPE1_DTl14r_net_1\, B => 
        \I2.PIPE1_DT_42l14r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854576__net_1\, 
        Y => \I2.PIPE1_DT_741_net_1\);
    
    \I2.STATE1_ns_i_o2l9r_966\ : OR3
      port map(A => FLUSH, B => \I2.FCNT_c1\, C => 
        \I2.FCNTL2R_599\, Y => \I2.N_3272_344\);
    
    \I2.L2TYPE_4_IL1R_1640\ : AND2
      port map(A => \I2.L2TYPE_i_0_il1r\, B => 
        \I2.N_4451_adt_net_68574_\, Y => 
        \I2.N_4451_adt_net_68617_\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__2842\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854736__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__200\);
    
    \I2.DT_TEMPl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_784_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl23r_net_1\);
    
    REGl227r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_128_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl227r\);
    
    \I3.PULSE_336\ : MUX2L
      port map(A => PULSEl6r, B => \I3.PULSE_46l6r\, S => 
        \I3.N_1409_adt_net_854740__net_1\, Y => 
        \I3.PULSE_336_net_1\);
    
    \I2.un1_tdc_res_43_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl409r, Y => 
        \I2.N_4624_i_0\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I122_Y_0\ : AOI21
      port map(A => \I2.N_64_0_adt_net_855028__net_1\, B => 
        \I2.N_93_0\, C => \I2.N_84_0\, Y => \I2.N537_i_0\);
    
    \I2.MIC_REG2l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_310_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2l1r_net_1\);
    
    \I2.CHAIN_ERR_DIS_448_1713\ : AOI21TTF
      port map(A => BNC_RES_E, B => \I2.CHAIN_RDY_net_1\, C => 
        REGl26r, Y => \I2.CHAIN_ERR_DIS_448_adt_net_92599_\);
    
    \I2.SUB9_576\ : MUX2H
      port map(A => \I2.SUB9l8r_net_1\, B => \I2.SUB9_1l8r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_576_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I154_Y_0\ : OAI21
      port map(A => \I2.PIPE4_DTl15r_net_1\, B => 
        \I2.PIPE4_DTl16r_net_1\, C => \I2.RAMDT4L12R_795\, Y => 
        \I2.N502_i_0_adt_net_490246_\);
    
    \I2.WOFFSETl12r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl12r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl12r_Rd1__net_1\);
    
    \I2.REG_1_n2\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => \I2.REG_1_n2_0_net_1\, Y => \I2.REG_1_n2_net_1\);
    
    \I2.SUB9_578\ : MUX2H
      port map(A => \I2.SUB9l10r_net_1\, B => \I2.SUB9_1l10r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_578_net_1\);
    
    \I2.L2TYPE_602\ : MUX2L
      port map(A => \I2.L2TYPE_i_0_il13r\, B => \I2.N_4439\, S
         => \I2.N_4482_0\, Y => \I2.L2TYPE_602_net_1\);
    
    DPR_padl25r : IB33
      port map(PAD => DPR(25), Y => DPR_cl25r);
    
    REGl250r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_151_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl250r\);
    
    \I2.PIPE8_DT_21_i_0l30r\ : AOI21
      port map(A => \I2.PIPE7_DTl31r_net_1\, B => 
        \I2.PIPE8_DTl30r_net_1\, C => 
        \I2.PIPE7_DTl30r_adt_net_855172__net_1\, Y => 
        \I2.PIPE8_DT_21_i_0_il30r\);
    
    \I3.VDBi_57_0_ivl31r\ : OAI21FTF
      port map(A => \I3.VDBi_31l31r_net_1\, B => \I3.N_1905\, C
         => \I3.VDBi_57l31r_adt_net_137844_\, Y => 
        \I3.VDBi_57l31r\);
    
    \I2.DT_TEMP_7l9r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, B => 
        \I2.N_4047\, Y => \I2.DT_TEMP_7l9r_net_1\);
    
    \I3.VADm_0_a3l8r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl8r_net_1\, Y => \I3.VADml8r\);
    
    \I1.REG_74_0_IVL397R_1792\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_30_sqmuxa_adt_net_854372__net_1\, Y => 
        \I1.REG_74l397r_adt_net_110358_\);
    
    \I2.SRAM_FULL\ : DFFC
      port map(CLK => CLK_c, D => \I2.SRAM_FULL_488_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.SRAM_FULL_net_1\);
    
    \I3.un1_STATE2_15_1_adt_net_1342_\ : OR2
      port map(A => \I3.STATE2_nsl0r_adt_net_136048_\, B => 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\, Y => 
        \I3.un1_STATE2_15_1_adt_net_1342__net_1\);
    
    \I3.un1_NOEDTKi_0_sqmuxa_adt_net_4101_\ : AO21
      port map(A => \I3.DSS_net_1\, B => \I3.STATE1_ipl7r\, C => 
        \I3.un1_NOEDTKi_0_sqmuxa_adt_net_135826__net_1\, Y => 
        \I3.un1_NOEDTKi_0_sqmuxa_adt_net_4101__net_1\);
    
    \I2.ROFFSET_n1\ : XOR2
      port map(A => \I2.N_1355\, B => \I2.N_1357\, Y => 
        \I2.ROFFSET_n1_net_1\);
    
    \I3.VDBoffa_48\ : OR3
      port map(A => \I3.VDBoffa_48_adt_net_163928_\, B => 
        \I3.VDBoffa_31l4r_adt_net_163889_\, C => 
        \I3.VDBoffa_31l4r_adt_net_163890_\, Y => 
        \I3.VDBoffa_48_net_1\);
    
    ADE_padl0r : OB33PH
      port map(PAD => ADE(0), A => ADE_cl0r);
    
    \I3.un141_reg_ads_0_a2_0_a2\ : OR3FFT
      port map(A => \I3.VASl2r_net_1\, B => \I3.N_548\, C => 
        \I3.N_586_adt_net_165970_\, Y => \I3.N_639\);
    
    \I2.REG_0L3R_ADT_NET_19771_RD1__3101\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.REG_0l3r_adt_net_19771_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.REG_0L3R_ADT_NET_19771_RD1__887\);
    
    REGl332r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_233_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl332r\);
    
    INT_ERRA_pad : IB33
      port map(PAD => INT_ERRA, Y => INT_ERRA_c);
    
    \I2.DT_SRAM_0l16r\ : MUX2L
      port map(A => \I2.PIPE10_DTl16r_net_1\, B => 
        \I2.PIPE5_DTl16r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854224__net_1\, Y => 
        \I2.N_884\);
    
    \I2.PIPE1_DT_42_1_IVL6R_1489\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855756__net_1\, B => 
        \I2.PIPE1_DT_30l6r_net_1\, C => 
        \I2.PIPE1_DT_42l6r_adt_net_50924_\, Y => 
        \I2.PIPE1_DT_42l6r_adt_net_50940_\);
    
    \I2.DTE_21_1_IV_0L8R_1312\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, 
        B => \I2.DT_TEMPl8r_net_1\, C => 
        \I2.DTE_21_1l8r_adt_net_38737_\, Y => 
        \I2.DTE_21_1l8r_adt_net_38752_\);
    
    \I2.STATE3l9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_i_il10r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE3l9r_net_1\);
    
    \I2.PIPE4_DTl5r_adt_net_854412__adt_net_855600_\ : BFR
      port map(A => \I2.PIPE4_DTl5r_adt_net_854412__net_1\, Y => 
        \I2.PIPE4_DTl5r_adt_net_854412__adt_net_855600__net_1\);
    
    \I2.MIC_ERR_REGS_372\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl44r_net_1\, B => 
        \I2.MIC_ERR_REGSl43r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_372_net_1\);
    
    \I1.REG_74_0_IVL404R_1785\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_30_sqmuxa_adt_net_854372__net_1\, Y => 
        \I1.REG_74l404r_adt_net_109656_\);
    
    \I5.BITCNTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.BITCNT_84_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.BITCNTl2r_net_1\);
    
    \I2.PIPE4_DTl12r_1249_1748\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL12R_855\);
    
    \I2.PIPE1_DT_42_0_IVL31R_1351\ : NOR2FT
      port map(A => \I2.TDCDASl31r_net_1\, B => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        Y => \I2.PIPE1_DT_42l31r_adt_net_45035_\);
    
    \I3.un2_clear_stat_i_a3\ : NAND2
      port map(A => EVRDY_c, B => CLEAR_STAT_12, Y => 
        \I3.N_2137_i_0\);
    
    \I1.REG_74_0_IVL328R_1888\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l328r_adt_net_118260_\);
    
    \I4.bcnt_i_0_il2r\ : DFFC
      port map(CLK => CLK_c, D => \I4.bcnt_7_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I4.bcnt_i_0_il2r_net_1\);
    
    \I1.PAGECNTL5R_2877\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_322_adt_net_854384__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL5R_309\);
    
    \I2.TDCTRGi_266\ : MUX2L
      port map(A => TDCTRG_c, B => \I2.STATE4_il0r\, S => 
        \I2.STATE4l2r_net_1\, Y => \I2.TDCTRGi_266_net_1\);
    
    \I2.TDCDASl25r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl25r, Q => 
        \I2.TDCDASl25r_net_1\);
    
    \I2.TOKENB_CNT_i_0l1r\ : NAND2
      port map(A => CLEAR_STAT_12, B => \I2.TOKENTOB_RES_net_1\, 
        Y => \I2.un12_clear_stat_i\);
    
    \I3.REG_1_174\ : MUX2L
      port map(A => VDB_inl25r, B => REGl73r, S => 
        \I3.N_1935_adt_net_855320__net_1\, Y => \I3.REG_1_174_0\);
    
    \I2.STATEel2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATEe_nsl2r\, CLR => 
        \I2.STATEe_i_0l0r_net_1\, Q => \I2.STATEe_ipl2r\);
    
    \I2.MIC_ERR_REGS_353\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl25r_net_1\, B => 
        \I2.MIC_ERR_REGSl24r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_353_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL22R_1382\ : NOR2FT
      port map(A => REGl426r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, Y => 
        \I2.PIPE1_DT_42l22r_adt_net_46757_\);
    
    \I1.REG_27_sqmuxa_adt_net_854808_\ : BFR
      port map(A => \I1.REG_27_sqmuxa\, Y => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\);
    
    \I2.N_4646_1_adt_net_19637_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_19637_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_adt_net_19637_Rd1__net_1\);
    
    \I3.VDBI_57_0_IVL11R_2210\ : AO21
      port map(A => \I3.PIPEAl11r_net_1\, B => \I3.N_90_i_0_1\, C
         => \I3.VDBi_57l11r_adt_net_141431_\, Y => 
        \I3.VDBi_57l11r_adt_net_141440_\);
    
    \I3.VDBOFFB_30_IV_0L3R_2421\ : AND2
      port map(A => \REGl352r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162508_\);
    
    \I2.un1_END_EVNT1_0_sqmuxa_i_0_m3\ : MUX2L
      port map(A => \I2.N_3882\, B => \I2.STATE1L9R_631\, S => 
        \I2.STATE1L18R_628\, Y => \I2.N_3888\);
    
    \I2.DTO_9_iv_0_o2l2r\ : OAI21TTF
      port map(A => \I2.N_4283_i_0_adt_net_854972__net_1\, B => 
        \I2.DT_TEMPl2r_net_1\, C => 
        \I2.DTO_9_ivl2r_adt_net_34812_\, Y => \I2.DTO_9_ivl2r\);
    
    \I2.DTE_21_1_IV_2L3R_1335\ : AND2
      port map(A => GA_cl3r, B => 
        \I2.STATE2l1r_adt_net_855120__net_1\, Y => 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39303_\);
    
    \I2.DTESl20r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl20r, Q => 
        \I2.DTESl20r_net_1\);
    
    \I2.CRC32_802\ : MUX2L
      port map(A => \I2.CRC32l7r_net_1\, B => \I2.N_3924\, S => 
        \I2.N_2826_1_ADT_NET_794__332\, Y => \I2.CRC32_802_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2399\ : OR2
      port map(A => \I3.VDBoffb_30l5r_adt_net_162171_\, B => 
        \I3.VDBoffb_30l5r_adt_net_162172_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162177_\);
    
    NRDMEB_pad : OB33PH
      port map(PAD => NRDMEB, A => NRDMEB_c);
    
    \I2.RAMAD1_669\ : MUX2L
      port map(A => \I2.RAMAD1_12l15r_net_1\, B => 
        \I2.RAMAD1l15r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__170\, Y => 
        \I2.RAMAD1_669_net_1\);
    
    \I2.STATE1l12r_adt_net_855180_\ : BFR
      port map(A => \I2.STATE1L12R_646\, Y => 
        \I2.STATE1l12r_adt_net_855180__net_1\);
    
    \I2.OFFSET_37_15l1r\ : MUX2L
      port map(A => \REGl230r\, B => \REGl166r\, S => 
        \I2.PIPE7_DTL27R_73\, Y => \I2.N_748\);
    
    \I2.REG_1_C12_I_1737\ : AND2
      port map(A => REGl44r, B => \I2.N_3856\, Y => 
        \I2.N_3841_i_0_adt_net_101174_\);
    
    \I2.BNCID_VECT_tile_DOUTl3r\ : MUX2L
      port map(A => \I2.DIN_REG1_0l3r\, B => \I2.DOUT_TMP_0l3r\, 
        S => \I2.N_13\, Y => \I2.BNCID_VECTrxl3r\);
    
    \I1.REG_74_4_I_A2_404_N_4_I_ADT_NET_1465__2838\ : AND2
      port map(A => \I1.N_268_Rd1__net_1\, B => \I1.N_254_195\, Y
         => \I1.REG_74_4_I_A2_404_N_4_I_ADT_NET_1465__193\);
    
    \I2.REG_1_c13_i_o2\ : NAND3
      port map(A => REGl45r, B => REGl44r, C => \I2.N_3856\, Y
         => \I2.N_3859\);
    
    \I2.PHASE_i_0\ : INV
      port map(A => NOESRAME_C_243, Y => \I2.NOESRAME_c_i_0\);
    
    \I2.DT_TEMP_7l15r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854244__net_1\, B => 
        \I2.DT_SRAMl15r_net_1\, Y => \I2.DT_TEMP_7l15r_net_1\);
    
    \I2.PIPE10_DT_633\ : MUX2L
      port map(A => \I2.PIPE10_DTl28r_net_1\, B => 
        \I2.PIPE9_DTl28r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_633_net_1\);
    
    \I3.un206_reg_ads_0_a2_1_a2\ : OR2FT
      port map(A => \I3.VASl5r_net_1\, B => \I3.VASl3r_net_1\, Y
         => \I3.N_554\);
    
    \I1.N_1193_adt_net_1562_\ : OAI21FTF
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.N_368\, C => 
        \I1.N_1193_adt_net_133987__net_1\, Y => 
        \I1.N_1193_adt_net_1562__net_1\);
    
    \I2.PIPE1_DTl20r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_747_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl20r_net_1\);
    
    \I3.PIPEA_8_0l20r\ : MUX2L
      port map(A => DPR_cl20r, B => \I3.PIPEA1l20r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855360__net_1\, Y => \I3.N_229\);
    
    \I5.SBYTE_72\ : MUX2H
      port map(A => \I5.SBYTEl7r_net_1\, B => \I5.SBYTE_9l7r\, S
         => \I5.N_406\, Y => \I5.SBYTE_72_net_1\);
    
    \I2.DTE_21_1l21r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l21r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l21r_Rd1__net_1\);
    
    \I3.N_1935_adt_net_855320_\ : BFR
      port map(A => \I3.N_1935\, Y => 
        \I3.N_1935_adt_net_855320__net_1\);
    
    \I1.REG_74_0_IVL268R_1955\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, Y => 
        \I1.REG_74l268r_adt_net_124027_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I121_Y_i_a2\ : NAND2FT
      port map(A => \I2.N_2360_tz_tz\, B => \I2.N_17\, Y => 
        \I2.N_158_0\);
    
    \I2.PIPE3_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl14r_net_1\);
    
    \I3.N_1414_i_i_o3_i_o2_0\ : OR2
      port map(A => \I3.STATE1_IPL2R_885\, B => \I3.N_1764\, Y
         => \I3.N_1910_0\);
    
    TDCDB_padl13r : IB33
      port map(PAD => TDCDB(13), Y => TDCDB_cl13r);
    
    \I2.OFFSET_37_20l1r\ : MUX2L
      port map(A => \I2.N_780\, B => \I2.N_772\, S => 
        \I2.PIPE7_DTL26R_359\, Y => \I2.N_788\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I202_Y\ : XOR2FT
      port map(A => \I2.N513\, B => \I2.SUB_21x21_fast_I202_Y_0\, 
        Y => \I2.SUB8_2l6r\);
    
    \I2.END_EVNT5_1143\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT5_405\);
    
    \I2.PIPE5_DTl21r_1519_1787\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_697_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL21R_893\);
    
    REGl372r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_273_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl372r\);
    
    \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776_\ : BFR
      port map(A => \I2.MIC_REG1_0_sqmuxa_0_net_1\, Y => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\);
    
    \I2.PIPE7_DTL27R_2793\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_86\);
    
    \I2.ADE_4l8r\ : MUX2H
      port map(A => \I2.WOFFSETl9r\, B => \I2.ROFFSETl9r_net_1\, 
        S => NOESRAME_c, Y => \I2.ADE_4l8r_net_1\);
    
    \I2.UN1_NWPIPE7_2_1670\ : OAI21TTF
      port map(A => \I2.CHA_DATA8_net_1\, B => 
        \I2.CHB_DATA8_net_1\, C => 
        \I2.un1_NWPIPE7_2_adt_net_73600_\, Y => 
        \I2.un1_NWPIPE7_2_adt_net_73606_\);
    
    \I2.FIDl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_418_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl2r);
    
    \I1.REG_1_235\ : MUX2H
      port map(A => \REGl334r\, B => \I1.REG_74l334r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y => 
        \I1.REG_1_235_net_1\);
    
    \I2.ROFFSET_910\ : MUX2H
      port map(A => \I2.ROFFSETl8r_net_1\, B => 
        \I2.ROFFSET_n8_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_910_net_1\);
    
    \I2.DTO_16_1_IVL15R_1140\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855680__net_1\, B => 
        \I2.DTO_9l15r\, Y => \I2.DTO_16_1l15r_adt_net_31948_\);
    
    \I2.WPAGE_c1\ : AND2
      port map(A => \I2.WPAGEl13r_net_1\, B => 
        \I2.WPAGEl12r_net_1\, Y => \I2.WPAGE_c1_net_1\);
    
    \I2.PIPE8_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_551_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl23r_net_1\);
    
    REGl386r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_287_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl386r\);
    
    \I2.END_CHAINB1_709_adt_net_2397_\ : OR2
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855240__net_1\, 
        B => \I2.TOKOUTBS_629\, Y => 
        \I2.END_CHAINB1_709_adt_net_2397__net_1\);
    
    \I2.PIPE1_DT_2_sqmuxa_1_1\ : NOR2FT
      port map(A => \I2.TDCGDB1_580\, B => \I2.N_3889_178\, Y => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_net_1\);
    
    \I1.REG_74_0_ivl338r\ : AO21
      port map(A => \REGl338r\, B => \I1.N_209\, C => 
        \I1.REG_74l338r_adt_net_117400_\, Y => \I1.REG_74l338r\);
    
    \I2.MIC_ERR_REGS_345\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl17r_net_1\, B => 
        \I2.MIC_ERR_REGSl16r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\, Y => 
        \I2.MIC_ERR_REGS_345_net_1\);
    
    \I1.REG_74_0_IVL166R_2068\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l166r_adt_net_133579_\);
    
    \I3.VDBI_57_0_IV_0L19R_2174\ : AO21
      port map(A => \I3.VDBil19r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l19r_adt_net_139383_\, Y => 
        \I3.VDBi_57l19r_adt_net_139393_\);
    
    \I2.PIPE4_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl20r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl20r_net_1\);
    
    \I2.TDCGDB1\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => TDCGDB_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.TDCGDB1_net_1\);
    
    \I2.PIPE8_DT_21_i_o2l30r\ : OR2
      port map(A => \I2.PIPE7_DTl31r_net_1\, B => 
        \I2.PIPE7_DTl30r_adt_net_855172__net_1\, Y => \I2.N_4401\);
    
    \I3.REGMAPl0r_1159\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un2_reg_ads_0_a2_0_a3_net_1\, Q => \I3.REGMAPL0R_421\);
    
    \I2.PIPE5_DT_6l7r\ : MUX2L
      port map(A => 
        \I2.PIPE4_DTl7r_adt_net_854552__adt_net_854948__net_1\, B
         => \I2.N_1076\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\, Y => 
        \I2.PIPE5_DT_6l7r_net_1\);
    
    \I2.PIPE5_DTl31r_1513\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_707_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL31R_620\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I42_Y_1647\ : AO21
      port map(A => \I2.N_3539_i_i\, B => \I2.G_1_2\, C => 
        \I2.N_3541_i_i\, Y => \I2.N307_1_adt_net_69278_\);
    
    \I2.N_4186_i_0_o2\ : NAND2
      port map(A => NOESRAME_C_239, B => 
        \I2.WOFFSETl0r_adt_net_854644__net_1\, Y => \I2.N_237\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I11_P0N_i_a4\ : OR2
      port map(A => \I2.RAMDT4L5R_821\, B => 
        \I2.PIPE4_DTl11r_net_1\, Y => \I2.N_91\);
    
    \I2.RAMDT4l5r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l5r_net_1\);
    
    \I1.N_311_i_i_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_311_i_i_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.N_311_i_i_Rd1__net_1\);
    
    \I2.REG_0l3r_adt_net_19773_Ra1_\ : OA21
      port map(A => \I3.REG1_136_net_1\, B => \I3.REG2_144_net_1\, 
        C => \I3.REG3_128_net_1\, Y => 
        \I2.REG_0l3r_adt_net_19773_Ra1__net_1\);
    
    \I1.REG_2_sqmuxa_0_a2_0\ : OR2FT
      port map(A => \I1.PAGECNTL5R_311\, B => 
        \I1.N_237_adt_net_854804__net_1\, Y => \I1.N_259\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I189_Y\ : XOR2
      port map(A => \I2.N498_0\, B => 
        \I2.ADD_21x21_fast_I189_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l19r\);
    
    \I3.TCNT4_388\ : XOR2
      port map(A => \I3.TCNT4_i_0_il0r_net_1\, B => 
        \I3.TICKl2r_net_1\, Y => \I3.TCNT4_388_net_1\);
    
    \I2.FID_7_0_IVL8R_1717\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl56r, C => 
        \I2.FID_7l8r_adt_net_92739_\, Y => 
        \I2.FID_7l8r_adt_net_92747_\);
    
    \I1.N_50_0_ADT_NET_1409__2870\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__541\, B => 
        \I1.N_50_0_ADT_NET_109751__258\, Y => 
        \I1.N_50_0_ADT_NET_1409__292\);
    
    \I3.VDBI_57_IV_0_0L7R_2230\ : AO21
      port map(A => \I3.PIPEAl7r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l7r_adt_net_143093_\, Y => 
        \I3.VDBi_57l7r_adt_net_143110_\);
    
    \I2.PIPE4_DTl12r_1249_1749\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL12R_856\);
    
    \I2.STOP_RDSRAM\ : DFFC
      port map(CLK => CLK_c, D => \I2.STOP_RDSRAM_453_i_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STOP_RDSRAM_net_1\);
    
    \I2.DT_SRAMl4r\ : MUX2L
      port map(A => \I2.N_872\, B => \I2.PIPE2_DTl4r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.DT_SRAMl4r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I139_Y_i_a4\ : OA21
      port map(A => \I2.PIPE4_DTl10r_net_1\, B => 
        \I2.PIPE4_DTL11R_410\, C => \I2.RAMDT4L12R_146\, Y => 
        \I2.N_96_0_adt_net_58152_\);
    
    \I2.un7_bnc_id_1_I_38\ : XOR2
      port map(A => \I2.BNC_IDl7r_net_1\, B => \I2.N_24_1\, Y => 
        \I2.I_38_0\);
    
    \I2.DT_TEMP_7l2r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, B => 
        \I2.N_4193\, Y => \I2.DT_TEMP_7l2r_net_1\);
    
    \I2.DTE_21_1_IV_0L26R_1240\ : AND2
      port map(A => \I2.DT_TEMPl26r_net_1\, B => \I2.N_4038_233\, 
        Y => \I2.DTE_21_1l26r_adt_net_36951_\);
    
    VAD_padl22r : OTB33PH
      port map(PAD => VAD(22), A => \I3.VADml22r\, EN => 
        NOEAD_c_i_0);
    
    \I2.PIPE1_DT_42_1_ivl15r\ : OR3
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48707_\, B => 
        \I2.PIPE1_DT_42l15r_adt_net_48716_\, C => 
        \I2.PIPE1_DT_42l15r_adt_net_48717_\, Y => 
        \I2.PIPE1_DT_42l15r\);
    
    \I2.CRC32_800\ : MUX2L
      port map(A => \I2.CRC32l5r_net_1\, B => \I2.N_3922\, S => 
        \I2.N_2826_1_adt_net_794__net_1\, Y => 
        \I2.CRC32_800_net_1\);
    
    \I3.VDBOFFA_44_2636\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal0r_net_1\, Y => 
        \I3.VDBoffa_44_adt_net_164688_\);
    
    \I2.MIC_REG2_316\ : MUX2H
      port map(A => \I2.MIC_REG2l7r_net_1\, B => 
        \I2.MTDIAS_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768__net_1\, Y => 
        \I2.MIC_REG2_316_net_1\);
    
    \I3.VDBi_57_0_ivl16r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855380__net_1\, B => 
        \I3.VDBi_31l16r_net_1\, C => 
        \I3.VDBi_57l16r_adt_net_139767_\, Y => \I3.VDBi_57l16r\);
    
    \I2.PIPE3_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl17r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl17r_net_1\);
    
    \I1.REG_74l276r\ : OR3FFT
      port map(A => \I1.REG_74_1l268r\, B => \I1.N_145_12\, C => 
        \I1.REG_13_sqmuxa\, Y => \I1.N_145\);
    
    \I1.REG_1_222\ : MUX2H
      port map(A => \REGl321r\, B => \I1.REG_74l321r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y => 
        \I1.REG_1_222_net_1\);
    
    \I3.VDBi_57_0_iv_0_a2_0l8r\ : AND2
      port map(A => \I3.STATE1_IPL2R_886\, B => \I3.N_57_i_0_0\, 
        Y => \I3.N_2034\);
    
    \I2.G_EVNT_NUM_n10_0_a2_1\ : AND2FT
      port map(A => EV_RES_C_568, B => \I2.G_EVNT_NUMl10r_net_1\, 
        Y => \I2.N_285_1\);
    
    \I2.SUB8_1_sqmuxa_0_adt_net_855160_\ : BFR
      port map(A => \I2.SUB8_1_sqmuxa_0\, Y => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855160__net_1\);
    
    \I2.PIPE1_DT_30l17r\ : MUX2L
      port map(A => \I2.TDCDBSl17r_net_1\, B => 
        \I2.TDCDBSl15r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, Y
         => \I2.PIPE1_DT_30l17r_net_1\);
    
    \I2.DTE_21_1_iv_0_o2_1_0l21r_855\ : OAI21FTT
      port map(A => \I2.STATE2L3R_439\, B => \I2.N_4283_I_0_234\, 
        C => \I2.DTO_cl_0_sqmuxa_0\, Y => \I2.N_4038_233\);
    
    \I2.TDCGDBi_673\ : MUX2H
      port map(A => TDCGDB_c, B => \I2.un1_STATE1_24\, S => 
        \I2.N_3866\, Y => \I2.TDCGDBi_673_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I151_Y_I_A2_2_1551\ : AO21
      port map(A => \I2.RAMDT4L5R_820\, B => 
        \I2.PIPE4_DTl19r_net_1\, C => 
        \I2.N_152_i_adt_net_4109__net_1\, Y => 
        \I2.N_152_i_adt_net_54890_\);
    
    REGl241r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_142_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl241r\);
    
    \I2.DTE_1l30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_868_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l30r_net_1\);
    
    \I3.REG_1l145r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_193_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl145r\);
    
    \I2.MIC_ERR_REGSl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_360_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl31r_net_1\);
    
    \I1.N_113_ADT_NET_3714__2866\ : OR2
      port map(A => \I1.N_41_9\, B => 
        \I1.N_113_adt_net_126306__net_1\, Y => 
        \I1.N_113_ADT_NET_3714__271\);
    
    \I1.REG_74_0_ivl344r\ : AO21
      port map(A => \REGl344r\, B => \I1.N_217\, C => 
        \I1.REG_74l344r_adt_net_116670_\, Y => \I1.REG_74l344r\);
    
    \I3.STATE2_ns_o3_1l3r\ : AND2FT
      port map(A => \I3.STATE2L2R_721\, B => 
        \I3.N_1463_i_adt_net_1279__net_1\, Y => \I3.N_1463_i_1\);
    
    \I2.PIPE1_DT_742\ : MUX2L
      port map(A => \I2.PIPE1_DTl15r_net_1\, B => 
        \I2.PIPE1_DT_42l15r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854576__net_1\, 
        Y => \I2.PIPE1_DT_742_net_1\);
    
    \I2.DTE_21_1_IV_0L12R_1291\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, 
        B => \I2.DT_TEMPl12r_net_1\, C => 
        \I2.DTE_21_1l12r_adt_net_38281_\, Y => 
        \I2.DTE_21_1l12r_adt_net_38296_\);
    
    \I2.TDCl0r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TDC_650_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TDCl0r_net_1\);
    
    \I2.FID_7_0_ivl19r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl19r_net_1\, 
        C => \I2.FID_7l19r_adt_net_17525_\, Y => \I2.FID_7l19r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I201_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl5r\, B => 
        \I2.PIPE7_DTl5r_net_1\, Y => \I2.SUB_21x21_fast_I201_Y_0\);
    
    \I1.REG_1_224\ : MUX2H
      port map(A => \REGl323r\, B => \I1.REG_74l323r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y => 
        \I1.REG_1_224_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I138_Y_0_o2_1\ : OA21
      port map(A => \I2.PIPE4_DTL11R_843\, B => 
        \I2.PIPE4_DTL12R_858\, C => \I2.RAMDT4L5R_138\, Y => 
        \I2.N_75\);
    
    FID_padl20r : OB33PH
      port map(PAD => FID(20), A => FID_cl20r);
    
    \I3.STATE1_423\ : OR2
      port map(A => \I3.STATE1_ipl1r\, B => \I3.N_1186\, Y => 
        \I3.N_1189\);
    
    \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272_\ : BFR
      port map(A => \I3.un1_STATE2_7_1_adt_net_1473__net_1\, Y
         => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\);
    
    \I2.STATE4l2r\ : DFFS
      port map(CLK => CLK_c, D => \I2.STATE4_ns_a3_il0r_net_1\, 
        SET => CLEAR_STAT_i_0, Q => \I2.STATE4l2r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I109_Y\ : OAI21
      port map(A => \I2.N321_0\, B => \I2.N324\, C => \I2.N320\, 
        Y => \I2.N363\);
    
    \I3.NDTKIN\ : OR2
      port map(A => \I3.CLOSEDTK_net_1\, B => NOEDTK_C_14, Y => 
        NDTKIN_c);
    
    \I2.EVNT_NUM_n9_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl9r_net_1\, B => 
        \I2.EVNT_NUM_c8_net_1\, Y => \I2.EVNT_NUM_n9_tz_i\);
    
    \I2.DTE_21_1_IV_0L13R_1284\ : AND2
      port map(A => \I2.N_4048\, B => 
        \I2.N_199_0_ADT_NET_1054__36\, Y => 
        \I2.DTE_21_1l13r_adt_net_38169_\);
    
    \I2.PIPE10_DT_17_il17r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l4r_net_1\, C => \I2.PIPE10_DT_17_i_0l17r_net_1\, 
        Y => \I2.N_3803\);
    
    \I2.DT_TEMPl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_761_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl0r_net_1\);
    
    \I2.DT_SRAMl12r\ : MUX2L
      port map(A => \I2.N_880\, B => \I2.PIPE2_DTl12r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672__net_1\, 
        Y => \I2.DT_SRAMl12r_net_1\);
    
    \I1.REG_74_0_iv_0l223r\ : AO21
      port map(A => \FBOUTl2r\, B => \I1.N_12233_i\, C => 
        \I1.REG_74l223r_adt_net_128394_\, Y => \I1.REG_74l223r\);
    
    \I2.DTO_9_IVL7R_1184\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl7r_net_1\, C => \I2.DTO_9l7r_adt_net_33660_\, 
        Y => \I2.DTO_9l7r_adt_net_33668_\);
    
    \I3.VDBOFFB_52_2492\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl0r_net_1\, Y => 
        \I3.VDBoffb_52_adt_net_163170_\);
    
    \I3.PIPEBl5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_84_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl5r_net_1\);
    
    \I2.PIPE1_DT_42_1_iv_1l24r\ : OAI21TTF
      port map(A => REGl428r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_1_il24r_adt_net_46469_\, Y => 
        \I2.PIPE1_DT_42_1_iv_1_il24r\);
    
    \I2.ROFFSET_n8\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\, B => 
        \I2.ROFFSET_n8_tz_i\, Y => \I2.ROFFSET_n8_net_1\);
    
    \I1.REG_74_0_ivl289r\ : AO21
      port map(A => \REGl289r\, B => \I1.N_161\, C => 
        \I1.REG_74l289r_adt_net_121947_\, Y => \I1.REG_74l289r\);
    
    \I2.RAMDT4L12R_3047\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_801\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I54_Y_1684\ : AND2FT
      port map(A => \I2.LSRAM_OUTl12r\, B => 
        \I2.PIPE7_DTl12r_net_1\, Y => \I2.N304_0_adt_net_87004_\);
    
    \I3.VDBI_57_0_IV_0L20R_2169\ : AO21
      port map(A => REGl68r, B => \I3.N_1839\, C => 
        \I3.VDBi_57l20r_adt_net_139285_\, Y => 
        \I3.VDBi_57l20r_adt_net_139290_\);
    
    \I3.STATE1_ns_0l0r\ : OR2
      port map(A => \I3.STATE1_nsl0r_adt_net_135920_\, B => 
        \I3.un1_NOEDTKi_0_sqmuxa_adt_net_4101__net_1\, Y => 
        \I3.STATE1_nsl0r\);
    
    \I3.VDBI_57_0_IV_0L18R_2175\ : AND2FT
      port map(A => \I3.N_1917_adt_net_855336__net_1\, B => 
        \I3.REGl151r\, Y => \I3.VDBi_57l18r_adt_net_139485_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I140_Y_0\ : AO21FTF
      port map(A => \I2.N_74_I_0_I_132\, B => 
        \I2.N519_adt_net_54631_\, C => \I2.N_70\, Y => \I2.N519\);
    
    \I3.VDBi_355\ : MUX2L
      port map(A => \I3.VDBil15r_net_1\, B => \I3.VDBi_57l15r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_355_net_1\);
    
    \I2.un1_tdc_res_44_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl411r, Y => 
        \I2.N_4625_i_0\);
    
    F_SI_pad : OB33PH
      port map(PAD => F_SI, A => F_SI_c);
    
    \I3.VDBml2r\ : MUX2L
      port map(A => \I3.VDBil2r_net_1\, B => \I3.N_144\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml2r_net_1\);
    
    \I2.TRGSERVl2r_1477\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l2r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVL2R_584\);
    
    \I2.LEAD_FLAG6_7_i_0l5r\ : AOI21
      port map(A => \I2.N_219\, B => \I2.N_483\, C => \I2.N_222\, 
        Y => \I2.N_4530_adt_net_64028_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I151_Y_i_a2_3\ : AOI21TTF
      port map(A => \I2.RAMDT4L12R_793\, B => 
        \I2.PIPE4_DTl16r_net_1\, C => \I2.N_163_0_adt_net_55087_\, 
        Y => \I2.N_163_0\);
    
    \I3.PULSE_46_0_IV_0_0L9R_2288\ : AND3
      port map(A => VDB_inl1r, B => \I3.REGMAPl56r_net_1\, C => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\, 
        Y => \I3.PULSE_46l9r_adt_net_146747_\);
    
    \I3.VDBi_57l2r_adt_net_1614_\ : OR2
      port map(A => \I3.VDBi_57l2r_adt_net_145218__net_1\, B => 
        \I3.VDBi_57l2r_adt_net_145227__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_1614__net_1\);
    
    \I2.DTE_21_1_IV_0_0L7R_1317\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855208__net_1\, 
        B => \I2.DT_TEMPl7r_net_1\, C => 
        \I2.DTE_21_1l7r_adt_net_38855_\, Y => 
        \I2.DTE_21_1l7r_adt_net_38870_\);
    
    \I2.ADE_4l6r\ : MUX2H
      port map(A => \I2.WOFFSETl7r\, B => \I2.ROFFSETl7r_net_1\, 
        S => NOESRAME_c, Y => \I2.ADE_4l6r_net_1\);
    
    \I1.SSTATEL2R_3004\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_289\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL2R_758\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855036_\ : BFR
      port map(A => \I2.PIPE1_DT_2_SQMUXA_ADT_NET_803__299\, Y
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855036__net_1\);
    
    \I3.VDBi_57l0r_adt_net_1621_\ : AO21
      port map(A => REGl32r, B => \I3.REGMAPl7r_net_1\, C => 
        \I3.REGMAPl8r_net_1\, Y => 
        \I3.VDBi_57l0r_adt_net_1621__net_1\);
    
    \I2.CRC32_812\ : MUX2L
      port map(A => \I2.CRC32l17r_net_1\, B => \I2.N_3934\, S => 
        \I2.N_2826_1_ADT_NET_794__331\, Y => \I2.CRC32_812_net_1\);
    
    \I2.OFFSET_37_9l6r\ : MUX2L
      port map(A => \REGl395r\, B => \REGl331r\, S => 
        \I2.PIPE7_DTL27R_76\, Y => \I2.N_705\);
    
    \I2.TEMPF_760\ : MUX2H
      port map(A => 
        \I2.TEMPF_adt_net_855740__adt_net_855896__net_1\, B => 
        \I2.N_2849\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.TEMPF_760_net_1\);
    
    \I2.INT_ERRAS_526\ : MUX2L
      port map(A => \I2.INT_ERRAS_net_1\, B => 
        \I2.INT_ERRAF1_net_1\, S => 
        \I2.N_3877_adt_net_855268__net_1\, Y => 
        \I2.INT_ERRAS_526_net_1\);
    
    \I1.REG_74_0_ivl374r\ : AO21
      port map(A => \REGl374r\, B => \I1.N_249\, C => 
        \I1.REG_74l374r_adt_net_113001_\, Y => \I1.REG_74l374r\);
    
    \I2.NWEN\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWEN_450_net_1\, SET => 
        CLEAR_STAT_i_0, Q => NWEN_c);
    
    \I1.PAGECNT_n4_0_0\ : OAI21
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_854520__net_1\, 
        B => \I1.N_394_i_i_0_i\, C => \I1.N_473\, Y => 
        \I1.PAGECNT_n4\);
    
    \I2.PIPE4_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl4r_net_1\);
    
    NPWON_pad : IB33
      port map(PAD => NPWON, Y => NPWON_c);
    
    \I5.SBYTE_66\ : MUX2H
      port map(A => \I5.SBYTEl1r_net_1\, B => \I5.N_16\, S => 
        \I5.N_406\, Y => \I5.SBYTE_66_net_1\);
    
    \I1.REG_74_0_IVL287R_1932\ : NOR2FT
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l287r_adt_net_122119_\);
    
    \I2.WOFFSET_834\ : MUX2L
      port map(A => \I2.WOFFSETl7r_Rd1__net_1\, B => 
        \I2.N_4250_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835308_Rd1__net_1\, Y
         => \I2.WOFFSETl7r\);
    
    \I2.UN1_NWPIPE7_2_1668\ : AND3
      port map(A => \I2.un1_NWPIPE7_2_adt_net_73604_\, B => 
        \I2.PIPE7_DTL25R_681\, C => \I2.PIPE7_DTl24r_net_1\, Y
         => \I2.un1_NWPIPE7_2_adt_net_73600_\);
    
    \I2.OFFSET_37_25l1r\ : MUX2L
      port map(A => \REGl254r\, B => \REGl190r\, S => 
        \I2.PIPE7_DTl27r_net_1\, Y => \I2.N_828\);
    
    \I3.VDBi_57_0_iv_0_0_a2l8r_941\ : NOR2
      port map(A => \I3.N_2015_120\, B => \I3.REGMAPL55R_782\, Y
         => \I3.N_2016_319\);
    
    \I2.L2TYPEl4r_1544\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_593_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL4R_651\);
    
    \I3.un57_reg_ads_0_a2_3_a3\ : NOR2
      port map(A => \I3.N_632\, B => \I3.N_581\, Y => 
        \I3.un57_reg_ads_0_a2_3_a3_net_1\);
    
    \I2.MIC_ERR_REGS_352\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl24r_net_1\, B => 
        \I2.MIC_ERR_REGSl23r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_352_net_1\);
    
    \I2.un21_pipe5_dt_3\ : XOR2
      port map(A => \I2.un21_pipe5_dt_1_net_1\, B => 
        \I2.un21_pipe5_dt_0_net_1\, Y => 
        \I2.un21_pipe5_dt_3_net_1\);
    
    \I3.VDBI_57_IV_0_0L2R_2264\ : AO21
      port map(A => \I3.N_2034_adt_net_854684__net_1\, B => 
        \I3.RAMDTSl2r_net_1\, C => 
        \I3.VDBi_57l2r_adt_net_145379_\, Y => 
        \I3.VDBi_57l2r_adt_net_145380_\);
    
    \I2.un6_tdcgdb1_3\ : XOR2
      port map(A => \I2.TDCl3r_net_1\, B => \I2.TDCDBSl27r_net_1\, 
        Y => \I2.un6_tdcgdb1_3_net_1\);
    
    \I2.PIPE8_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_535_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl7r_net_1\);
    
    \I5.SDAout_12_iv_0_a2\ : OR2FT
      port map(A => \I5.N_70\, B => \I5.N_150_adt_net_9847_\, Y
         => \I5.N_150\);
    
    \I2.resyn_0_I2_BITCNT_935\ : MUX2H
      port map(A => \I2.BITCNTl5r_net_1\, B => \I2.N_4326\, S => 
        \I2.BITCNTe\, Y => \I2.BITCNT_935\);
    
    \I2.un28_sram_empty_2_0\ : MUX2L
      port map(A => \I2.L2TYPEL12R_652\, B => \I2.L2TYPEL4R_651\, 
        S => \I2.RPAGEL15R_515\, Y => \I2.N_621\);
    
    \I2.PIPE7_DTL27R_2771\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_64\);
    
    \I2.RAMAD1_12l13r\ : MUX2L
      port map(A => \I2.TDCDASl24r_net_1\, B => 
        \I2.TDCDBSl24r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855184__net_1\, Y => 
        \I2.RAMAD1_12l13r_net_1\);
    
    \I1.REG_74_0_iv_0_0_a2l245r\ : NOR2
      port map(A => \I1.N_240\, B => \I1.N_254_196\, Y => 
        \I1.N_592\);
    
    \I2.DTOSl4r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl4r, Q => 
        \I2.DTOSl4r_net_1\);
    
    AMB_padl1r : IB33
      port map(PAD => AMB(1), Y => AMB_cl1r);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__2820\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__148\);
    
    \I3.VDBOFFB_30_IV_0L1R_2471\ : OR2
      port map(A => \I3.VDBoffb_30l1r_adt_net_162931_\, B => 
        \I3.VDBoffb_30l1r_adt_net_162932_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162937_\);
    
    \I2.un28_sram_empty_5_0\ : MUX2L
      port map(A => \I2.L2TYPEL14R_656\, B => \I2.L2TYPEL6R_655\, 
        S => \I2.RPAGEL15R_518\, Y => \I2.N_624\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_adt_net_803__net_1\, Y
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\);
    
    \I2.CHAINB_EN244_c_0_adt_net_855240_\ : BFR
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\, 
        Y => \I2.CHAINB_EN244_c_0_adt_net_855240__net_1\);
    
    \I2.PIPE9_DT_271\ : MUX2L
      port map(A => \I2.PIPE9_DTl2r_net_1\, B => 
        \I2.PIPE8_DTl2r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_271_net_1\);
    
    \I2.OFFSETl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_565_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl5r_net_1\);
    
    \I3.PIPEA_259\ : MUX2L
      port map(A => \I3.PIPEAl28r_net_1\, B => 
        \I3.PIPEA_8l28r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854652__net_1\, Y
         => \I3.PIPEA_259_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I6_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L12R_798\, B => 
        \I2.PIPE4_DTl6r_net_1\, Y => \I2.N_61_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I177_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl7r_adt_net_854552__adt_net_854948__net_1\, Y
         => \I2.ADD_21x21_fast_I177_Y_0\);
    
    \I2.UN1_STATE3_12_I_1710\ : OR2
      port map(A => \I2.STATE3_i_il10r\, B => \I2.STATE3_i_il12r\, 
        Y => \I2.N_2989_adt_net_92422_\);
    
    \I2.PIPE4_DTl5r_adt_net_854420_\ : BFR
      port map(A => \I2.PIPE4_DTl5r_net_1\, Y => 
        \I2.PIPE4_DTl5r_adt_net_854420__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I142_Y_0\ : XOR2
      port map(A => \I2.N_3537_i_i\, B => \I2.G_1_3\, Y => 
        \I2.ADD_18x18_fast_I142_Y_0\);
    
    \I1.REG_74_1_380_m8_i_0\ : OA21TTF
      port map(A => \I1.REG_74_1_396_m7_i_a5_0\, B => 
        \I1.REG_74_1_380_N_16\, C => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536__net_1\, 
        Y => \I1.REG_74_1_380_m8_i_0_0\);
    
    \I1.REG_0_sqmuxa_i_0_a4_1\ : NAND2
      port map(A => \I1.N_598_322\, B => 
        \I1.SSTATE_NS_IL5R_ADT_NET_107266__323\, Y => 
        \I1.N_435_1\);
    
    \I3.un6_asb_3_0_x2\ : XOR2FT
      port map(A => VAD_inl31r, B => GA_cl3r, Y => \I3.N_262_i_0\);
    
    \I2.INC_EVNT_NUM_759\ : AO21FTT
      port map(A => \I2.STATE2l1r_adt_net_855116__net_1\, B => 
        \I2.INC_EVNT_NUM_net_1\, C => 
        \I2.N_2864_0_adt_net_854268__net_1\, Y => 
        \I2.INC_EVNT_NUM_759_net_1\);
    
    \I2.REG_1_n7_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855788__net_1\, B
         => REGl39r, Y => \I2.REG_1_n7_0_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_4\ : AND2
      port map(A => \I2.RAMDT4L5R_821\, B => 
        \I2.N_140_0_adt_net_947__net_1\, Y => \I2.N_140\);
    
    \I2.FID_7_IVL2R_1729\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl2r_net_1\, 
        Y => \I2.FID_7l2r_adt_net_93351_\);
    
    \I2.PIPE9_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_283_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl14r_net_1\);
    
    \I2.TEMPF\ : DFFC
      port map(CLK => CLK_c, D => \I2.TEMPF_760_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TEMPF_net_1\);
    
    \I2.DTO_9_IVL14R_1145\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        B => \I2.N_126_i_0\, Y => \I2.DTO_9l14r_adt_net_32134_\);
    
    REGl261r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_162_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl261r\);
    
    \I2.DTE_cl_63l31r\ : DFFS
      port map(CLK => CLK_c, D => \I2.DTE_cl_63_870_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.DTE_cl_32l31r\);
    
    \I3.REG_1_294\ : MUX2L
      port map(A => VDB_inl12r, B => REGl113r, S => 
        \I3.N_318_adt_net_855884__net_1\, Y => \I3.REG_1_294_0\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2389\ : AND2
      port map(A => \REGl346r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        Y => \I3.VDBoffb_30l5r_adt_net_162144_\);
    
    \I3.PULSEl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_332_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl2r);
    
    \I1.REG_74_0_ivl356r\ : AO21
      port map(A => \REGl356r\, B => \I1.N_225\, C => 
        \I1.REG_74l356r_adt_net_115601_\, Y => 
        \I1.REG_74l356r_net_1\);
    
    \I2.RAMADl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l1r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl1r);
    
    \I2.DTE_21_1_IV_0L16R_1270\ : AND2
      port map(A => \I2.DT_TEMPl16r_net_1\, B => \I2.N_4038_233\, 
        Y => \I2.DTE_21_1l16r_adt_net_37825_\);
    
    \I1.REG_74_0_ivl331r\ : AO21
      port map(A => \REGl331r\, B => \I1.N_201\, C => 
        \I1.REG_74l331r_adt_net_118002_\, Y => \I1.REG_74l331r\);
    
    \I2.DTOSl27r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl27r, Q => 
        \I2.DTOSl27r_net_1\);
    
    \I2.PIPE5_DTl23r_1516\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_699_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL23R_623\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_2678\ : AND2
      port map(A => \I2.N_128_adt_net_54290_\, B => \I2.N_95\, Y
         => \I2.N525_adt_net_336000_\);
    
    \I2.RAMDT4L5R_3066\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_820\);
    
    \I2.SUB9_1_ADD_18x18_fast_I101_Y\ : AO21
      port map(A => \I2.N308\, B => \I2.N346_adt_net_4075__net_1\, 
        C => \I2.N307_1\, Y => \I2.N469\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I99_Y\ : AOI21FTT
      port map(A => \I2.N311_0\, B => \I2.N314\, C => \I2.N310_0\, 
        Y => \I2.N353\);
    
    \I2.CRC32_12_i_m2l13r\ : MUX2L
      port map(A => \I2.DT_TEMPl13r_net_1\, B => \I2.N_4048\, S
         => \I2.N_4667_1_ADT_NET_1046__35\, Y => \I2.N_3958_i_i\);
    
    \I2.RAMDT4L12R_2812\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_140\);
    
    \I2.I_1340_G_1\ : XOR2FT
      port map(A => \I2.OFFSETL5R_674\, B => \I2.SUB8l8r_net_1\, 
        Y => \I2.G_1_1\);
    
    \I2.TDCDBSl25r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl25r, Q => 
        \I2.TDCDBSl25r_net_1\);
    
    \I3.majority_0_reg_5_i_il0r\ : AO21
      port map(A => \I3.REG2l0r_net_1\, B => \I3.REG3l0r_net_1\, 
        C => \REGl0r_adt_net_53773_\, Y => REGl0r);
    
    \I2.N_587_adt_net_1201_\ : NAND3
      port map(A => \I2.PIPE7_DTL31R_502\, B => 
        \I2.PIPE7_DTl30r_net_1\, C => \I2.PIPE7_DT_i_0l33r\, Y
         => \I2.N_587_adt_net_1201__net_1\);
    
    \I2.ENDF_1139\ : DFFC
      port map(CLK => CLK_c, D => \I2.ENDF_712_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ENDF_401\);
    
    \I3.REG_1l157r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_205_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl157r\);
    
    \I2.DTE_21_1_IV_2L3R_1337\ : OAI21TTF
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_290\, B => 
        \I2.DT_SRAMl3r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39312_\, Y => 
        \I2.DTE_21_1_iv_2_il3r_adt_net_39313_\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I140_Y_0_O2_1_1545\ : 
        AOI21
      port map(A => \I2.PIPE4_DTl8r_adt_net_854556__net_1\, B => 
        \I2.PIPE4_DTL9R_846\, C => \I2.RAMDT4L5R_811\, Y => 
        \I2.N_74_i_0_i_adt_net_54331_\);
    
    \I3.EVREADi\ : DFFC
      port map(CLK => CLK_c, D => \I3.EVREADi_225_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => EVREAD);
    
    \I2.PIPE1_DT_42_1_IVL5R_1495\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855756__net_1\, B => 
        \I2.PIPE1_DT_30l5r_net_1\, C => 
        \I2.PIPE1_DT_42l5r_adt_net_51171_\, Y => 
        \I2.PIPE1_DT_42l5r_adt_net_51187_\);
    
    \I4.STATE1l2r\ : DFFS
      port map(CLK => CLK_c, D => \I4.STATE1_nsl0r_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I4.STATE1l2r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L7R_2358\ : AO21
      port map(A => \REGl300r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l7r_adt_net_161756_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161791_\);
    
    \I2.G_EVNT_NUM_n6_i_o2\ : AND2FT
      port map(A => \I2.N_4669_adt_net_855052__net_1\, B => 
        \I2.G_EVNT_NUMl5r_net_1\, Y => \I2.N_4672\);
    
    \I2.MIC_REG3_323\ : MUX2L
      port map(A => \I2.MIC_REG3l7r_net_1\, B => 
        \I2.MIC_REG3l6r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG3_323_net_1\);
    
    \I2.RAMAD1_12l14r\ : MUX2L
      port map(A => \I2.TDCDASl25r_net_1\, B => 
        \I2.TDCDBSl25r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855184__net_1\, Y => 
        \I2.RAMAD1_12l14r_net_1\);
    
    \I2.PIPE6_DT_478\ : MUX2H
      port map(A => \I2.PIPE5_DTl24r_net_1\, B => 
        \I2.PIPE6_DTl24r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_478_net_1\);
    
    \I1.PAGECNT_n3_0_0\ : OAI21
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_854520__net_1\, 
        B => \I1.N_393_i_i_0_i\, C => \I1.N_473\, Y => 
        \I1.PAGECNT_n3\);
    
    \I3.VDBI_57_0_IVL12R_2206\ : AO21
      port map(A => \I3.PIPEAl12r_net_1\, B => \I3.N_90_i_0_1\, C
         => \I3.VDBi_57l12r_adt_net_140988_\, Y => 
        \I3.VDBi_57l12r_adt_net_140997_\);
    
    REGl316r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_217_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl316r\);
    
    \I2.N507_adt_net_283110_\ : OA21
      port map(A => \I2.PIPE4_DTL11R_843\, B => 
        \I2.PIPE4_DTL12R_857\, C => \I2.RAMDT4L5R_815\, Y => 
        \I2.N507_adt_net_283110__net_1\);
    
    \I2.N_140_0_ADT_NET_947__2886\ : OR2
      port map(A => \I2.PIPE4_DTl5r_adt_net_854420__net_1\, B => 
        \I2.PIPE4_DTL6R_479\, Y => \I2.N_140_0_ADT_NET_947__327\);
    
    \I2.un1_tdc_res_24_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl406r, Y => 
        \I2.N_4605_i_0\);
    
    \I5.SDAOUT_12_IV_0_A2_918\ : OR3
      port map(A => \I5.sstate1l6r_net_1\, B => \I5.N_74\, C => 
        \I5.N_150_adt_net_9846_\, Y => \I5.N_150_adt_net_9847_\);
    
    \I2.CRC32_810\ : MUX2L
      port map(A => \I2.CRC32l15r_net_1\, B => \I2.N_3932\, S => 
        \I2.N_2826_1_ADT_NET_794__331\, Y => \I2.CRC32_810_net_1\);
    
    \I2.N_3_adt_net_940_\ : OR2
      port map(A => \I2.PIPE4_DTl6r_net_1\, B => 
        \I2.PIPE4_DTl7r_adt_net_854552__adt_net_854948__net_1\, Y
         => \I2.N_3_adt_net_940__net_1\);
    
    \I2.un1_DTE_1_sqmuxa_i_a6_0_a2_0_a2_1\ : NOR2
      port map(A => \I2.N_237\, B => \I2.N_4641\, Y => 
        \I2.N_2868_1\);
    
    \I2.PIPE5_DTl21r_1518\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_697_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL21R_625\);
    
    \I2.EVNT_NUM_102\ : NAND2FT
      port map(A => EV_RES_c, B => \I2.EVNT_NUMl11r_net_1\, Y => 
        \I2.N_1233\);
    
    \I2.END_CHAINA1_708\ : OR2FT
      port map(A => \I2.N_3273\, B => 
        \I2.END_CHAINA1_708_adt_net_53513_\, Y => 
        \I2.END_CHAINA1_708_net_1\);
    
    \I3.un146_reg_ads_0_a2_1_a2_0\ : OR3FFT
      port map(A => \I3.VASl2r_net_1\, B => \I3.N_548\, C => 
        \I3.N_555\, Y => \I3.N_641\);
    
    \I1.N_50_0_ADT_NET_1409__2868\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__541\, B => 
        \I1.N_50_0_ADT_NET_109751__256\, Y => 
        \I1.N_50_0_ADT_NET_1409__282\);
    
    \I2.STATE4l0r\ : DFFS
      port map(CLK => CLK_c, D => \I2.STATE4_ns_il2r_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.STATE4_il0r\);
    
    \I3.VDBoffb_58\ : OR3
      port map(A => \I3.VDBoffb_58_adt_net_162030_\, B => 
        \I3.VDBoffb_30l6r_adt_net_161989_\, C => 
        \I3.VDBoffb_30l6r_adt_net_161990_\, Y => 
        \I3.VDBoffb_58_net_1\);
    
    \I2.END_CHAINA1\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.END_CHAINA1_708_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.END_CHAINA1_net_1\);
    
    REGl333r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_234_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl333r\);
    
    \I3.PULSE_46_0_iv_0_0l6r\ : OR2FT
      port map(A => \I3.REG_1_sqmuxa_3\, B => 
        \I3.PULSE_46l6r_adt_net_147015_\, Y => \I3.PULSE_46l6r\);
    
    \I1.REG_1_144\ : MUX2H
      port map(A => \REGl243r\, B => \I1.REG_74l243r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_144_net_1\);
    
    \I2.STATE1l14r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_il4r_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.STATE1l14r_net_1\);
    
    \I3.VDBi_31l1r\ : NOR3
      port map(A => \I3.REGMAPl17r_adt_net_854292__net_1\, B => 
        \I3.REGMAPL14R_735\, C => \I3.REGMAPl11r_net_1\, Y => 
        \I3.VDBi_31l1r_adt_net_506111_\);
    
    \I2.MAJORITY_REG_I_0L1R_896\ : AOI21
      port map(A => \I2.MIC_REG3L1R_454\, B => 
        \I2.MIC_REG1L1R_455\, C => \I2.MIC_REG2L1R_536\, Y => 
        \I2.N_3877_adt_net_4725_\);
    
    \I2.STATE1_1_sqmuxa_3_0_a3\ : NAND3FFT
      port map(A => \I2.CHAINA_EN244_i_adt_net_855264__net_1\, B
         => \I2.TOKOUTAS_net_1\, C => \I2.STATE1l11r_net_1\, Y
         => \I2.STATE1_1_sqmuxa_3\);
    
    \I3.VDBi_40_1l14r\ : MUX2L
      port map(A => REGl131r, B => \I3.VDBi_31l14r_net_1\, S => 
        \I3.REGMAPl16r_net_1\, Y => \I3.N_352\);
    
    \I2.STATE4_ns_i_0_o2_0l1r\ : NOR2
      port map(A => \I2.L2AS_adt_net_855720__net_1\, B => 
        PULSEl2r, Y => \I2.N_4462\);
    
    LSRAM_FL_RADDRl2r : DFFC
      port map(CLK => CLK_c, D => \I4.LSRAM_FL_RADDR_11\, CLR => 
        CLEAR_STAT_i_0, Q => \LSRAM_FL_RADDRl2r\);
    
    \I1.REG_74_0_IVL299R_1919\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l299r_adt_net_120954_\);
    
    \I3.MBLTCYC_1161\ : DFFC
      port map(CLK => CLK_c, D => \I3.MBLTCYC_114_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.MBLTCYC_423\);
    
    \I1.REG_74_0_iv_0_0l245r\ : AO21
      port map(A => \REGl245r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l245r_adt_net_126207_\, Y => \I1.REG_74l245r\);
    
    \I2.DTE_21_1_IV_0L27R_1239\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.G_EVNT_NUMl11r_net_1\, 
        C => \I2.DTE_21_1l27r_adt_net_36860_\, Y => 
        \I2.DTE_21_1l27r_adt_net_36861_\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I108_Y_1659\ : AND2FT
      port map(A => \I2.SUB8l19r_net_1\, B => 
        \I2.N436_adt_net_1185__net_1\, Y => 
        \I2.N436_adt_net_70753_\);
    
    \I3.un21_reg_ads_0_a2_0_a3_1\ : NAND3FFT
      port map(A => \I3.WRITES_8\, B => 
        \I3.un60_reg_ads_3_adt_net_166295_\, C => 
        \I3.VASl1r_net_1\, Y => \I3.un60_reg_ads_3\);
    
    \I1.ISCK_0_SQMUXA_0_0_2076\ : AND3FFT
      port map(A => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854908__net_1\, B
         => \I1.sstatel4r_net_1\, C => \I1.N_628\, Y => 
        \I1.ISCK_0_sqmuxa_adt_net_134155_\);
    
    \I3.VDBOFFB_30_IV_0L6R_2367\ : AND2
      port map(A => \REGl355r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161938_\);
    
    \I1.sstatel0r\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_ns_il10r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel0r_net_1\);
    
    \I2.resyn_0_I2_FID_438\ : MUX2H
      port map(A => FID_cl22r, B => \I2.FID_7l22r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        Y => \I2.FID_438\);
    
    \I2.PIPE2_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl11r_net_1\);
    
    \I2.FIDl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_447\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl31r);
    
    \I3.PIPEB_88_2335\ : NOR2FT
      port map(A => \I3.PIPEBl9r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_88_adt_net_160335_\);
    
    \I2.PIPE8_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_548_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl20r_net_1\);
    
    N_1_I3_TCNT2_n6 : XOR2
      port map(A => \I3.TCNT2_i_0_il6r_net_1\, B => 
        \N_1.I3.TCNT2_c5\, Y => \N_1.I3.TCNT2_n6\);
    
    \I2.DTE_21_1_iv_0l5r\ : AO21
      port map(A => \I2.DTE_1l5r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\, C => 
        \I2.DTE_21_1l5r_adt_net_39101_\, Y => \I2.DTE_21_1l5r\);
    
    \I2.PIPE9_DTl29r_1562\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_298_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTL29R_669\);
    
    \I2.CRC32_12_i_0l10r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_249_i_i_0\, Y => 
        \I2.N_3927\);
    
    \I3.un196_reg_ads_0_a2_2_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_584\, Y => 
        \I3.un196_reg_ads_0_a2_2_a3_net_1\);
    
    \I1.REG_74_12_284_m10_i_0_0\ : AO21
      port map(A => \I1.REG_74_12_348_m9_i_adt_net_115429_\, B
         => \I1.REG_74_12_284_m10_i_o6_net_1\, C => 
        \I1.REG_74_12_284_m10_i_0_i_adt_net_121593_\, Y => 
        \I1.REG_74_12_284_m10_i_0_i\);
    
    \I2.WOFFSETl6r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl6r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl6r_Rd1__net_1\);
    
    \I1.REG_74_8_308_m9_i_x2\ : XOR2FT
      port map(A => \I1.PAGECNTl8r_net_1\, B => 
        \I1.REG_74_8_308_m6_e_net_1\, Y => 
        \I1.REG_74_8_308_N_6_i\);
    
    \I1.REG_74_0_ivl324r\ : AO21
      port map(A => \REGl324r\, B => \I1.N_193\, C => 
        \I1.REG_74l324r_adt_net_118701_\, Y => 
        \I1.REG_74l324r_net_1\);
    
    \I3.VDBoffa_46\ : OR3
      port map(A => \I3.VDBoffa_46_adt_net_164308_\, B => 
        \I3.VDBoffa_31l2r_adt_net_164269_\, C => 
        \I3.VDBoffa_31l2r_adt_net_164270_\, Y => 
        \I3.VDBoffa_46_net_1\);
    
    \I2.G_EVNT_NUM_n3_i_0_a2\ : NOR2FT
      port map(A => \I2.N_187\, B => \I2.G_EVNT_NUMl3r_net_1\, Y
         => \I2.N_317\);
    
    \I2.DTO_16_1_iv_0_o2_2tt_21_m3\ : AO21FTT
      port map(A => \I2.MIC_REG1l3r_adt_net_834596_Rd1__net_1\, B
         => \I2.DTO_16_1_iv_0_o2_2tt_21_N_8\, C => 
        \I2.DTO_16_1_iv_0_o2_2tt_21_m3_adt_net_27978_\, Y => 
        \I2.DTO_16_1_iv_0_o2_2tt_21_m3_net_1\);
    
    \I2.DTO_16_1_IV_0_0L16R_1135\ : AND2
      port map(A => \I2.DTO_1l16r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l16r_adt_net_31708_\);
    
    VDB_padl1r : IOB33PH
      port map(PAD => VDB(1), A => \I3.VDBml1r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl1r);
    
    \I3.VDBOFFB_30_IV_0L0R_2485\ : AO21
      port map(A => \REGl325r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l0r_adt_net_163090_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163122_\);
    
    \I3.STATE2l1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE2_nsl3r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I3.STATE2l1r_net_1\);
    
    \I2.un1_tdc_res_40_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl406r, Y => 
        \I2.N_4621_i_0\);
    
    \I3.PIPEA1l27r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_325_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l27r_net_1\);
    
    \I3.REGMAPL34R_2929\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un151_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL34R_446\);
    
    \I3.VDBoff_4_i_il7r\ : MUX2L
      port map(A => \I3.VDBoffbl7r_net_1\, B => 
        \I3.VDBoffal7r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_81\);
    
    \I3.PIPEB_81\ : AO21
      port map(A => DPR_cl2r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_81_adt_net_160629_\, Y => 
        \I3.PIPEB_81_net_1\);
    
    \I1.REG_74_0_IV_0_0L258R_1967\ : AND2
      port map(A => \FBOUTl5r\, B => \I1.N_596\, Y => 
        \I1.REG_74l258r_adt_net_124970_\);
    
    \I1.REG_74_0_ivl345r\ : AO21
      port map(A => \REGl345r\, B => \I1.N_217\, C => 
        \I1.REG_74l345r_adt_net_116584_\, Y => \I1.REG_74l345r\);
    
    \I1.REG_74_8_0_324_m9_i_x2\ : XOR2
      port map(A => \I1.PAGECNTL8R_457\, B => 
        \I1.REG_74_8_0_324_m6_e_net_1\, Y => 
        \I1.REG_74_8_0_N_6_i_i_0\);
    
    \I2.L2SERVl3r_1254\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_516\);
    
    \I2.BNC_IDl6r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_31_0\, CLR => 
        \I2.N_4623_i_0\, SET => \I2.N_4615_i_0\, Q => 
        \I2.BNC_IDl6r_net_1\);
    
    \I1.PAGECNT_320_adt_net_854872_\ : BFR
      port map(A => \I1.PAGECNT_320_net_1\, Y => 
        \I1.PAGECNT_320_adt_net_854872__net_1\);
    
    DTE_padl20r : IOB33PH
      port map(PAD => DTE(20), A => \I2.DTE_1l20r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl20r);
    
    \I2.REG_1l35r_1457\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n3_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL35R_564);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I140_Y_0_o2\ : AOI21
      port map(A => \I2.N_45_1_106\, B => 
        \I2.ADD_21x21_fast_I140_Y_0_a2_0_0_0\, C => 
        \I2.N_152_i_0_adt_net_502546_\, Y => \I2.N_70_0\);
    
    \I3.VADm_0_a3l23r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl23r_net_1\, Y => \I3.VADml23r\);
    
    \I2.SUB8l6r_1599\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_509_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8L6R_706\);
    
    \I5.REG_1_38\ : MUX2L
      port map(A => \I5.TEMPDATAl5r_net_1\, B => REGl425r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_38_net_1\);
    
    \I0.CLEAR_STATi_634\ : DFFC
      port map(CLK => CLK_c, D => \I0.CLEAR_STATi_4_net_1\, CLR
         => \I0.un12_clear_i\, Q => CLEAR_STAT_12);
    
    REGl254r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_155_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl254r\);
    
    \I2.PIPE1_DT_42_1_IVL14R_1437\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044__net_1\, 
        B => \I2.PIPE1_DT_12l14r_net_1\, Y => 
        \I2.PIPE1_DT_42l14r_adt_net_48948_\);
    
    \I5.SDAOUT_12_IV_0_919\ : AO21
      port map(A => \I5.sstate1l6r_net_1\, B => 
        \I5.SBYTEl7r_net_1\, C => \I5.sstate1l9r_net_1\, Y => 
        \I5.SDAout_12_adt_net_9914_\);
    
    \I2.DT_SRAM_0_i_m2l9r\ : MUX2L
      port map(A => \I2.PIPE10_DTl9r_net_1\, B => 
        \I2.PIPE5_DTl9r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854216__net_1\, Y => 
        \I2.N_4045\);
    
    \I2.FID_7_0_IVL31R_973\ : AND2
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl31r_net_1\, 
        Y => \I2.FID_7l31r_adt_net_18457_\);
    
    \I2.un2_evnt_word_I_65\ : AND2
      port map(A => \I2.WOFFSETl10r\, B => \I2.N_16_1\, Y => 
        \I2.N_9_1\);
    
    \I3.un1_NRDMEBi_2_sqmuxa_3_0\ : OAI21
      port map(A => \I3.N_203_adt_net_854976__net_1\, B => 
        DTEST_FIFO, C => \I3.STATE2l4r_net_1\, Y => 
        \I3.un1_NRDMEBi_2_sqmuxa_3_0_adt_net_153527_\);
    
    \I2.DTE_21_1_IV_0L5R_1325\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855120__net_1\, B => 
        \I2.EVNT_WORDl1r_net_1\, Y => 
        \I2.DTE_21_1l5r_adt_net_39083_\);
    
    \I3.END_PK_229\ : MUX2H
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854456__net_1\, B => 
        \I3.END_PK_net_1\, S => \I3.un1_STATE2_11\, Y => 
        \I3.END_PK_229_net_1\);
    
    \I2.STATE2l1r_adt_net_855132_\ : BFR
      port map(A => \I2.STATE2l1r\, Y => 
        \I2.STATE2l1r_adt_net_855132__net_1\);
    
    \I2.PIPE1_DT_42_0_ivl31r\ : OR2
      port map(A => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__169\, B => 
        \I2.PIPE1_DT_42l31r_adt_net_45041_\, Y => 
        \I2.PIPE1_DT_42l31r\);
    
    \I2.OFFSET_37_11l3r\ : MUX2L
      port map(A => \REGl376r\, B => \REGl312r\, S => 
        \I2.PIPE7_DTL27R_81\, Y => \I2.N_718\);
    
    \I2.PIPE10_DT_634\ : MUX2L
      port map(A => \I2.PIPE10_DTl29r_net_1\, B => 
        \I2.PIPE10_DT_17l29r\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_634_net_1\);
    
    \I2.DTO_16_1_iv_1l3r\ : AO21FTT
      port map(A => \I2.DTO_1l3r_net_1\, B => \I2.N_196_53\, C
         => \I2.DTO_16_1_iv_1l3r_adt_net_34608_\, Y => 
        \I2.DTO_16_1_iv_1l3r_net_1\);
    
    \I3.PIPEA_252\ : MUX2L
      port map(A => \I3.PIPEAl21r_net_1\, B => 
        \I3.PIPEA_8l21r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854660__net_1\, Y
         => \I3.PIPEA_252_net_1\);
    
    \I3.NRDMEBi_0_sqmuxa\ : OR2
      port map(A => \I3.N_1463_i_adt_net_1279__net_1\, B => 
        \I3.END_PK_879\, Y => \I3.NRDMEBi_0_sqmuxa_net_1\);
    
    REGl373r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_274_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl373r\);
    
    \I3.VDBil2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_342_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil2r_net_1\);
    
    \I1.REG_74_0_ivl402r\ : AO21
      port map(A => \REGl402r\, B => \I1.N_273\, C => 
        \I1.REG_74l402r_adt_net_109928_\, Y => \I1.REG_74l402r\);
    
    \I1.REG_74_0_ivl218r\ : AO21
      port map(A => \REGl218r\, B => \I1.N_89_165\, C => 
        \I1.REG_74l218r_adt_net_128948_\, Y => \I1.REG_74l218r\);
    
    \I2.WOFFSET_13_i_o2l1r\ : AND2FT
      port map(A => \I2.WPAGEe\, B => \I2.N_4262_adt_net_39852_\, 
        Y => \I2.N_4262\);
    
    \I1.REG_74_0_IVL332R_1884\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l332r_adt_net_117916_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I3_G0N_0_o3\ : NAND2
      port map(A => \I2.RAMDT4L3R_765\, B => 
        \I2.PIPE4_DTl3r_adt_net_854548__net_1\, Y => \I2.N_17\);
    
    \I2.SUB9l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_571_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l3r_net_1\);
    
    \I2.CRC32_12_i_m2l15r\ : MUX2H
      port map(A => \I2.DT_SRAMl15r_net_1\, B => 
        \I2.DT_TEMPl15r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854432__net_1\, Y => 
        \I2.N_3960_i_i\);
    
    FID_padl4r : OB33PH
      port map(PAD => FID(4), A => FID_cl4r);
    
    \I2.PIPE1_DT_42_0l27r\ : NAND2FT
      port map(A => \I2.PIPE1_DT_1_sqmuxa\, B => \I2.N_3273\, Y
         => \I2.PIPE1_DT_42_0l27r_net_1\);
    
    \I3.REGMAPl14r_1625\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un57_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL14R_732\);
    
    VAD_padl24r : OTB33PH
      port map(PAD => VAD(24), A => \I3.VADml24r\, EN => 
        NOEAD_c_i_0);
    
    \I1.REG_74_3_i_a2l172r\ : NAND2FT
      port map(A => \I1.N_1370_adt_net_112317_\, B => 
        \I1.N_273_6_i_0\, Y => \I1.N_1370\);
    
    \I2.N475_adt_net_442369_\ : OA21
      port map(A => \I2.N296_0\, B => \I2.N479_adt_net_642266_\, 
        C => \I2.N285\, Y => \I2.N475_adt_net_442369__net_1\);
    
    \I3.VDBI_57_0_IVL31R_2139\ : AND2
      port map(A => \I3.PIPEAl31r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l31r_adt_net_137838_\);
    
    \I2.WOFFSET_837\ : MUX2L
      port map(A => \I2.WOFFSETl10r_Rd1__net_1\, B => 
        \I2.N_4253_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835304_Rd1__net_1\, Y
         => \I2.WOFFSETl10r\);
    
    \I1.ISI_0_SQMUXA_1_0_I_2074\ : NOR2FT
      port map(A => \I1.N_346\, B => \I1.N_368\, Y => 
        \I1.N_1375_adt_net_134063_\);
    
    \I2.DTO_cl_0_sqmuxa_0_adt_net_855200_\ : BFR
      port map(A => \I2.DTO_cl_0_sqmuxa_0\, Y => 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855200__net_1\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__2834\ : NOR3FFT
      port map(A => \I2.END_EVNT5_406\, B => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\, C => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m3_net_1\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__183\);
    
    \I1.PAGECNT_318_adt_net_854856_\ : BFR
      port map(A => \I1.PAGECNT_318_net_1\, Y => 
        \I1.PAGECNT_318_adt_net_854856__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I142_Y\ : XOR2
      port map(A => \I2.N313_0\, B => 
        \I2.ADD_18x18_fast_I142_Y_0\, Y => \I2.SUB9_1l5r\);
    
    \I3.VDBI_57_IVL4R_2253\ : AO21
      port map(A => 
        \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344__net_1\, 
        B => \I3.VDBi_52l4r_net_1\, C => 
        \I3.VDBi_57l4r_adt_net_144440_\, Y => 
        \I3.VDBi_57l4r_adt_net_144441_\);
    
    \I2.SUB9_0_sqmuxa_0_a2_0_0\ : NOR3FFT
      port map(A => \I2.SUB9_0_sqmuxa_0_adt_net_20771_\, B => 
        \I2.PIPE8_DTl31r_net_1\, C => \I2.PIPE8_DTl29r_net_1\, Y
         => \I2.SUB9_0_sqmuxa_0\);
    
    \I2.PIPE2_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl3r_net_1\);
    
    \I1.REG_74_0_ivl375r\ : AO21
      port map(A => \REGl375r\, B => \I1.N_249\, C => 
        \I1.REG_74l375r_adt_net_112915_\, Y => \I1.REG_74l375r\);
    
    \I2.CRC32_12_i_0_m2l19r\ : MUX2L
      port map(A => \I2.DT_TEMPl19r_net_1\, B => 
        \I2.DT_SRAMl19r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854196__net_1\, Y => 
        \I2.N_229_i_i\);
    
    \I2.STATE1l18r\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_o2_0l0r_net_1\, SET => CLEAR_STAT_i_0, Q
         => \I2.STATE1l18r_net_1\);
    
    \I3.VDBoffb_30_iv_0l6r\ : AND2
      port map(A => \REGl371r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161934_\);
    
    \I2.PIPE1_DT_42_1_ivl29r\ : OR2
      port map(A => \I2.PIPE1_DT_42l29r_adt_net_45838_\, B => 
        \I2.PIPE1_DT_42l29r_adt_net_45839_\, Y => 
        \I2.PIPE1_DT_42l29r\);
    
    \I2.OFFSET_37_13l3r\ : MUX2L
      port map(A => \I2.N_726\, B => \I2.N_710\, S => 
        \I2.PIPE7_DTL25R_685\, Y => \I2.N_734\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855428_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__22\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\);
    
    \I2.DTE_2_1l10r\ : XOR2
      port map(A => \I2.CRC32l30r_net_1\, B => 
        \I2.DTE_2_1_0l10r_net_1\, Y => \I2.DTE_2_1l10r_net_1\);
    
    \I2.G_EVNT_NUM_m_1_i_0_o2l8r\ : OR2FT
      port map(A => \I2.N_176_I_157\, B => \I2.N_4641_55\, Y => 
        \I2.N_223\);
    
    \I3.STATE1l6r_1623\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl4r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL6R_730\);
    
    \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__2824\ : OR3
      port map(A => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_N_20_i\, B
         => \I2.DTE_cl_0_sqmuxa_2_adt_net_20059__net_1\, C => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20061__net_1\, Y => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\);
    
    \I1.REG_3_sqmuxa_0_a2_0\ : NAND2FT
      port map(A => \I1.PAGECNTl9r_net_1\, B => 
        \I1.N_238_Rd1__adt_net_854884__net_1\, Y => \I1.N_254\);
    
    \I2.PIPE6_DT_458\ : MUX2H
      port map(A => \I2.PIPE5_DTl4r_net_1\, B => 
        \I2.PIPE6_DTl4r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_458_net_1\);
    
    \I1.PAGECNT_n6_i_i_a2_851\ : AND2FT
      port map(A => \I1.PAGECNTl6r_net_1\, B => 
        \I1.PAGECNTL5R_311\, Y => \I1.N_590_229\);
    
    \I2.FID_419\ : MUX2H
      port map(A => FID_cl3r, B => \I2.FID_7l3r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        Y => \I2.FID_419_net_1\);
    
    \I2.TOKENA_TIMOUT\ : DFFC
      port map(CLK => CLK_c, D => \I2.TOKENA_TIMOUT_2_net_1\, CLR
         => \I2.un6_clear_stat_i\, Q => \I2.TOKENA_TIMOUT_net_1\);
    
    \I1.BYTECNTlde_i_a2_i_m2\ : MUX2H
      port map(A => \I1.SSTATEL6R_714\, B => \I1.SSTATEL4R_715\, 
        S => \I1.BYTECNTl8r_net_1\, Y => \I1.N_332\);
    
    \I5.AIR_WDATA_59\ : MUX2L
      port map(A => \I5.AIR_WDATAl9r_net_1\, B => 
        \I5.AIR_WDATA_9l9r_net_1\, S => \I5.N_461\, Y => 
        \I5.AIR_WDATA_59_net_1\);
    
    \I3.REG2l2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG2_143_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l2r_net_1\);
    
    \I3.VDBi_354\ : MUX2L
      port map(A => \I3.VDBil14r_net_1\, B => \I3.VDBi_57l14r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_354_net_1\);
    
    \I3.PIPEA_8l8r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854480__net_1\, B => 
        \I3.N_217\, Y => \I3.PIPEA_8l8r_net_1\);
    
    \I2.NWPIPE5_1470\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE4_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE5_577\);
    
    \I3.VDBml9r\ : MUX2L
      port map(A => \I3.VDBil9r_net_1\, B => \I3.N_151\, S => 
        \I3.SINGCYC_881\, Y => \I3.VDBml9r_net_1\);
    
    \I1.REG_74_0_ivl290r\ : AO21
      port map(A => \REGl290r\, B => \I1.N_161\, C => 
        \I1.REG_74l290r_adt_net_121861_\, Y => \I1.REG_74l290r\);
    
    \I2.PIPE1_DT_42_1_IVL3R_1504\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl35r_net_1\, C => 
        \I2.PIPE1_DT_42l3r_adt_net_51617_\, Y => 
        \I2.PIPE1_DT_42l3r_adt_net_51634_\);
    
    \I3.VDBI_20_IVL8R_2219\ : AND2FT
      port map(A => \I3.N_1907\, B => \I3.VDBi_16l8r_net_1\, Y
         => \I3.VDBi_20l8r_adt_net_142456_\);
    
    \I3.un151_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_583\, Y => 
        \I3.un151_reg_ads_0_a2_0_a3_net_1\);
    
    \I3.PIPEA1_329\ : MUX2L
      port map(A => \I3.PIPEA1l31r_net_1\, B => 
        \I3.PIPEA1_12l31r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, Y => 
        \I3.PIPEA1_329_net_1\);
    
    \I3.REG_1l7r\ : AO21
      port map(A => \I3.REG1l7r_net_1\, B => \I3.REG2l7r_net_1\, 
        C => \REGl7r_adt_net_8466_\, Y => REGl7r);
    
    VAD_padl31r : IOB33PH
      port map(PAD => VAD(31), A => \I3.VADml31r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl31r);
    
    \I2.DTO_16_1_IV_0_O2_0L12R_1156\ : AND2FT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl12r_net_1\, Y => \I2.N_3966_adt_net_32562_\);
    
    \I1.REG_1_299\ : MUX2H
      port map(A => \REGl398r\, B => \I1.REG_74l398r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y => 
        \I1.REG_1_299_net_1\);
    
    \I3.VDBi_366\ : MUX2L
      port map(A => \I3.VDBil26r_net_1\, B => \I3.VDBi_57l26r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_366_net_1\);
    
    \I3.PIPEA1l2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_300_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l2r_net_1\);
    
    \I1.PAGECNTl6r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_321_adt_net_854880__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTl6r_net_1\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2524\ : AO21
      port map(A => \REGl187r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.N_2070_adt_net_163498_\, Y => 
        \I3.N_2070_adt_net_163505_\);
    
    \I2.TOKINBi_326\ : OA21TTF
      port map(A => TOKINB_c, B => \I2.STATE1l8r_net_1\, C => 
        \I2.STATE1l7r_net_1\, Y => \I2.TOKINBi_326_net_1\);
    
    NOELUT_pad : OB33PH
      port map(PAD => NOELUT, A => NOELUT_c);
    
    \I2.PIPE6_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_482_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl28r_net_1\);
    
    \I2.ADO_3l9r\ : MUX2L
      port map(A => \I2.WOFFSETl10r\, B => \I2.ROFFSETl10r_net_1\, 
        S => NOESRAME_C_243, Y => \I2.ADO_3l9r_net_1\);
    
    \I2.un2_tdcgdb1_0_adt_net_21805_\ : OR2
      port map(A => \I2.TDCDBSl31r_net_1\, B => 
        \I2.TDCDBSl29r_net_1\, Y => 
        \I2.un2_tdcgdb1_0_adt_net_21805__net_1\);
    
    REGl221r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_122_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl221r\);
    
    \I5.SDAnoe\ : DFFS
      port map(CLK => CLK_c, D => \I5.SDAnoe_83_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SDAnoe_net_1\);
    
    RAMAD_padl6r : OB33PH
      port map(PAD => RAMAD(6), A => RAMAD_cl6r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I62_Y\ : AO21
      port map(A => \I2.N258_0_adt_net_854936__net_1\, B => 
        \I2.N312_0_adt_net_86450_\, C => 
        \I2.N312_0_adt_net_86445_\, Y => \I2.N312_0\);
    
    \I2.DTOSl0r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl0r, Q => 
        \I2.DTOSl0r_net_1\);
    
    PAF_c_i : INV
      port map(A => PAF_c, Y => PAF_c_i_0);
    
    \I3.TCNT4l3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT4_385_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT4l3r_net_1\);
    
    \I1.BITCNT_n2_i_i_o2_646\ : AND2
      port map(A => \I1.BITCNTL0R_18\, B => \I1.BITCNTl1r_net_1\, 
        Y => \I1.N_324_24\);
    
    \I2.SUB9l16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_584_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l16r_net_1\);
    
    \I1.REG_74l236r\ : OR3
      port map(A => \I1.N_201_9\, B => \I1.REG_10_sqmuxa\, C => 
        \I1.N_113_adt_net_3714__net_1\, Y => \I1.N_105\);
    
    \I2.RESYN_0_I2_LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_950\ : AO21
      port map(A => \I2.PIPE4_DTl23r_net_1\, B => 
        \I2.N_4524_adt_net_16596_\, C => 
        \I2.N_4524_adt_net_16803_\, Y => 
        \I2.N_4524_adt_net_16804_\);
    
    \I2.L2TYPE_4_i_o2_0l6r\ : AND2FT
      port map(A => \I2.L2ARRl3r_net_1\, B => \I2.L2ARRl2r_net_1\, 
        Y => \I2.N_4460\);
    
    \I1.N_1377_adt_net_106750_\ : AO21FTT
      port map(A => \I1.N_310_Rd1__net_1\, B => \I1.N_590\, C => 
        \I1.N_238_Rd1__adt_net_854884__net_1\, Y => 
        \I1.N_1377_adt_net_106750__net_1\);
    
    \I2.RAMADl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l5r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl5r);
    
    \I2.DTO_9_ivl22r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl22r_net_1\, 
        C => \I2.DTO_9l22r_adt_net_30294_\, Y => \I2.DTO_9l22r\);
    
    \I2.DTO_1l7r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l7r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l7r_Rd1__net_1\);
    
    \I2.TDCDBSl23r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl23r, Q => 
        \I2.TDCDBSl23r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I145_Y\ : XOR2
      port map(A => \I2.N469\, B => \I2.ADD_18x18_fast_I145_Y_0\, 
        Y => \I2.SUB9_1l8r\);
    
    \I2.FID_7_0_IVL12R_967\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl12r_net_1\, 
        Y => \I2.FID_7l12r_adt_net_18175_\);
    
    \I3.VDBoffbl6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_58_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl6r_net_1\);
    
    \I5.AIR_START\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_START_16_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_START_net_1\);
    
    \I5.SENS_ADDR_1_sqmuxa\ : OR2
      port map(A => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\, B
         => \I5.SENS_ADDR_1_sqmuxa_adt_net_14344_\, Y => 
        \I5.SENS_ADDR_1_sqmuxa_net_1\);
    
    \I2.DTE_21_1_IV_0L24R_1247\ : AO21FTT
      port map(A => \I2.DTE_cl_0_sqmuxa_2_0\, B => \I2.N_4194\, C
         => \I2.DTE_21_1l24r_adt_net_37173_\, Y => 
        \I2.DTE_21_1l24r_adt_net_37174_\);
    
    \I3.REG_1_ml77r\ : AND2
      port map(A => REGl77r, B => 
        \I3.REGMAPl9r_adt_net_854304__net_1\, Y => 
        \I3.VDBi_20l29r\);
    
    \I3.REG2_148\ : MUX2L
      port map(A => VDB_inl7r, B => \I3.REG2l7r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG2_148_net_1\);
    
    \I2.MIC_REG2l6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_315_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2l6r_net_1\);
    
    \I2.ADO_3l13r\ : MUX2H
      port map(A => \I2.RPAGEl13r\, B => \I2.WPAGEl13r_net_1\, S
         => NOESRAME_c, Y => \I2.ADO_3l13r_net_1\);
    
    \I2.FID_7_0_IVL29R_978\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl77r, C => 
        \I2.FID_7l29r_adt_net_18645_\, Y => 
        \I2.FID_7l29r_adt_net_18653_\);
    
    \I1.PAGECNT_n1_0_0\ : OAI21
      port map(A => \I1.un1_sbyte13_1_i_1\, B => \I1.N_388_i_0_i\, 
        C => \I1.N_473_205\, Y => \I1.PAGECNT_n1\);
    
    \I3.TCNT_0_sqmuxa_0_a2_0_a3\ : NOR3FFT
      port map(A => \I3.REGMAPl51r_net_1\, B => \I3.WRITES_8\, C
         => \I3.N_276\, Y => \I3.TCNT_0_sqmuxa\);
    
    \I2.DTO_1l28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_902_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l28r_net_1\);
    
    \I2.CHB_DATA8\ : DFFC
      port map(CLK => CLK_c, D => \I2.CHB_DATA8_503_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.CHB_DATA8_net_1\);
    
    \I1.sstate_ns_1_iv_0_0l7r\ : OR2FT
      port map(A => \I1.N_485\, B => 
        \I1.sstate_nsl7r_adt_net_107578_\, Y => \I1.sstate_nsl7r\);
    
    \I2.PIPE10_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_617_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl12r_net_1\);
    
    \I3.TICKil0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.un6_tcnt1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TICKl0r);
    
    \I2.DTE_21_1_IVL15R_1273\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855128__net_1\, B => 
        \I2.EVNT_WORDl11r_net_1\, Y => 
        \I2.DTE_21_1l15r_adt_net_37935_\);
    
    \I2.un7_bnc_id_1_I_30\ : AND2
      port map(A => \I2.BNC_IDl5r_net_1\, B => \I2.N_34_0\, Y => 
        \I2.N_29_0\);
    
    \I1.REG_1_296\ : MUX2H
      port map(A => \REGl395r\, B => \I1.REG_74l395r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y => 
        \I1.REG_1_296_net_1\);
    
    \I1.N_50_0_adt_net_1409_\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__200\, B => 
        \I1.N_50_0_adt_net_109751__net_1\, Y => 
        \I1.N_50_0_adt_net_1409__net_1\);
    
    \I2.DTE_21_1_IV_2L2R_1338\ : AND2
      port map(A => GA_cl2r, B => 
        \I2.STATE2l1r_adt_net_855120__net_1\, Y => 
        \I2.DTE_21_1_iv_2_il2r_adt_net_39443_\);
    
    \I2.CHAIN_ERR_DIS_448\ : OR2FT
      port map(A => \I2.N_3510\, B => 
        \I2.CHAIN_ERR_DIS_448_adt_net_92599_\, Y => 
        \I2.CHAIN_ERR_DIS_448_net_1\);
    
    \I2.TRGARRl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGARR_3l2r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGARRl2r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I155_Y_0\ : XOR2FT
      port map(A => \I2.N_3562_i\, B => \I2.SUB8l19r_net_1\, Y
         => \I2.ADD_18x18_fast_I155_Y_0\);
    
    \I1.PAGECNTl4r_adt_net_835120_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.PAGECNT_323_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNTl4r_adt_net_835120_Rd1__net_1\);
    
    \I2.STATE1_nsl6r\ : NAND3FTT
      port map(A => \I2.STATE1_nsl6r_adt_net_23511_\, B => 
        \I2.STATE1_1_sqmuxa_3\, C => \I2.un1_STATE1_28\, Y => 
        \I2.STATE1_nsl6r_net_1\);
    
    VDB_padl28r : IOB33PH
      port map(PAD => VDB(28), A => \I3.VDBml28r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl28r);
    
    \I2.DTO_16_1_IV_0L20R_1119\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854616__net_1\, 
        B => \I2.DT_TEMPl20r_net_1\, C => 
        \I2.DTO_16_1l20r_adt_net_30786_\, Y => 
        \I2.DTO_16_1l20r_adt_net_30792_\);
    
    \I2.MTDCRESA\ : DFFC
      port map(CLK => CLK_c, D => \I2.MTDCRESA_378_net_1\, CLR
         => \I2.un9_clear_stat_i\, Q => MTDCRESA_c);
    
    \I2.PIPE1_DTl7r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_734_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl7r_net_1\);
    
    \I3.PIPEA1l20r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_318_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l20r_net_1\);
    
    \I2.G_EVNT_NUM_929\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl5r_net_1\, B => \I2.N_4345\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_929_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I113_un1_Y\ : AND3
      port map(A => \I2.N346_adt_net_4075__net_1\, B => 
        \I2.N463_adt_net_70886_\, C => \I2.N331\, Y => 
        \I2.I113_un1_Y\);
    
    \I2.BNCID_VECT_tile_DOUTl0r\ : MUX2L
      port map(A => \I2.DIN_REG1_0l0r\, B => \I2.DOUT_TMP_0l0r\, 
        S => \I2.N_13\, Y => \I2.BNCID_VECTrxl0r\);
    
    \I2.L2TYPE_4_il5r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4447_adt_net_68073_\, C => 
        \I2.N_4447_adt_net_68116_\, Y => \I2.N_4447\);
    
    \I3.PIPEA1_12l0r\ : AND2
      port map(A => DPR_cl0r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854488__net_1\, Y => 
        \I3.PIPEA1_12l0r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL28R_1362\ : AND3
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, B => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, C
         => \I2.TDCDBSl28r_net_1\, Y => 
        \I2.PIPE1_DT_42l28r_adt_net_45931_\);
    
    \I2.BNCID_VECT_tile_I_1\ : RAM256x9SA
      port map(DO8 => OPEN, DO7 => \I2.DOUT_TMPl7r\, DO6 => 
        \I2.DOUT_TMPl6r\, DO5 => \I2.DOUT_TMPl5r\, DO4 => 
        \I2.DOUT_TMPl4r\, DO3 => \I2.DOUT_TMP_0l3r\, DO2 => 
        \I2.DOUT_TMP_0l2r\, DO1 => \I2.DOUT_TMP_0l1r\, DO0 => 
        \I2.DOUT_TMP_0l0r\, WPE => OPEN, RPE => OPEN, DOS => OPEN, 
        WADDR7 => \GND\, WADDR6 => \GND\, WADDR5 => \GND\, WADDR4
         => \GND\, WADDR3 => \I2.TRGARRl3r_net_1\, WADDR2 => 
        \I2.TRGARRl2r_net_1\, WADDR1 => \I2.TRGARRl1r_net_1\, 
        WADDR0 => \I2.TRGARRl0r_net_1\, RADDR7 => \GND\, RADDR6
         => \GND\, RADDR5 => \GND\, RADDR4 => \GND\, RADDR3 => 
        \I2.TRGSERVl3r_net_1\, RADDR2 => \I2.TRGSERVL2R_584\, 
        RADDR1 => \I2.TRGSERVl1r_net_1\, RADDR0 => 
        \I2.TRGSERVl0r_net_1\, DI8 => \GND\, DI7 => 
        \I2.BNC_IDl7r_net_1\, DI6 => \I2.BNC_IDl6r_net_1\, DI5
         => \I2.BNC_IDl5r_net_1\, DI4 => \I2.BNC_IDl4r_net_1\, 
        DI3 => \I2.BNC_IDl3r_net_1\, DI2 => \I2.BNC_IDl2r_net_1\, 
        DI1 => \I2.BNC_IDl1r_net_1\, DI0 => \I2.BNC_IDl0r_net_1\, 
        WRB => \I2.TDCTRG_c_i_0\, RDB => \GND\, WBLKB => \GND\, 
        RBLKB => \GND\, PARODD => \VCC\, WCLKS => CLK_c, DIS => 
        \VCC\);
    
    \I2.STATE3l13r\ : DFFS
      port map(CLK => CLK_c, D => \GND\, SET => CLEAR_STAT_i_0, Q
         => \I2.STATE3l13r_net_1\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3\ : AO21
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__806\, B => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_a5_2_i_adt_net_2404__net_1\, C
         => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__161\, 
        Y => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_net_1\);
    
    \I2.OFFSET_37_21l3r\ : MUX2L
      port map(A => \I2.N_790\, B => \I2.N_766\, S => 
        \I2.PIPE7_DTL25R_685\, Y => \I2.N_798\);
    
    \I2.DTO_16_1_IVL15R_1141\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.DTE_2_1l15r_net_1\, Y
         => \I2.DTO_16_1l15r_adt_net_31956_\);
    
    \I3.VDBI_20_IVL10R_2212\ : AND2
      port map(A => REGl58r, B => 
        \I3.REGMAPl9r_adt_net_854320__net_1\, Y => 
        \I3.VDBi_20l10r_adt_net_141609_\);
    
    \I3.un146_reg_ads_0_a2_1_a2\ : NAND2FT
      port map(A => \I3.VASl5r_net_1\, B => \I3.VASl3r_net_1\, Y
         => \I3.N_551\);
    
    \I1.REG_74_0_1l332r\ : NOR3FFT
      port map(A => \I1.N_57_9_i\, B => \I1.REG_74_1L268R_187\, C
         => \I1.N_73_10\, Y => \I1.REG_74_0l332r\);
    
    \I2.SRAM_EVNT_n1\ : XOR2
      port map(A => \I2.N_3825\, B => \I2.SRAM_EVNT_n1_0_net_1\, 
        Y => \I2.SRAM_EVNT_n1_net_1\);
    
    \I2.RESYN_0_I2_LSRAM_RADDRI_1_SQMUXA_0_A4_I_O2_947\ : 
        OAI21TTF
      port map(A => \I2.PIPE4_DTl22r_net_1\, B => \I2.N_2330_tz\, 
        C => \I2.N_4524_adt_net_16740_\, Y => 
        \I2.N_4524_adt_net_16701_\);
    
    \I2.L2TYPEl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_590_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_i_0_il1r\);
    
    \I2.PIPE1_DT_42_1_IVL2R_1509\ : AND2FT
      port map(A => \I2.N_3279_0_adt_net_855232__net_1\, B => 
        \I2.MIC_ERR_REGSl2r_net_1\, Y => 
        \I2.PIPE1_DT_42l2r_adt_net_51829_\);
    
    \I2.ADOl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl4r);
    
    \I2.RAMDT4l3r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl3r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l3r_net_1\);
    
    \I3.REG3_128\ : MUX2L
      port map(A => VDB_inl3r, B => \I3.REG3l3r_net_1\, S => 
        \I3.REG3_0_sqmuxa\, Y => \I3.REG3_128_net_1\);
    
    \I1.sstate_ns_0_iv_0_i_m2l3r\ : MUX2L
      port map(A => \I1.sstatel7r_net_1\, B => 
        \I1.sstatel8r_net_1\, S => 
        \I1.N_321_adt_net_855540__net_1\, Y => \I1.N_420_i\);
    
    \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35789_\ : AND2
      port map(A => \I2.STATE2l5r_net_1\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35702__net_1\, Y => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35789__net_1\);
    
    \I1.REG_74_12_284_m10_i_o6\ : AND2FT
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854396__net_1\, 
        B => \I1.REG_74_1_380_N_16\, Y => 
        \I1.REG_74_12_284_m10_i_o6_net_1\);
    
    \I2.WOFFSET_829\ : MUX2L
      port map(A => \I2.WOFFSETl2r_Rd1__net_1\, B => 
        \I2.N_4245_Rd1__net_1\, S => 
        \I2.N_2828_ADT_NET_1062__ADT_NET_835312_RD1__379\, Y => 
        \I2.WOFFSETl2r\);
    
    \I2.DTE_1l15r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l15r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l15r_Rd1__net_1\);
    
    \I2.PIPE1_DT_42_1_IVL23R_1379\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, B => 
        \I2.TDCDBSl23r_net_1\, C => 
        \I2.PIPE1_DT_42l23r_adt_net_46639_\, Y => 
        \I2.PIPE1_DT_42l23r_adt_net_46654_\);
    
    \I2.STATE1_ns_il14r\ : OA21
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855244__net_1\, 
        B => \I2.END_CHAINB1_net_1\, C => \I2.N_158\, Y => 
        \I2.STATE1_ns_il14r_net_1\);
    
    \I1.REG_74_0_ivl343r\ : AO21
      port map(A => \REGl343r\, B => \I1.N_217\, C => 
        \I1.REG_74l343r_adt_net_116756_\, Y => \I1.REG_74l343r\);
    
    \I3.PIPEA1_12l5r\ : AND2
      port map(A => DPR_cl5r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854508__net_1\, Y => 
        \I3.PIPEA1_12l5r_net_1\);
    
    \I2.BNCID_VECTrff_11\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_11_254_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_11\);
    
    \I1.REG_74_0_ivl325r\ : AO21
      port map(A => \REGl325r\, B => \I1.N_201\, C => 
        \I1.REG_74l325r_adt_net_118518_\, Y => \I1.REG_74l325r\);
    
    \I2.un1_end_flush_9_1_adt_net_1193_\ : OR2
      port map(A => END_FLUSH_559, B => \I2.un1_NWPIPE5_1_i\, Y
         => \I2.un1_end_flush_9_1_adt_net_1193__net_1\);
    
    \I2.PIPE4_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl12r_net_1\);
    
    \I2.DTOSl5r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl5r, Q => 
        \I2.DTOSl5r_net_1\);
    
    \I3.PULSE_46_0_IV_I_IL4R_2293\ : AND2
      port map(A => PULSEL4R_15, B => 
        \I3.N_311_adt_net_854752__net_1\, Y => 
        \I3.N_55_adt_net_147183_\);
    
    \I1.REG_74_0_ivl233r\ : AO21
      port map(A => \REGl233r\, B => \I1.N_105\, C => 
        \I1.REG_74l233r_adt_net_127366_\, Y => \I1.REG_74l233r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I186_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_800\, B => 
        \I2.PIPE4_DTl16r_net_1\, Y => 
        \I2.ADD_21x21_fast_I186_Y_0_0\);
    
    \I2.BNCID_VECTrff_12_253_0\ : AO21
      port map(A => \I2.BNCID_VECTwa12_1_net_1\, B => 
        \I2.BNCID_VECTrff_12_253_0_a2_0\, C => 
        \I2.BNCID_VECTro_12\, Y => 
        \I2.BNCID_VECTrff_12_253_0_net_1\);
    
    REGl240r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_141_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl240r\);
    
    \I5.sstate1se_5_0_0_m2\ : MUX2H
      port map(A => \I5.sstate1l7r_net_1\, B => 
        \I5.sstate1l8r_net_1\, S => TICKl0r, Y => 
        \I5.sstate1_ns_el6r\);
    
    TDCDB_padl18r : IB33
      port map(PAD => TDCDB(18), Y => TDCDB_cl18r);
    
    \I3.STATE1_0l8r_1158\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl2r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL8R_420\);
    
    \I3.VDBOFFA_31_IV_0L7R_2495\ : AND2
      port map(A => \REGl220r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.VDBoffa_31l7r_adt_net_163276_\);
    
    \I1.REG_74_0_IV_I_A2L199R_2035\ : AND2
      port map(A => \REGl199r\, B => \I1.N_182_i\, Y => 
        \I1.N_1338_adt_net_130619_\);
    
    TDCDA_padl24r : IB33
      port map(PAD => TDCDA(24), Y => TDCDA_cl24r);
    
    \I2.OFFSET_37_23l3r\ : MUX2L
      port map(A => \REGl272r\, B => \REGl208r\, S => 
        \I2.PIPE7_DTL27R_90\, Y => \I2.N_814\);
    
    \I3.NRDMEBI_2_SQMUXA_I_0_O3_2300\ : NOR3
      port map(A => NOEAD_c, B => \I3.N_281_255\, C => 
        \I3.END_PK_net_1\, Y => \I3.N_297_adt_net_147649_\);
    
    \I3.VDBi_20_ivl14r\ : AO21
      port map(A => REGl62r, B => 
        \I3.REGMAPl9r_adt_net_854316__net_1\, C => 
        \I3.VDBi_20l14r_adt_net_140054_\, Y => \I3.VDBi_20l14r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I182_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_801\, B => 
        \I2.PIPE4_DTl12r_net_1\, Y => 
        \I2.ADD_21x21_fast_I182_Y_0_0\);
    
    \I2.CRC32_12_il3r\ : OA21
      port map(A => 
        \I2.N_4667_1_adt_net_1046__adt_net_854424__net_1\, B => 
        \I2.CRC32_2l3r_net_1\, C => \I2.N_3920_adt_net_43068_\, Y
         => \I2.N_3920\);
    
    \I2.SUB9_1_ADD_18x18_fast_I98_Y\ : NAND2FT
      port map(A => \I2.N460_adt_net_70355_\, B => \I2.N336\, Y
         => \I2.N460\);
    
    \I2.N_4540_i_0_o2\ : AND2FT
      port map(A => \I2.PIPE5_DTL23R_624\, B => 
        \I2.PIPE5_DTL21R_893\, Y => \I2.N_4673\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I189_Y\ : XOR2FT
      port map(A => \I2.N498\, B => \I2.ADD_21x21_fast_I189_Y_0\, 
        Y => \I2.un27_pipe5_dt0l19r\);
    
    \I2.PIPE1_DT_42_1_IVL21R_1389\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, B => 
        \I2.TDCDBSl21r_net_1\, C => 
        \I2.PIPE1_DT_42l21r_adt_net_46859_\, Y => 
        \I2.PIPE1_DT_42l21r_adt_net_46874_\);
    
    \I2.un7_tdcgda1_2\ : XOR2
      port map(A => \I2.TDCDASl26r_net_1\, B => \I2.TDCl2r_net_1\, 
        Y => \I2.un7_tdcgda1_2_i_i\);
    
    \I2.PIPE8_DT_16_0l14r\ : MUX2H
      port map(A => \I2.PIPE8_DTl14r_net_1\, B => 
        \I2.PIPE7_DTl14r_net_1\, S => 
        \I2.N_565_0_adt_net_855736__net_1\, Y => \I2.N_580\);
    
    \I3.STATE1_ILLEGAL_2133\ : AO21
      port map(A => 
        \I3.STATE1_ipl3r_adt_net_854364__adt_net_855344__net_1\, 
        B => \I3.N_1186_adt_net_1488__net_1\, C => 
        \I3.N_1193_ip_adt_net_136555_\, Y => 
        \I3.N_1193_ip_adt_net_136556_\);
    
    \I2.DTO_16_1_iv_0l13r\ : OR2
      port map(A => \I2.DTO_16_1l13r_adt_net_32395_\, B => 
        \I2.DTO_16_1l13r_adt_net_32396_\, Y => \I2.DTO_16_1l13r\);
    
    \I2.STATE2l1r_adt_net_855116_\ : BFR
      port map(A => \I2.STATE2l1r_adt_net_855120__net_1\, Y => 
        \I2.STATE2l1r_adt_net_855116__net_1\);
    
    \I2.CRC32l14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_809_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l14r_net_1\);
    
    \I1.REG_1_298\ : MUX2H
      port map(A => \REGl397r\, B => \I1.REG_74l397r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y => 
        \I1.REG_1_298_net_1\);
    
    \I2.PIPE6_DT_461\ : MUX2H
      port map(A => \I2.PIPE5_DTl7r_net_1\, B => 
        \I2.PIPE6_DTl7r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_461_net_1\);
    
    \I2.DTO_16_1_IVL11R_1168\ : AO21
      port map(A => \I2.DTO_1l11r\, B => \I2.N_196\, C => 
        \I2.DTO_16_1l11r_adt_net_32864_\, Y => 
        \I2.DTO_16_1l11r_adt_net_32880_\);
    
    \I5.un1_AIR_PULSE_0_sqmuxa_i_a3\ : OR2
      port map(A => \I5.N_463\, B => \I5.N_480\, Y => \I5.N_479\);
    
    \I2.REG_1_c13_i_a2_0\ : AND2FT
      port map(A => REGl45r, B => \I2.N_136_1\, Y => \I2.N_138\);
    
    \I2.DTO_16_1l4r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l4r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l4r_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L0R_2620\ : AND2
      port map(A => \REGl229r\, B => \I3.REGMAPl26r_net_1\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164602_\);
    
    \I3.VDBm_i_i_m2l5r\ : MUX2L
      port map(A => \I3.VDBil5r_net_1\, B => \I3.N_284\, S => 
        \I3.SINGCYC_net_1\, Y => VDBm_i_i_m2l5r);
    
    \I2.un1_TOKENA_CNT_I_1\ : AND2
      port map(A => TICKL0R_557, B => \I2.TOKENA_CNTl0r_net_1\, Y
         => \I2.DWACT_ADD_CI_0_TMP_2l0r\);
    
    \I1.REG_74_0_ivl373r\ : AO21
      port map(A => \REGl373r\, B => \I1.N_249\, C => 
        \I1.REG_74l373r_adt_net_113087_\, Y => \I1.REG_74l373r\);
    
    \I1.BYTECNTl2r_adt_net_855020_\ : BFR
      port map(A => \I1.BYTECNTl2r_net_1\, Y => 
        \I1.BYTECNTl2r_adt_net_855020__net_1\);
    
    \I2.L2ARRl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_944_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRl0r_net_1\);
    
    \I2.DTE_21_1l24r_adt_net_37175_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.DTE_21_1l24r_adt_net_37175_\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.DTE_21_1l24r_adt_net_37175_Rd1__net_1\);
    
    \I2.REG_1l44r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n12_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl44r);
    
    \I1.REG_74_0_ivl295r\ : AO21
      port map(A => \REGl295r\, B => \I1.N_169\, C => 
        \I1.REG_74l295r_adt_net_121298_\, Y => \I1.REG_74l295r\);
    
    \I3.REG_1l70r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_171_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl70r);
    
    \I2.LSRAM_IN_402\ : MUX2L
      port map(A => \I2.PIPE5_DTl18r_net_1\, B => 
        \I2.LSRAM_INl18r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_402_net_1\);
    
    \I2.DT_SRAMl30r\ : MUX2L
      port map(A => \I2.N_898\, B => \I2.PIPE2_DTl30r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl30r_net_1\);
    
    \I1.COMMAND_0_sqmuxa_1_0_0_a2_i\ : OR2
      port map(A => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854908__net_1\, B
         => \I1.N_606_Rd1__net_1\, Y => \I1.N_1384\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_A2_2_1544\ : AND2
      port map(A => \I2.N_64\, B => \I2.N_89\, Y => 
        \I2.N_128_adt_net_54291_\);
    
    \I2.UN1_STATE1_38_0_O2_1526\ : OA21FTT
      port map(A => \I2.ERR_WORDS_RDY_net_1\, B => \I2.N_3277\, C
         => \I2.STATE1l14r_net_1\, Y => 
        \I2.N_3292_adt_net_52393_\);
    
    \I2.DTO_16_1_IV_0L8R_1181\ : AO21
      port map(A => \I2.N_457\, B => \I2.DTE_2_1l8r_net_1\, C => 
        \I2.DTO_16_1l8r_adt_net_33480_\, Y => 
        \I2.DTO_16_1l8r_adt_net_33489_\);
    
    TDCDA_padl13r : IB33
      port map(PAD => TDCDA(13), Y => TDCDA_cl13r);
    
    \I3.UN5_NOE16RI_0_I_O2_898\ : AND3FFT
      port map(A => DS0B_c, B => DS1B_c, C => \I3.WRITES_8\, Y
         => \I3.N_290_adt_net_4891_\);
    
    \I1.REG_74l228r\ : OAI21
      port map(A => \I1.REG_74_2_4_il228r\, B => 
        \I1.REG_74_2_3_il228r\, C => 
        \I1.REG_74_12_220_m9_i_net_1\, Y => \I1.N_97\);
    
    TDCDB_padl27r : IB33
      port map(PAD => TDCDB(27), Y => TDCDB_cl27r);
    
    \I2.BNCID_VECTror_8_tz\ : AOI21
      port map(A => \I2.BNCID_VECTra14_1_net_1\, B => 
        \I2.BNCID_VECTro_10\, C => \I2.BNCID_VECTria_11_0_i\, Y
         => \I2.BNCID_VECTror_8_tz_i_adt_net_48039_\);
    
    \I1.REG_74_1l276r_809\ : NOR3FFT
      port map(A => \I1.N_273_5_i\, B => 
        \I1.N_273_6_i_0_adt_net_854796__net_1\, C => 
        \I1.N_201_9_189\, Y => \I1.REG_74_1L268R_187\);
    
    \I2.PIPE7_DTl30r_adt_net_855172_\ : BFR
      port map(A => \I2.PIPE7_DTl30r_net_1\, Y => 
        \I2.PIPE7_DTl30r_adt_net_855172__net_1\);
    
    \I2.ADOl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l5r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl5r);
    
    \I2.DTE_21_1_IV_2L2R_1340\ : OAI21TTF
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_290\, B => 
        \I2.N_4193\, C => \I2.DTE_21_1_iv_2_il2r_adt_net_39452_\, 
        Y => \I2.DTE_21_1_iv_2_il2r_adt_net_39453_\);
    
    REGl337r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_238_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl337r\);
    
    \I5.DATA_12l13r\ : MUX2L
      port map(A => REGl130r, B => \I5.SBYTEl5r_net_1\, S => 
        \I5.DATA_1_sqmuxa_2\, Y => \I5.DATA_12l13r_net_1\);
    
    REGl174r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_75_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl174r\);
    
    \I3.PIPEA_8_0l28r\ : MUX2L
      port map(A => DPR_cl28r, B => \I3.PIPEA1l28r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855356__net_1\, Y => \I3.N_237\);
    
    \I2.TEMPF_7_i_a6\ : NAND2FT
      port map(A => \I2.STATE2l5r_net_1\, B => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, Y => 
        \I2.N_2849\);
    
    \I2.PIPE1_DT_42_1_IVL13R_1447\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\, B => 
        \I2.PIPE1_DT_30l13r_net_1\, C => 
        \I2.PIPE1_DT_42l13r_adt_net_49195_\, Y => 
        \I2.PIPE1_DT_42l13r_adt_net_49211_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_o2_728\ : AND3FFT
      port map(A => \I2.N_3_0_adt_net_1070__net_1\, B => 
        \I2.N_95_0\, C => \I2.N_45_1_adt_net_271427_\, Y => 
        \I2.N_45_1_106\);
    
    \I2.PIPE5_DTl30r_1515\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_706_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL30R_622\);
    
    \I2.REG_1_n10_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855788__net_1\, B
         => REG_i_0_il42r, Y => \I2.REG_1_n10_0_net_1\);
    
    \I3.PIPEA1l22r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_320_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l22r_net_1\);
    
    \I2.FIDl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_429\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl13r);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2276\ : AND2
      port map(A => \I3.N_2046\, B => \I3.REGl133r\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146424_\);
    
    FID_padl8r : OB33PH
      port map(PAD => FID(8), A => FID_cl8r);
    
    \I2.DTO_1_892\ : MUX2L
      port map(A => \I2.DTO_1l18r_Rd1__net_1\, B => 
        \I2.DTO_16_1l18r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834764_Rd1__net_1\, Y
         => \I2.DTO_1l18r\);
    
    \I2.BNCID_VECTrff_8_257_0\ : AO21
      port map(A => \I2.BNCID_VECTwa12_1_net_1\, B => 
        \I2.BNCID_VECTrff_8_257_0_a2_0\, C => \I2.BNCID_VECTro_8\, 
        Y => \I2.BNCID_VECTrff_8_257_0_net_1\);
    
    \I3.VDBoffb_56\ : OR3
      port map(A => \I3.VDBoffb_56_adt_net_162410_\, B => 
        \I3.VDBoffb_30l4r_adt_net_162369_\, C => 
        \I3.VDBoffb_30l4r_adt_net_162370_\, Y => 
        \I3.VDBoffb_56_net_1\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854452_\ : BFR
      port map(A => \I3.N_243_4_adt_net_1290__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\);
    
    \I3.VDBi_57l7r_adt_net_143017_\ : AND2
      port map(A => REGl413r, B => \I3.REGMAPl55r_net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_143017__net_1\);
    
    \I2.DT_TEMPl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_785_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl24r_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2393\ : AO21
      port map(A => \REGl386r\, B => \I3.REGMAP_i_0_il45r_net_1\, 
        C => \I3.VDBoffb_30l5r_adt_net_162132_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162170_\);
    
    \I2.TDCDBSl30r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl30r, Q => 
        \I2.TDCDBSl30r_net_1\);
    
    DTE_padl25r : IOB33PH
      port map(PAD => DTE(25), A => \I2.DTE_1l25r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl25r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I68_Y\ : AO21
      port map(A => \I2.N245\, B => \I2.N249_0\, C => 
        \I2.N316_i_i_adt_net_86582_\, Y => \I2.N318\);
    
    \I3.UN15_TCNT4_2645\ : AND3FFT
      port map(A => \I3.TCNT4l1r_net_1\, B => 
        \I3.TCNT4_i_0_il2r_net_1\, C => 
        \I3.un15_tcnt4_adt_net_165650_\, Y => 
        \I3.un15_tcnt4_adt_net_165652_\);
    
    \I5.TEMPDATA_77\ : MUX2L
      port map(A => \I5.TEMPDATAl3r_net_1\, B => REGl128r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_77_net_1\);
    
    \I3.REG_1_153\ : MUX2L
      port map(A => VDB_inl4r, B => REGl52r, S => 
        \I3.N_1935_adt_net_855332__net_1\, Y => \I3.REG_1_153_0\);
    
    \I2.DTE_21_1_IV_0_0L7R_1318\ : OR3
      port map(A => \I2.DTO_16_1l7r_adt_net_33728_\, B => 
        \I2.DTE_21_1l7r_adt_net_38863_\, C => 
        \I2.DTE_21_1l7r_adt_net_38870_\, Y => 
        \I2.DTE_21_1l7r_adt_net_38872_\);
    
    \I2.TOKENB_TIMOUT\ : DFFC
      port map(CLK => CLK_c, D => \I2.TOKENB_TIMOUT_2\, CLR => 
        \I2.un12_clear_stat_i\, Q => \I2.TOKENB_TIMOUT_i_i\);
    
    \I2.MIC_REG1_307\ : MUX2L
      port map(A => \I2.MIC_REG1l7r_net_1\, B => 
        \I2.MIC_REG1_i_il6r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG1_307_net_1\);
    
    \I3.VDBi_351\ : MUX2L
      port map(A => \I3.VDBil11r_net_1\, B => \I3.VDBi_57l11r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__116\, Y => 
        \I3.VDBi_351_net_1\);
    
    \I2.WREi_8_i_i_a2\ : AOI21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.N_2838_i_0\, C
         => \I2.WREi_8_i_i_a2_1_net_1\, Y => \I2.N_4203\);
    
    \I3.VDBi_31l26r\ : MUX2L
      port map(A => \I3.REGl159r\, B => \I3.VDBi_20l26r\, S => 
        \I3.REGMAPl17r_adt_net_854284__net_1\, Y => 
        \I3.VDBi_31l26r_net_1\);
    
    \I3.VDBi_23l1r_adt_net_145541_\ : OAI21FTF
      port map(A => REGl33r, B => \I3.N_2033\, C => 
        \I3.VDBi_23l1r_adt_net_145526__net_1\, Y => 
        \I3.VDBi_23l1r_adt_net_145541__net_1\);
    
    \I2.SUB8l9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_512_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l9r_net_1\);
    
    \I2.REG_0l3r_adt_net_848__adt_net_854204_\ : BFR
      port map(A => \I2.REG_0l3r_adt_net_848__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__adt_net_854204__net_1\);
    
    \I2.G_EVNT_NUM_n6_i\ : NOR3
      port map(A => EV_RES_C_569, B => \I2.N_280\, C => 
        \I2.N_198\, Y => \I2.N_4638\);
    
    \I2.CHAINA_ERRS\ : DFFC
      port map(CLK => CLK_c, D => \I2.CHAINA_ERRS_524_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.CHAINA_ERRS_net_1\);
    
    \I2.RAMDT4L5R_3065\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_819\);
    
    REGl260r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_161_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl260r\);
    
    \I3.REGMAPl37r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un166_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl37r_net_1\);
    
    \I3.REG2l0r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG2_141_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l0r_net_1\);
    
    \I3.REG1l4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG1_137_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l4r_net_1\);
    
    \I5.BITCNT_n0_i_a2\ : AND2FT
      port map(A => \I5.N_73\, B => \I5.N_94\, Y => \I5.N_144\);
    
    \I3.VDBI_57_IV_0_0L7R_2231\ : AO21
      port map(A => \I3.N_2034_adt_net_854684__net_1\, B => 
        \I3.RAMDTSl7r_net_1\, C => 
        \I3.VDBi_57l7r_adt_net_143110_\, Y => 
        \I3.VDBi_57l7r_adt_net_143111_\);
    
    \I1.N_127_i_0_a4\ : OR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835132_RD1__884\, B
         => \I1.N_299_adt_net_833868_Rd1__net_1\, Y => 
        \I1.N_127_i\);
    
    \I3.STATE1_ILLEGAL_2129\ : AO21
      port map(A => \I3.STATE1_ipl7r\, B => 
        \I3.N_1174_adt_net_1495__net_1\, C => 
        \I3.N_1193_ip_adt_net_136551_\, Y => 
        \I3.N_1193_ip_adt_net_136552_\);
    
    \I2.EVNT_NUM_c7\ : AND2
      port map(A => \I2.EVNT_NUMl7r_net_1\, B => 
        \I2.EVNT_NUM_c6_net_1\, Y => \I2.EVNT_NUM_c7_net_1\);
    
    \I2.INT_ERRAF1_494\ : OAI21TTF
      port map(A => \I2.N_3877_adt_net_855268__net_1\, B => 
        INT_ERRA_c, C => \I2.INT_ERRAF1_494_adt_net_90420_\, Y
         => \I2.INT_ERRAF1_494_net_1\);
    
    \I3.PIPEA_8_0l19r\ : MUX2L
      port map(A => DPR_cl19r, B => \I3.PIPEA1l19r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855360__net_1\, Y => \I3.N_228\);
    
    \I2.STATE3_ns_il11r\ : NOR2
      port map(A => \I2.STATE3_0_sqmuxa_1_0\, B => \I2.N_3019\, Y
         => \I2.STATE3_ns_il11r_net_1\);
    
    \I2.DTO_16_1_IV_0L5R_1194\ : AND2FT
      port map(A => \I2.N_223_156\, B => \I2.DTE_2_1l5r_net_1\, Y
         => \I2.DTO_16_1l5r_adt_net_34192_\);
    
    \I3.REG3l0r_1638\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG3_125_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3L0R_745\);
    
    \I2.FID_7_0_IVL17R_957\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl17r_net_1\, 
        Y => \I2.FID_7l17r_adt_net_17705_\);
    
    NWRLUT_pad : OB33PH
      port map(PAD => NWRLUT, A => NWRLUT_c);
    
    \I3.VDBI_57_0_IV_0_0L15R_2186\ : AO21
      port map(A => REGl132r, B => \I3.N_2058\, C => 
        \I3.VDBi_57l15r_adt_net_139961_\, Y => 
        \I3.VDBi_57l15r_adt_net_139970_\);
    
    \I1.REG_74_0_IV_I_A2_IL205R_2029\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_6_sqmuxa_adt_net_854708__net_1\, Y => 
        \I1.N_280_adt_net_130103_\);
    
    \I3.PIPEA_8_0l12r\ : MUX2L
      port map(A => DPR_cl12r, B => \I3.PIPEA1l12r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855352__net_1\, Y => \I3.N_221\);
    
    \I1.REG_1_180\ : MUX2H
      port map(A => \REGl279r\, B => \I1.REG_74l279r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\, Y => 
        \I1.REG_1_180_net_1\);
    
    \I2.OFFSET_37_14l3r\ : MUX2L
      port map(A => \I2.N_734\, B => \I2.N_686\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_742\);
    
    \I2.DTO_16_1_IV_0_1L2R_1207\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.DTO_9_ivl2r\, C => 
        \I2.DTO_16_1_iv_0_1l2r_adt_net_34862_\, Y => 
        \I2.DTO_16_1_iv_0_1l2r_adt_net_34868_\);
    
    \I1.REG_74_0_iv_0_0l247r\ : AO21
      port map(A => \REGl247r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l247r_adt_net_126035_\, Y => \I1.REG_74l247r\);
    
    \I2.PIPE1_DTl12r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_739_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl12r_net_1\);
    
    \I2.N291_adt_net_4302_\ : OR2
      port map(A => \I2.SUB8l15r_net_1\, B => \I2.SUB8l14r_net_1\, 
        Y => \I2.N291_adt_net_4302__net_1\);
    
    \I2.RAMAD_4_0l16r\ : MUX2H
      port map(A => \I2.RAMAD1l16r_net_1\, B => RAMAD_VMEl16r, S
         => \REG_i_il5r_adt_net_855552__net_1\, Y => \I2.N_543\);
    
    \I2.PIPE5_DT_6_0l6r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l6r\, B => 
        \I2.un27_pipe5_dt0l6r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1075\);
    
    \I2.DT_TEMP_790\ : MUX2H
      port map(A => \I2.DT_TEMPl29r_net_1\, B => 
        \I2.DT_TEMP_7l29r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_790_net_1\);
    
    DTO_padl19r : IOB33PH
      port map(PAD => DTO(19), A => \I2.DTO_1l19r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl19r);
    
    \I2.un7_tdcgda1_1\ : XOR2
      port map(A => \I2.TDCDASl25r_net_1\, B => \I2.TDCl1r_net_1\, 
        Y => \I2.un7_tdcgda1_1_i_i\);
    
    \I2.PIPE1_DT_739\ : MUX2L
      port map(A => \I2.PIPE1_DTl12r_net_1\, B => 
        \I2.PIPE1_DT_42l12r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854576__net_1\, 
        Y => \I2.PIPE1_DT_739_net_1\);
    
    \I2.RAMDT4L7R_2926\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl7r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L7R_443\);
    
    \I3.TCNT4_c1\ : AND2
      port map(A => \I3.TCNT4_i_0_il0r_net_1\, B => 
        \I3.TCNT4l1r_net_1\, Y => \I3.TCNT4_c1_net_1\);
    
    \I2.TDCDBSl10r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl10r, Q => 
        \I2.TDCDBSl10r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2548\ : AND2
      port map(A => \REGl233r\, B => \I3.REGMAPl26r_net_1\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163842_\);
    
    \I3.RAMAD_VMEl10r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_34_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl10r);
    
    \I2.MIC_REG1_302\ : MUX2H
      port map(A => \I2.MIC_REG1l1r_net_1\, B => 
        \I2.MIC_REG1l2r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG1_302_net_1\);
    
    \I3.VDBI_20_IVL4R_2702\ : AO21
      port map(A => REGl52r, B => 
        \I3.REGMAPl9r_adt_net_854320__net_1\, C => 
        \I3.VDBi_20l4r_adt_net_414879_\, Y => 
        \I3.VDBi_20l4r_adt_net_514155_\);
    
    \I2.DTO_16_1_IVL28R_1076\ : AOI21
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.DTO_9_iv_ml28r_adt_net_857__net_1\, C => 
        \I2.DT_SRAM_i_m_0l28r_net_1\, Y => 
        \I2.DTO_16_1_ivl28r_adt_net_28982_\);
    
    \I2.resyn_0_I2_FID_437\ : MUX2H
      port map(A => FID_cl21r, B => \I2.FID_7l21r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        Y => \I2.FID_437\);
    
    WRITEB_pad : IB33
      port map(PAD => WRITEB, Y => WRITEB_c);
    
    \I3.VDBi_20_ivl8r\ : AO21
      port map(A => REGl56r, B => 
        \I3.REGMAPl9r_adt_net_854316__net_1\, C => 
        \I3.VDBi_20l8r_adt_net_142456_\, Y => \I3.VDBi_20l8r\);
    
    \I2.DTO_16_1_IV_0L17R_1132\ : AO21
      port map(A => \I2.G_EVNT_NUMl1r_net_1\, B => \I2.N_457\, C
         => \I2.DTO_16_1l17r_adt_net_31520_\, Y => 
        \I2.DTO_16_1l17r_adt_net_31531_\);
    
    \I2.CRC32l26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_821_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l26r_net_1\);
    
    \I4.UN2_END_TDC_1_930\ : OR2
      port map(A => LEAD_FLAGl5r, B => LEAD_FLAGl4r, Y => 
        \I4.un2_end_tdc_1_adt_net_15219_\);
    
    \I2.DTO_16_1_IV_0_O2L8R_1177\ : AND2FT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl8r_net_1\, Y => \I2.N_3967_adt_net_33418_\);
    
    REGl377r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_278_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl377r\);
    
    ADO_padl14r : OB33PH
      port map(PAD => ADO(14), A => ADO_cl14r);
    
    \I2.STATE3l12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3l13r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE3_i_il12r\);
    
    \I4.END_FLUSH_1453\ : DFFC
      port map(CLK => CLK_c, D => \I4.END_FLUSH_2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => END_FLUSH_560);
    
    \I3.VDBi_20_ivl12r\ : AO21
      port map(A => \I3.N_280\, B => 
        \I3.VDBi_20l12r_adt_net_140770_\, C => 
        \I3.VDBi_20l12r_adt_net_140765_\, Y => \I3.VDBi_20l12r\);
    
    \I3.PIPEA1_12l23r\ : AND2
      port map(A => DPR_cl23r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854496__net_1\, Y => 
        \I3.PIPEA1_12l23r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2434\ : AO21
      port map(A => \REGl392r\, B => \I3.REGMAP_i_il46r_net_1\, C
         => \I3.VDBoffb_30l3r_adt_net_162548_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162555_\);
    
    \I1.REG_74_0_IVL325R_1891\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l325r_adt_net_118518_\);
    
    \I2.DTO_16_1_IVL22R_1108\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854616__net_1\, 
        B => \I2.DT_TEMPl22r_net_1\, C => 
        \I2.DTO_16_1l22r_adt_net_30352_\, Y => 
        \I2.DTO_16_1l22r_adt_net_30360_\);
    
    \I1.REG_1_239\ : MUX2H
      port map(A => \REGl338r\, B => \I1.REG_74l338r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\, Y => 
        \I1.REG_1_239_net_1\);
    
    \I2.DTO_1_874\ : MUX2L
      port map(A => \I2.DTO_1l0r_net_1\, B => \I2.DTO_16_1_ivl0r\, 
        S => \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => 
        \I2.DTO_1_874_net_1\);
    
    ADO_padl7r : OB33PH
      port map(PAD => ADO(7), A => ADO_cl7r);
    
    \I3.VDBI_10_I_M2L5R_2239\ : AND2FT
      port map(A => \I2.N_3876_adt_net_855256__net_1\, B => 
        \I3.REGMAPL2R_737\, Y => \I3.N_283_adt_net_143528_\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855504_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__294\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\);
    
    \I3.TCNT1l2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT1_n2_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT1l2r_net_1\);
    
    \I2.DTO_16_1_IV_0L4R_1199\ : AND2
      port map(A => \I2.N_4671_adt_net_854600__net_1\, B => 
        \I2.DT_TEMPl4r_net_1\, Y => 
        \I2.DTO_16_1l4r_adt_net_34376_\);
    
    \I1.REG_1_142\ : MUX2H
      port map(A => \REGl241r\, B => \I1.REG_74l241r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_142_net_1\);
    
    \I1.PAGECNT_326\ : MUX2H
      port map(A => \I1.PAGECNTl1r_adt_net_834904_Rd1__net_1\, B
         => \I1.PAGECNT_n1\, S => 
        \I1.PAGECNTe_adt_net_854896__net_1\, Y => 
        \I1.PAGECNT_326_net_1\);
    
    \I2.PIPE9_DT_285\ : MUX2L
      port map(A => \I2.PIPE9_DTl16r_net_1\, B => 
        \I2.PIPE8_DTl16r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_285_net_1\);
    
    \I2.CRC32_12_i_x2l4r\ : XOR2FT
      port map(A => \I2.CRC32l4r_net_1\, B => \I2.N_3955_i_i\, Y
         => \I2.N_118_i_i_0\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855416_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__321\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\);
    
    \I1.REG_1_66\ : MUX2H
      port map(A => \REGl165r\, B => \I1.REG_74l165r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, Y => 
        \I1.REG_1_66_net_1\);
    
    \I3.REGMAP_I_0_A2L52R_2089\ : NOR2
      port map(A => \I3.REGMAPl4r_net_1\, B => 
        \I3.REGMAP_i_0_il15r\, Y => \I3.N_638_adt_net_134637_\);
    
    \I1.REG_74_0_IVL241R_1985\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_10_sqmuxa_adt_net_854716__net_1\, Y => 
        \I1.REG_74l241r_adt_net_126641_\);
    
    \I2.DTO_cl_0_sqmuxa_0_adt_net_855208_\ : BFR
      port map(A => \I2.DTO_cl_0_sqmuxa_0\, Y => 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855208__net_1\);
    
    \I1.REG_74_0_ivl323r\ : AO21
      port map(A => \REGl323r\, B => \I1.N_193\, C => 
        \I1.REG_74l323r_adt_net_118787_\, Y => \I1.REG_74l323r\);
    
    \I2.SUB9l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_572_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l4r_net_1\);
    
    \I2.MIC_REG1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_306_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1l5r_net_1\);
    
    \I3.VDBi_57_ivl3r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855384__net_1\, B => 
        \I3.VDBi_43l3r_net_1\, C => 
        \I3.VDBi_57l3r_adt_net_145074_\, Y => \I3.VDBi_57l3r\);
    
    \I3.PIPEA1_311\ : MUX2L
      port map(A => \I3.PIPEA1l13r_net_1\, B => 
        \I3.PIPEA1_12l13r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__253\, Y => 
        \I3.PIPEA1_311_net_1\);
    
    \I2.PIPE8_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_557_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl29r_net_1\);
    
    \I2.PIPE3_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl6r_net_1\);
    
    \I2.DTE_cl_0_sqmuxa_2_adt_net_904_\ : OR3
      port map(A => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_N_20_i\, B
         => \I2.DTE_cl_0_sqmuxa_2_adt_net_20059__net_1\, C => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20061__net_1\, Y => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_904__net_1\);
    
    \I3.VDBoffa_44\ : OR3
      port map(A => \I3.VDBoffa_44_adt_net_164688_\, B => 
        \I3.VDBoffa_31l0r_adt_net_164649_\, C => 
        \I3.VDBoffa_31l0r_adt_net_164650_\, Y => 
        \I3.VDBoffa_44_net_1\);
    
    \I1.PAGECNT_0l9r_adt_net_835128_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854852__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\);
    
    \I2.UN1_REG80_I_1700\ : NOR3FTT
      port map(A => \I2.N_119\, B => REGl36r, C => REGl38r, Y => 
        \I2.N_3824_adt_net_90292_\);
    
    \I2.PIPE9_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_271_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl2r_net_1\);
    
    \I5.TEMPDATAl4r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_78_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl4r_net_1\);
    
    \I2.L2TYPE_4_il3r\ : OAI21FTF
      port map(A => \I2.L2TYPEl3r_net_1\, B => \I2.N_4465\, C => 
        \I2.N_4449_adt_net_68340_\, Y => \I2.N_4449\);
    
    \I2.LSRAM_INl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_386_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl2r_net_1\);
    
    \I1.NWRLUTi_0_sqmuxa_1_i_0\ : OAI21TTF
      port map(A => \I1.BYTECNTl8r_net_1\, B => \I1.N_435_1\, C
         => \I1.N_1192_adt_net_133761_\, Y => \I1.N_1192\);
    
    \I2.PIPE1_DT_42_0_IVL31R_1352\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\, B => 
        \I2.TDCDBSl31r_net_1\, C => 
        \I2.PIPE1_DT_42l31r_adt_net_45035_\, Y => 
        \I2.PIPE1_DT_42l31r_adt_net_45041_\);
    
    \I2.EVNT_NUM_n7\ : NOR2
      port map(A => EV_RES_c, B => \I2.EVNT_NUM_n7_tz_i\, Y => 
        \I2.EVNT_NUM_n7_net_1\);
    
    \I1.PAGECNT_n1_0_0_x2\ : XOR2FT
      port map(A => \I1.PAGECNTl1r_adt_net_834904_Rd1__net_1\, B
         => \I1.PAGECNTl0r_adt_net_833884_Rd1__net_1\, Y => 
        \I1.N_388_i_0_i\);
    
    TOKINB_pad : OB33PH
      port map(PAD => TOKINB, A => TOKINB_c);
    
    \I2.NWPIPE4\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE3_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE4_net_1\);
    
    \I2.OFFSET_37_5l0r\ : MUX2L
      port map(A => \REGl397r\, B => \REGl333r\, S => 
        \I2.PIPE7_DTL27R_85\, Y => \I2.N_667\);
    
    \I2.WPAGEL14R_2996\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_949_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEL14R_750\);
    
    \I2.CRC32_12_i_0_x2l10r\ : XOR2FT
      port map(A => \I2.CRC32l10r_net_1\, B => \I2.N_227_i_i\, Y
         => \I2.N_249_i_i_0\);
    
    \I3.STBMIC\ : DFFS
      port map(CLK => CLK_c, D => \I3.STBMIC_78_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => STBMIC_c);
    
    \I2.REG_1l38r\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n6_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGl38r);
    
    \I2.SUB9_1_ADD_18x18_fast_I111_un1_Y\ : NOR3FFT
      port map(A => \I2.N300\, B => \I2.N304\, C => \I2.N327\, Y
         => \I2.I111_un1_Y_adt_net_71419_\);
    
    \I2.LEAD_FLAG6_639\ : AO21
      port map(A => \I2.N_4533_adt_net_1164__net_1\, B => 
        \I2.N_4533_adt_net_64364_\, C => 
        \I2.LEAD_FLAG6_639_adt_net_64404_\, Y => 
        \I2.LEAD_FLAG6_639_net_1\);
    
    \I3.VDBI_57_0_IVL25R_2153\ : AND2
      port map(A => \I3.PIPEAl25r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l25r_adt_net_138707_\);
    
    \I2.DTE_21_1l10r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l10r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l10r_Rd1__net_1\);
    
    \I5.REG_1_28\ : MUX2H
      port map(A => \I5.SENS_ADDRl1r_net_1\, B => REGl445r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_28_net_1\);
    
    \I2.OFFSET_37_7l7r\ : MUX2L
      port map(A => \I2.N_682\, B => \I2.N_658\, S => 
        \I2.PIPE7_DTL25R_682\, Y => \I2.N_690\);
    
    \I2.DTE_21_1l9r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l9r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l9r_Rd1__net_1\);
    
    \I1.REG_74_0_IVL168R_2066\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l168r_adt_net_133407_\);
    
    \I2.OFFSET_37_19l6r\ : MUX2L
      port map(A => \REGl283r\, B => \REGl219r\, S => 
        \I2.PIPE7_DTL27R_87\, Y => \I2.N_785\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I39_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl18r\, B => 
        \I2.PIPE7_DTl18r_net_1\, Y => \I2.N285\);
    
    \I1.REG_1_236\ : MUX2H
      port map(A => \REGl335r\, B => \I1.REG_74l335r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y => 
        \I1.REG_1_236_net_1\);
    
    \I2.DTE_21_1_iv_0l12r\ : OR3
      port map(A => \I2.DTE_21_1l12r_adt_net_38283_\, B => 
        \I2.DTE_21_1l12r_adt_net_38297_\, C => 
        \I2.DTE_21_1l12r_adt_net_38298_\, Y => \I2.DTE_21_1l12r\);
    
    \I3.REG_1l99r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_280_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl99r\);
    
    \I2.RAMAD_4l14r\ : MUX2L
      port map(A => \I2.N_541\, B => 
        \I1.PAGECNTl6r_adt_net_854928__net_1\, S => LOAD_RES_1, Y
         => \I2.RAMAD_4l14r_net_1\);
    
    \I2.PIPE7_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl10r_net_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I23_Y_1643\ : OR2FT
      port map(A => \I2.N_3560_i_net_1\, B => \I2.N_3558_i_net_1\, 
        Y => \I2.N288_adt_net_68878_\);
    
    \I1.REG_74_0_IVL303R_1915\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l303r_adt_net_120610_\);
    
    \I2.FCNTl1r_1242\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_946_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.FCNTL1R_504\);
    
    \I2.RAMAD1_671\ : AO21FTT
      port map(A => 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_44987__net_1\, B => 
        \I2.RAMAD1l17r_net_1\, C => \I2.FIRST_TDC_1_sqmuxa_net_1\, 
        Y => \I2.RAMAD1_671_net_1\);
    
    \I2.STATE1l17r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3798\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1l17r_net_1\);
    
    \I2.BITCNT_n2_i_a5\ : NOR2
      port map(A => \I2.N_4327\, B => \I2.BITCNTl2r_net_1\, Y => 
        \I2.N_4335\);
    
    \I2.RAMAD1_12l15r\ : MUX2L
      port map(A => \I2.TDCDASl26r_net_1\, B => 
        \I2.TDCDBSl26r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855184__net_1\, Y => 
        \I2.RAMAD1_12l15r_net_1\);
    
    \I1.REG_1_188\ : MUX2H
      port map(A => \REGl287r\, B => \I1.REG_74l287r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\, Y => 
        \I1.REG_1_188_net_1\);
    
    \I1.PAGECNT_n3_0_0_o2\ : NAND2
      port map(A => \I1.PAGECNT_325_493\, B => \I1.N_300_Ra1_\, Y
         => \I1.N_305_Ra1_\);
    
    \I5.REG_1l420r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_33_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl420r);
    
    \I2.PIPE5_DT_6_0l9r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l9r\, B => 
        \I2.un27_pipe5_dt0l9r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1078\);
    
    \I2.BNCID_VECTrff_12\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_12_253_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_12\);
    
    \I1.N_145_adt_net_854768_\ : BFR
      port map(A => \I1.N_145\, Y => 
        \I1.N_145_adt_net_854768__net_1\);
    
    \I2.CRC32_806\ : MUX2L
      port map(A => \I2.CRC32l11r_net_1\, B => \I2.N_3928\, S => 
        \I2.N_2826_1_ADT_NET_794__332\, Y => \I2.CRC32_806_net_1\);
    
    \I2.DT_SRAMl10r\ : MUX2L
      port map(A => \I2.N_878\, B => \I2.PIPE2_DTl10r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.DT_SRAMl10r_net_1\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__2833\ : NAND3FFT
      port map(A => \I2.ENDF_838\, B => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__184\, C => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_60\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__181\);
    
    \I5.TEMP_ACK\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMP_ACK_73_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMP_ACK_net_1\);
    
    \I2.ADOl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl2r);
    
    \I1.SBYTE_64\ : MUX2L
      port map(A => \FBOUTl6r\, B => \I1.N_206\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_64_net_1\);
    
    \I3.REGMAPl16r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un64_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPl16r_net_1\);
    
    \I5.un1_tick_5_i\ : NAND2FT
      port map(A => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\, B => 
        \I5.N_479\, Y => \I5.N_461\);
    
    \I3.VDBi_43l1r\ : MUX2L
      port map(A => REGl407r, B => \I3.VDBi_40l1r_net_1\, S => 
        \I3.REGMAPl55r_net_1\, Y => \I3.VDBi_43l1r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2598\ : OR3
      port map(A => \I3.VDBoffa_31l2r_adt_net_164265_\, B => 
        \I3.VDBoffa_31l2r_adt_net_164259_\, C => 
        \I3.VDBoffa_31l2r_adt_net_164260_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164269_\);
    
    \I1.N_341_RD1__2970\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_341_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_341_RD1__487\);
    
    \HWRES_3_ADT_NET_738__2744\ : NAND2
      port map(A => NPWON_c, B => SYSRESB_c, Y => 
        \HWRES_3_ADT_NET_738__17\);
    
    \I1.PAGECNTLDE_0_1760\ : OAI21TTF
      port map(A => \I1.N_591_1\, B => \I1.N_328_I_0_212\, C => 
        \I1.N_370\, Y => \I1.PAGECNTe_adt_net_106660_\);
    
    \I1.REG_74_0_IVL214R_2020\ : AND2
      port map(A => \FBOUTl1r\, B => \I1.REG_7_sqmuxa\, Y => 
        \I1.REG_74l214r_adt_net_129292_\);
    
    \I3.UN15_ANYCYC_2299\ : NOR3FFT
      port map(A => \I3.MBLTCYC_844\, B => \I3.PIPEBl30r_net_1\, 
        C => \I3.PIPEBl29r_net_1\, Y => 
        \I3.un15_anycyc_adt_net_147620_\);
    
    \I2.ENDF_712\ : MUX2L
      port map(A => \I2.ENDF_net_1\, B => \I2.un1_STATE2_9\, S
         => \I2.un1_STATE2_7\, Y => \I2.ENDF_712_net_1\);
    
    \I2.MIC_ERR_REGS_364\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl36r_net_1\, B => 
        \I2.MIC_ERR_REGSl35r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_364_net_1\);
    
    \I2.TDCDRYAS\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDRYA_c, Q => 
        \I2.TDCDRYAS_net_1\);
    
    \I1.BYTECNT_N2_I_1778\ : XOR2
      port map(A => \I1.BYTECNTl2r_adt_net_855020__net_1\, B => 
        \I1.N_323_adt_net_108906_\, Y => 
        \I1.N_174_adt_net_108976_\);
    
    \I2.un1_STATE1_38_0_a2_1_0_a3\ : OR2
      port map(A => \I2.STATE1l18r_net_1\, B => 
        \I2.STATE1_i_0_il15r\, Y => \I2.N_3358\);
    
    \I1.REG_74_0_IVL353R_1860\ : NOR2FT
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_24_sqmuxa_adt_net_854776__net_1\, Y => 
        \I1.REG_74l353r_adt_net_115859_\);
    
    \I3.TCNT3_379\ : XOR2
      port map(A => \I3.TCNT3_i_0_il0r_net_1\, B => \TICKl1r\, Y
         => \I3.TCNT3_379_net_1\);
    
    \I3.VDBm_0l21r\ : MUX2L
      port map(A => \I3.PIPEAl21r_net_1\, B => 
        \I3.PIPEBl21r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_163\);
    
    \I1.REG_17_sqmuxa_0_a2_0_a3_0_a2_844\ : NAND2
      port map(A => \I1.N_590_231\, B => \I1.PAGECNTL9R_246\, Y
         => \I1.N_260_222\);
    
    \I2.DTE_21_1_IV_0L6R_1322\ : AND2
      port map(A => \I2.DTE_1l6r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\, Y => 
        \I2.DTE_21_1l6r_adt_net_38973_\);
    
    \I2.PIPE8_DT_21l12r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl12r\, B => \I2.N_578\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l12r_net_1\);
    
    \I2.CRC32_12_i_x2l0r\ : XOR2FT
      port map(A => \I2.CRC32l0r_net_1\, B => \I2.N_3954_i_i\, Y
         => \I2.N_4027_i_0\);
    
    \I3.VDBi_40_0_i_m2l5r\ : MUX2L
      port map(A => REGl423r, B => REGl439r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_137\);
    
    \I2.CHA_DATA8_2_i_o2\ : NOR2
      port map(A => \I2.N_4401\, B => \I2.PIPE7_DTl29r_net_1\, Y
         => \I2.N_4403\);
    
    REGl401r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_302_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl401r\);
    
    \I1.N_310_RD1__2892\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_310_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_310_RD1__335\);
    
    FID_padl18r : OB33PH
      port map(PAD => FID(18), A => FID_cl18r);
    
    \I3.TCNT1_n5\ : XOR2FT
      port map(A => \I3.TCNT1l5r_net_1\, B => \I3.TCNT1_c4_net_1\, 
        Y => \I3.TCNT1_n5_net_1\);
    
    \I2.OFFSET_37_24l3r\ : MUX2L
      port map(A => \I2.N_814\, B => \I2.N_806\, S => 
        \I2.PIPE7_DTL26R_358\, Y => \I2.N_822\);
    
    \I2.WMIC\ : DFFB
      port map(CLK => MWOK_c, D => \GND\, CLR => 
        \HWRES_3_adt_net_738__net_1\, SET => PULSEl4r, Q => 
        WMIC_c);
    
    DTE_padl3r : IOB33PH
      port map(PAD => DTE(3), A => \I2.DTE_1l3r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl3r);
    
    \I2.REG_1_c11_i_o2\ : AND3
      port map(A => REG_i_0_il42r, B => REGl43r, C => \I2.N_3853\, 
        Y => \I2.N_3856\);
    
    TDCDA_padl20r : IB33
      port map(PAD => TDCDA(20), Y => TDCDA_cl20r);
    
    \I2.PIPE1_DT_30l13r\ : MUX2L
      port map(A => \I2.TDCDBSl13r_net_1\, B => 
        \I2.TDCDBSl11r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, Y
         => \I2.PIPE1_DT_30l13r_net_1\);
    
    \I2.END_EVNT4\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT3_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT4_net_1\);
    
    \I2.SUB9l9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_577_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9_i_0_il9r\);
    
    \I1.N_50_0_ADT_NET_109751__2863\ : NOR3FFT
      port map(A => \I1.N_232_1_296\, B => 
        \I1.N_50_0_adt_net_109760__net_1\, C => \I1.N_435_1_285\, 
        Y => \I1.N_50_0_ADT_NET_109751__258\);
    
    \I2.N_4528_adt_net_1129_\ : AO21
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_219\, C
         => LEAD_FLAGl7r, Y => \I2.N_4528_adt_net_1129__net_1\);
    
    \I3.PIPEAl19r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_250_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl19r_net_1\);
    
    \I1.REG_30_sqmuxa_adt_net_854372_\ : BFR
      port map(A => \I1.REG_30_sqmuxa_adt_net_854376__net_1\, Y
         => \I1.REG_30_sqmuxa_adt_net_854372__net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I141_Y_0_o4\ : AOI21
      port map(A => \I2.N_13_0\, B => \I2.N525\, C => \I2.N_16\, 
        Y => \I2.N522\);
    
    \I2.PIPE4_DTL4R_2960\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL4R_477\);
    
    \I2.PIPE5_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_687_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl11r_net_1\);
    
    \I2.MIC_ERR_REGSl43r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_372_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl43r_net_1\);
    
    \I1.REG_1_238\ : MUX2H
      port map(A => \REGl337r\, B => \I1.REG_74l337r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855500__net_1\, Y => 
        \I1.REG_1_238_net_1\);
    
    \I3.VDBml4r\ : MUX2L
      port map(A => \I3.VDBil4r_net_1\, B => \I3.N_146\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml4r_net_1\);
    
    \I3.STATE1_illegal\ : OR2
      port map(A => \I3.N_1193_ip_adt_net_136557_\, B => 
        \I3.N_1193_ip_adt_net_136558_\, Y => \I3.N_1193_ip\);
    
    \I2.OFFSET_37_13l4r\ : MUX2L
      port map(A => \I2.N_727\, B => \I2.N_711\, S => 
        \I2.PIPE7_DTL25R_684\, Y => \I2.N_735\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854188_\ : BFR
      port map(A => \I2.N_4667_1_ADT_NET_1046__35\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854188__net_1\);
    
    REGl220r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_121_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl220r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I213_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl17r\, B => 
        \I2.PIPE7_DTl17r_net_1\, Y => 
        \I2.SUB_21x21_fast_I213_Y_0\);
    
    \I2.REG_1_c1_i\ : OAI21TTF
      port map(A => \I2.un8_evread_1_adt_net_855780__net_1\, B
         => \I2.N_3844\, C => \I2.N_3830_adt_net_101622_\, Y => 
        \I2.N_3830\);
    
    \I3.VDBi_57_iv_0_0_a2_13l2r\ : NOR2
      port map(A => \I3.N_1904\, B => 
        \I3.N_57_i_0_0_adt_net_854688__net_1\, Y => \I3.N_2048\);
    
    \I2.SUB9_1_ADD_18x18_fast_I157_Y\ : XOR2FT
      port map(A => \I2.SUB8l20r_net_1\, B => \I2.N434\, Y => 
        \I2.SUB9_1l20r\);
    
    \I2.RAMAD1l3r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_657_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l3r_net_1\);
    
    \I2.PIPE5_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_682_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl6r_net_1\);
    
    \I3.PIPEB_103\ : AO21
      port map(A => DPR_cl24r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855272__net_1\, 
        C => \I3.PIPEB_103_adt_net_159705_\, Y => 
        \I3.PIPEB_103_net_1\);
    
    \I2.PIPE5_DT_688\ : MUX2L
      port map(A => \I2.PIPE5_DTl12r_net_1\, B => 
        \I2.PIPE5_DT_6l12r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_688_net_1\);
    
    \I2.LEAD_FLAG6_7_i_0_a2_1l5r\ : NOR2FT
      port map(A => \I2.PIPE5_DTl30r_net_1\, B => 
        \I2.PIPE5_DTl22r_net_1\, Y => \I2.N_483\);
    
    \I1.NWRLUTi_0_sqmuxa_1_i_0_o2\ : NOR2
      port map(A => \I1.sstatel8r_net_1\, B => 
        \I1.sstatel5r_net_1\, Y => \I1.N_380\);
    
    \I3.PIPEA_231\ : MUX2L
      port map(A => \I3.PIPEAl0r_net_1\, B => 
        \I3.PIPEA_8l0r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854680__net_1\, Y
         => \I3.PIPEA_231_net_1\);
    
    TDCDB_padl1r : IB33
      port map(PAD => TDCDB(1), Y => TDCDB_cl1r);
    
    \I2.PIPE2_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl17r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl17r_net_1\);
    
    \I2.LEAD_FLAG6_642\ : AO21
      port map(A => \I2.N_4530_adt_net_1143__net_1\, B => 
        \I2.N_4530_adt_net_64028_\, C => 
        \I2.LEAD_FLAG6_642_adt_net_64068_\, Y => 
        \I2.LEAD_FLAG6_642_net_1\);
    
    \I2.L2TYPE_597\ : MUX2L
      port map(A => \I2.L2TYPEl8r_net_1\, B => \I2.N_4444\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_597_net_1\);
    
    \I3.REG_1_263_e\ : AND3
      port map(A => \I3.REGMAPl12r_net_1\, B => 
        \I3.STATE1_IPL8R_10\, C => \I3.N_127\, Y => \I3.N_2277_i\);
    
    \I2.un1_sram_evnt12_i\ : OR2
      port map(A => \I2.N_3823_adt_net_90689_\, B => \I2.N_132\, 
        Y => \I2.N_3823\);
    
    \I1.sstate_tr28_0_a2_0_a4\ : NOR2FT
      port map(A => \I1.sstatel2r_net_1\, B => 
        \PULSE_0l0r_adt_net_834380_Rd1__net_1\, Y => 
        \I1.sstate_nsl9r\);
    
    \I2.OFFSET_37_10l5r\ : MUX2L
      port map(A => \I2.N_704\, B => \I2.N_696\, S => 
        \I2.PIPE7_DTL26R_352\, Y => \I2.N_712\);
    
    \I2.N_4283_i_0_adt_net_854972_\ : BFR
      port map(A => \I2.N_4283_I_0_235\, Y => 
        \I2.N_4283_i_0_adt_net_854972__net_1\);
    
    \I5.N_155_0_adt_net_983__adt_net_855864_\ : BFR
      port map(A => \I5.N_155_0_adt_net_983__net_1\, Y => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\);
    
    \I3.VDBi_57l7r_adt_net_143035_\ : AO21
      port map(A => \I3.REGl140r\, B => \I3.N_2046\, C => 
        \I3.VDBi_57l7r_adt_net_143034__net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_143035__net_1\);
    
    \I2.STATE1l2r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1l3r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1l2r_net_1\);
    
    \I4.un1_lead_flag_1_7_0\ : MUX2L
      port map(A => \I4.N_6\, B => \I4.N_3\, S => 
        \I4.bcntl0r_net_1\, Y => \I4.un1_lead_flag_1\);
    
    \I2.PIPE10_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_630_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl25r_net_1\);
    
    \I3.REG_1_ml76r\ : AND2
      port map(A => REGl76r, B => 
        \I3.REGMAPl9r_adt_net_854304__net_1\, Y => 
        \I3.VDBi_20l28r\);
    
    \I2.MIC_ERR_REGSl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_333_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl4r_net_1\);
    
    \I1.REG_74_0_iv_0l369r\ : AO21
      port map(A => \REGl369r\, B => \I1.N_660\, C => 
        \I1.REG_74l369r_adt_net_113568_\, Y => \I1.REG_74l369r\);
    
    \I2.PIPE4_DTl5r_adt_net_854412_\ : BFR
      port map(A => \I2.PIPE4_DTl5r_adt_net_854416__net_1\, Y => 
        \I2.PIPE4_DTl5r_adt_net_854412__net_1\);
    
    \I2.STATE1l18r_1769\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_o2_0l0r_net_1\, SET => CLEAR_STAT_i_0, Q
         => \I2.STATE1L18R_875\);
    
    GA_padl1r : IB33
      port map(PAD => GA(1), Y => GA_cl1r);
    
    \I2.FIDl26r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_442\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl26r);
    
    \I3.VDBI_57_0_IV_0_0L13R_2193\ : AO21FTT
      port map(A => \I3.N_354_0_adt_net_855368__net_1\, B => 
        \I3.N_2276\, C => \I3.VDBi_57l13r_adt_net_140499_\, Y => 
        \I3.VDBi_57l13r_adt_net_140454_\);
    
    \I2.L2TYPEl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_602_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_i_0_il13r\);
    
    \I2.PIPE2_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl13r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl13r_net_1\);
    
    \I2.PIPE4_DTl11r_1147_1735\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL11R_842\);
    
    \I2.PIPE8_DT_21l15r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl15r\, B => 
        \I2.PIPE8_DT_16l15r_net_1\, S => \I2.NWPIPE7_net_1\, Y
         => \I2.PIPE8_DT_21l15r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I144_Y_0\ : XOR2
      port map(A => \I2.N_3541_i_i\, B => \I2.G_1_1\, Y => 
        \I2.ADD_18x18_fast_I144_Y_0\);
    
    \I2.resyn_0_I2_BITCNT_939\ : MUX2H
      port map(A => \I2.BITCNTl1r_net_1\, B => \I2.N_4322\, S => 
        \I2.BITCNTe\, Y => \I2.BITCNT_939\);
    
    \I2.PIPE8_DT_21l22r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl22r\, B => 
        \I2.PIPE7_DTl22r_net_1\, S => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l22r_net_1\);
    
    \I2.N_3279_0_adt_net_855228_\ : BFR
      port map(A => \I2.N_3279_0_adt_net_855236__net_1\, Y => 
        \I2.N_3279_0_adt_net_855228__net_1\);
    
    \I3.TCNT_N2_0_0_2137\ : XOR2FT
      port map(A => \I3.N_1911\, B => \I3.TCNTl2r_net_1\, Y => 
        \I3.TCNT_n2_adt_net_137234_\);
    
    \I2.un28_sram_empty_1_0\ : MUX2L
      port map(A => \I2.L2TYPEL8R_650\, B => \I2.L2TYPEL0R_649\, 
        S => \I2.RPAGEL15R_515\, Y => \I2.N_620\);
    
    \I2.FIFO_END_EVNT\ : DFFC
      port map(CLK => CLK_c, D => \I2.FIFO_END_EVNT_489_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.FIFO_END_EVNT_net_1\);
    
    \I2.DT_SRAM_0l5r\ : MUX2L
      port map(A => \I2.PIPE10_DTl5r_net_1\, B => 
        \I2.PIPE5_DTl5r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854228__net_1\, Y => 
        \I2.N_873\);
    
    \I2.PIPE5_DT_6_0l11r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l11r\, B => 
        \I2.un27_pipe5_dt0l11r\, S => 
        \I2.dataout_0_adt_net_855804__net_1\, Y => \I2.N_1080\);
    
    \I3.PIPEA1l25r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_323_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l25r_net_1\);
    
    \I2.RAMAD_4_0l0r\ : MUX2H
      port map(A => \I2.RAMAD1l0r_net_1\, B => RAMAD_VMEl0r, S
         => \REG_i_il5r_adt_net_855560__net_1\, Y => \I2.N_527\);
    
    \I1.BYTECNT_n5_i_0_o2_0\ : AND2
      port map(A => \I1.BYTECNTl3r_net_1\, B => \I1.N_323\, Y => 
        \I1.N_327\);
    
    \I3.VDBoffa_31_iv_0l1r\ : AND2
      port map(A => \REGl206r\, B => 
        \I3.REGMAPl23r_adt_net_855016__net_1\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164404_\);
    
    \I2.PIPE9_DT_278\ : MUX2L
      port map(A => \I2.PIPE9_DTl9r_net_1\, B => 
        \I2.PIPE8_DTl9r_net_1\, S => \I2.NWPIPE8_i_0_i_0_0\, Y
         => \I2.PIPE9_DT_278_net_1\);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_1_sqmuxa_0_a4_i_o2_47_tz\ : 
        AO21FTT
      port map(A => LEAD_FLAGl7r, B => \I2.PIPE4_DTl21r_net_1\, C
         => \I2.N_2329_tz_adt_net_16479_\, Y => \I2.N_2329_tz\);
    
    \I2.RAMAD1_12l7r\ : MUX2L
      port map(A => \I2.TDCDASl5r_net_1\, B => 
        \I2.TDCDBSl5r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855180__net_1\, Y => 
        \I2.RAMAD1_12l7r_net_1\);
    
    \I3.REG2l6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG2_147_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l6r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I146_Y_0\ : XOR2
      port map(A => \I2.N_3545_i_i\, B => \I2.G_1\, Y => 
        \I2.ADD_18x18_fast_I146_Y_0\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I120_Y_0_1587\ : AO21FTT
      port map(A => \I2.N_72_0\, B => \I2.N_93_0\, C => 
        \I2.N531_0_adt_net_60100_\, Y => 
        \I2.N531_0_adt_net_60059_\);
    
    \I3.un41_reg_ads_0_a2_3_a3\ : NOR2
      port map(A => \I3.un41_reg_ads_0_a2_3_a3_0\, B => 
        \I3.un41_reg_ads_2\, Y => 
        \I3.un41_reg_ads_0_a2_3_a3_net_1\);
    
    VAD_padl30r : IOB33PH
      port map(PAD => VAD(30), A => \I3.VADml30r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl30r);
    
    TDCDB_padl19r : IB33
      port map(PAD => TDCDB(19), Y => TDCDB_cl19r);
    
    \I2.DTOSl21r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl21r, Q => 
        \I2.DTOSl21r_net_1\);
    
    \I1.PAGECNT_326_824\ : MUX2H
      port map(A => \I1.PAGECNTl1r_adt_net_834904_Rd1__net_1\, B
         => \I1.PAGECNT_n1\, S => 
        \I1.PAGECNTe_adt_net_854900__net_1\, Y => 
        \I1.PAGECNT_326_202\);
    
    \I2.OFFSET_37_29l6r\ : MUX2L
      port map(A => \I2.N_857\, B => \I2.N_745\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l6r\);
    
    \I2.RAMAD_4_0l15r\ : MUX2H
      port map(A => \I2.RAMAD1l15r_net_1\, B => RAMAD_VMEl15r, S
         => \REG_i_il5r_adt_net_855552__net_1\, Y => \I2.N_542\);
    
    \I5.SENS_ADDR_1_sqmuxa_1_0\ : NAND2
      port map(A => REGL117R_390, B => TICKL0R_2, Y => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_net_1\);
    
    \I3.PULSE_46_0_iv_i_i_o2_0l3r\ : NOR2
      port map(A => \I3.STATE1_IPL9R_427\, B => 
        \I3.STATE1_IPL8R_426\, Y => \I3.N_291\);
    
    \I3.PIPEB_82_2341\ : NOR2FT
      port map(A => \I3.PIPEBl3r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_82_adt_net_160587_\);
    
    \I2.DT_TEMP_7l30r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854232__net_1\, B => 
        \I2.DT_SRAMl30r_adt_net_854200__net_1\, Y => 
        \I2.DT_TEMP_7l30r_net_1\);
    
    \I1.BYTECNTlde_i_a2_i\ : AO21
      port map(A => \I1.N_628\, B => 
        \I1.sstate_ns_i_0_a4_0_1l0r_adt_net_107171_\, C => 
        \I1.N_223_226\, Y => \I1.N_1383\);
    
    \I2.N_128_adt_net_54291__adt_net_854408_\ : BFR
      port map(A => \I2.N_128_adt_net_54291_\, Y => 
        \I2.N_128_adt_net_54291__adt_net_854408__net_1\);
    
    REGl244r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_145_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl244r\);
    
    \I3.REG_1l139r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_187_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl139r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I144_Y\ : XOR2FT
      port map(A => \I2.N344\, B => \I2.ADD_18x18_fast_I144_Y_0\, 
        Y => \I2.SUB9_1l7r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I199_Y\ : XOR2FT
      port map(A => \I2.N510_adt_net_220925_\, B => 
        \I2.SUB_21x21_fast_I199_Y_0\, Y => \I2.SUB8_2l3r\);
    
    \I2.un1_DTO_cl_1_sqmuxa_2_0_o2_1_0_x2\ : XOR2FT
      port map(A => NOESRAME_C_240, B => 
        \I2.WOFFSETl0r_adt_net_854648__net_1\, Y => \I2.N_176_i\);
    
    \I2.CRC32_816\ : MUX2L
      port map(A => \I2.CRC32l21r_net_1\, B => \I2.N_3938\, S => 
        \I2.N_2826_1_ADT_NET_794__330\, Y => \I2.CRC32_816_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I34_Y\ : OA21TTF
      port map(A => \I2.SUB8l11r_net_1\, B => \I2.N_3547_i_i\, C
         => \I2.SUB8l12r_net_1\, Y => \I2.N299\);
    
    \I2.EVNT_NUM_959\ : MUX2L
      port map(A => \I2.EVNT_NUMl4r_net_1\, B => 
        \I2.EVNT_NUM_n4_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_959_net_1\);
    
    \I2.PIPE7_DTL27R_2781\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_74\);
    
    \I2.PIPE5_DT_6_sl19r\ : OR2
      port map(A => \I2.dataout_0_adt_net_855800__net_1\, B => 
        \I2.N_4547_1_adt_net_1209__net_1\, Y => 
        \I2.PIPE5_DT_6_sl19r_net_1\);
    
    \I2.L2TYPE_4_i_o2l11r\ : NOR2
      port map(A => \I2.N_4454\, B => \I2.N_4459\, Y => 
        \I2.N_4467\);
    
    \I3.REG_1l63r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_164_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl63r);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854672_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854672__net_1\);
    
    \I2.OFFSETl5r_1567\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_565_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL5R_674\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I29_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl8r\, B => \I2.PIPE7_DTL8R_697\, 
        Y => \I2.N255_0\);
    
    \I2.TDCDBSl16r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl16r, Q => 
        \I2.TDCDBSl16r_net_1\);
    
    \I3.PIPEA_8l4r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854484__net_1\, B => 
        \I3.N_213\, Y => \I3.PIPEA_8l4r_net_1\);
    
    \I3.VDBi_362\ : MUX2L
      port map(A => \I3.VDBil22r_net_1\, B => \I3.VDBi_57l22r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_362_net_1\);
    
    \I3.REG_1l406r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_213_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl406r);
    
    \I3.VADm_0_a3l26r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl26r_net_1\, Y => \I3.VADml26r\);
    
    \I1.REG_74_12_220_M9_I_1998\ : OAI21TTF
      port map(A => \I1.REG_74_12_220_m9_i_a6_0\, B => 
        \I1.REG_74_12_220_N_13\, C => 
        \I1.N_1169_adt_net_854824__net_1\, Y => 
        \I1.REG_74_12_220_m9_i_adt_net_127882_\);
    
    \I5.SDAOUT_12_IV_0_O4_0_906\ : NOR2
      port map(A => \I5.N_64\, B => \I5.COMMANDl1r_net_1\, Y => 
        \I5.N_75_adt_net_8973_\);
    
    \I3.VDBoff_4_i_il3r\ : MUX2L
      port map(A => \I3.VDBoffbl3r_net_1\, B => 
        \I3.VDBoffal3r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_2067\);
    
    \I1.N_308_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_308_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_308_Rd1__net_1\);
    
    \I2.TOKOUTBS_3_i\ : MUX2H
      port map(A => TOKOUTB_BP_c, B => TOKOUTB_c, S => 
        \I2.N_4431\, Y => \I2.TOKOUTBS_3_i_net_1\);
    
    \I2.PIPE6_DT_464\ : MUX2H
      port map(A => \I2.PIPE5_DTl10r_net_1\, B => 
        \I2.PIPE6_DTl10r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_464_net_1\);
    
    \I2.PIPE5_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_695_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl19r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I57_Y\ : NAND2
      port map(A => \I2.N267_0_868\, B => \I2.N264_0_866\, Y => 
        \I2.N307_2\);
    
    \I2.DTE_21_1_0_IV_0_0L29R_1231\ : AND2FT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855192__net_1\, 
        B => \I2.DT_TEMPl29r_net_1\, Y => 
        \I2.DTE_21_1l29r_adt_net_36645_\);
    
    \I2.SRAM_FULL_488\ : MUX2H
      port map(A => \I2.SRAM_FULL_net_1\, B => 
        \I2.START_GIRO_net_1\, S => \I2.N_3823\, Y => 
        \I2.SRAM_FULL_488_net_1\);
    
    \I2.ADE_4l2r\ : MUX2H
      port map(A => \I2.WOFFSETl3r_adt_net_854988__net_1\, B => 
        \I2.ROFFSETl3r_net_1\, S => NOESRAME_c, Y => 
        \I2.ADE_4l2r_net_1\);
    
    \I2.TDCDBSl18r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl18r, Q => 
        \I2.TDCDBSl18r_net_1\);
    
    N_1_I3_TCNT2_c1 : AND2
      port map(A => \I3.TCNT2_i_0_il0r_net_1\, B => 
        \I3.TCNT2l1r_net_1\, Y => \I3.TCNT2_c1\);
    
    \I2.REG_1_n11\ : XOR2FT
      port map(A => \I2.N_3839_i_0\, B => \I2.REG_1_n11_0_net_1\, 
        Y => \I2.REG_1_n11_net_1\);
    
    \I1.N_113_ADT_NET_3714__2865\ : OR2
      port map(A => \I1.N_41_9_adt_net_854784__net_1\, B => 
        \I1.N_113_adt_net_126306__net_1\, Y => 
        \I1.N_113_ADT_NET_3714__270\);
    
    \I3.REG_1l148r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_196_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl148r\);
    
    \I3.VDBOFFB_30_IV_0L3R_2435\ : OR2
      port map(A => \I3.VDBoffb_30l3r_adt_net_162551_\, B => 
        \I3.VDBoffb_30l3r_adt_net_162552_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162557_\);
    
    \I2.LSRAM_INl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_391_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl7r_net_1\);
    
    \I2.RESYN_0_I2_UN1_TRGCNT14_I_939\ : NOR2
      port map(A => \I2.TRGCNT_i_0_il3r\, B => 
        \I2.TRGCNTl2r_net_1\, Y => \I2.N_3760_adt_net_15913_\);
    
    \I2.L2ARR_c1_i_o2\ : NAND2
      port map(A => \I2.L2ARRl1r_net_1\, B => \I2.L2ARRl0r_net_1\, 
        Y => \I2.N_4454\);
    
    \I2.PIPE8_DT_21l25r\ : MUX2H
      port map(A => \I2.PIPE7_DTl25r_net_1\, B => 
        \I2.LSRAM_OUTl25r\, S => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l25r_net_1\);
    
    \I2.REG_1_n5_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855784__net_1\, B
         => REGl37r, Y => \I2.REG_1_n5_0_net_1\);
    
    \I2.FID_7_0_IVL16R_960\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl64r, C => 
        \I2.FID_7l16r_adt_net_17799_\, Y => 
        \I2.FID_7l16r_adt_net_17807_\);
    
    \I2.DTE_1_864\ : MUX2L
      port map(A => \I2.DTE_1l26r_Rd1__net_1\, B => 
        \I2.DTE_21_1l26r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\, Y => 
        \I2.DTE_1l26r\);
    
    \I1.REG_1_179\ : MUX2H
      port map(A => \REGl278r\, B => \I1.REG_74l278r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\, Y => 
        \I1.REG_1_179_net_1\);
    
    \I2.DTO_16_1_IV_0_0L18R_1127\ : NOR3
      port map(A => \I2.DTO_16_1_iv_0_a2_4_18_N_12_i\, B => 
        \I2.DTO_16_1_iv_0_a2_4_18_N_14_i\, C => 
        \I2.DTO_16_1_iv_0_a2_4_18_m7_0_0_i\, Y => 
        \I2.DTO_16_1l18r_adt_net_31339_\);
    
    \I1.REG_74_0_IVL213R_2021\ : AND2
      port map(A => \FBOUTl0r\, B => \I1.REG_7_sqmuxa\, Y => 
        \I1.REG_74l213r_adt_net_129378_\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2395\ : AO21
      port map(A => \REGl330r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l5r_adt_net_162140_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162172_\);
    
    \I2.un2_evnt_word_I_8\ : AND2
      port map(A => \I2.WOFFSETl0r_adt_net_854636__net_1\, B => 
        \I2.WOFFSETl1r_adt_net_854992__net_1\, Y => \I2.N_50\);
    
    \I2.PIPE1_DT_12l0r\ : MUX2H
      port map(A => \I2.TDCDASl19r_net_1\, B => 
        \I2.TDCDASl0r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855100__net_1\, Y
         => \I2.PIPE1_DT_12l0r_net_1\);
    
    \I2.PIPE8_DT_21l14r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl14r_adt_net_854944__net_1\, B
         => \I2.PIPE8_DT_16l14r_net_1\, S => \I2.NWPIPE7_net_1\, 
        Y => \I2.PIPE8_DT_21l14r_net_1\);
    
    \I2.DTE_1_842\ : MUX2L
      port map(A => \I2.DTE_1l2r_net_1\, B => 
        \I2.DTE_21_1_iv_i_0l2r\, S => \I2.N_2868_1\, Y => 
        \I2.DTE_1_842_net_1\);
    
    \I5.sstate1l12r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el1r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l12r_net_1\);
    
    \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_N_8_RD1__2968\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_N_8_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_N_8_RD1__485\);
    
    \I3.PIPEAl26r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_257_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl26r_net_1\);
    
    \I3.N_264_0_ADT_NET_1653_RD1__2819\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.N_264_0_adt_net_1653_Ra1__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.N_264_0_ADT_NET_1653_RD1__147\);
    
    \I3.REG_1l58r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_159_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl58r);
    
    DTO_padl27r : IOB33PH
      port map(PAD => DTO(27), A => \I2.DTO_1l27r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl27r);
    
    \I2.RMIC\ : DFFLB
      port map(CLK => MROK_c, D => \GND\, CLR => \I2.un8_hwres_i\, 
        SET => PULSEl5r, Q => RMIC_c);
    
    \I2.DTE_21_1_0_IVL31R_1228\ : AO21
      port map(A => \I2.STATE2L3R_440\, B => \I2.DTO_9l31r\, C
         => \I2.DTE_21_1l31r_adt_net_36416_\, Y => 
        \I2.DTE_21_1l31r_adt_net_36417_\);
    
    \I5.COMMAND_4l13r\ : AND2FT
      port map(A => REGl7r, B => REGl114r, Y => 
        \I5.COMMAND_4l13r_net_1\);
    
    \I1.REG_74_0_iv_0_0l254r\ : AO21
      port map(A => \REGl254r\, B => \I1.N_658\, C => 
        \I1.REG_74l254r_adt_net_125314_\, Y => \I1.REG_74l254r\);
    
    \I2.DTO_16_1_IVL10R_1170\ : AND2
      port map(A => \I2.N_4671_adt_net_854596__net_1\, B => 
        \I2.DT_TEMPl10r_net_1\, Y => 
        \I2.DTO_16_1l10r_adt_net_33056_\);
    
    \I1.REG_74_0_IV_0_0L255R_1970\ : AND2
      port map(A => \FBOUTl2r\, B => \I1.N_596\, Y => 
        \I1.REG_74l255r_adt_net_125228_\);
    
    \I2.CHAINB_ERRF1\ : DFFC
      port map(CLK => CLK_c, D => \I2.CHAINB_ERRF1_493_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.CHAINB_ERRF1_net_1\);
    
    \I2.DTE_21_1_IV_0L16R_1269\ : AND2
      port map(A => \I2.DTE_1l16r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1l16r_adt_net_37823_\);
    
    \I2.OFFSET_37_23l4r\ : MUX2L
      port map(A => \REGl273r\, B => \REGl209r\, S => 
        \I2.PIPE7_DTL27R_89\, Y => \I2.N_815\);
    
    \I2.PIPE9_DT_277\ : MUX2L
      port map(A => \I2.PIPE9_DTl8r_net_1\, B => 
        \I2.PIPE8_DTl8r_net_1\, S => \I2.NWPIPE8_i_0_i_0_0\, Y
         => \I2.PIPE9_DT_277_net_1\);
    
    \I1.REG_74_0_ivl387r\ : AO21
      port map(A => \REGl387r\, B => \I1.N_257\, C => 
        \I1.REG_74l387r_adt_net_111405_\, Y => \I1.REG_74l387r\);
    
    \I3.VDBOFFA_31_IV_0L1R_2606\ : AND2
      port map(A => \REGl278r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        Y => \I3.VDBoffa_31l1r_adt_net_164428_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I138_Y_0\ : AND2FT
      port map(A => \I2.N_100_0\, B => 
        \I2.N513_i_0_adt_net_58712_\, Y => \I2.N513_i_0\);
    
    \I2.L2ARRl2r_1497\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_942_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRL2R_604\);
    
    \I2.PIPE10_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_628_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl23r_net_1\);
    
    \I2.ROFFSET_226\ : NAND2FT
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855704__net_1\, B => 
        \I2.ROFFSETl1r_net_1\, Y => \I2.N_1357\);
    
    \I5.REG_1_44\ : MUX2L
      port map(A => \I5.REG_12l431r_net_1\, B => REGl431r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_44_net_1\);
    
    \I3.VDBI_57_0_IVL29R_2144\ : AO21
      port map(A => \I3.VDBil29r_net_1\, B => 
        \I3.N_1910_0_adt_net_854340__net_1\, C => 
        \I3.VDBi_57l29r_adt_net_138169_\, Y => 
        \I3.VDBi_57l29r_adt_net_138175_\);
    
    \I2.STATE3_NS_A7L9R_1042\ : AND2
      port map(A => \I2.STATE3l5r_net_1\, B => 
        \I3.N_203_adt_net_854976__net_1\, Y => 
        \I2.N_12254_i_adt_net_24491_\);
    
    \I3.VDBI_57_IV_0_0L2R_2261\ : NOR2FT
      port map(A => \FBOUTl2r\, B => \I3.N_2047\, Y => 
        \I3.VDBi_57l2r_adt_net_145368_\);
    
    \I2.SUB8l6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_509_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l6r_net_1\);
    
    \I2.RAMAD_4_0l9r\ : MUX2H
      port map(A => \I2.RAMAD1l9r_net_1\, B => RAMAD_VMEl9r, S
         => \REG_i_il5r_adt_net_855556__net_1\, Y => \I2.N_536\);
    
    \I2.STATE3l8r\ : DFFS
      port map(CLK => CLK_c, D => \I2.STATE3_il9r\, SET => 
        CLEAR_STAT_i_0, Q => \I2.STATE3_il8r\);
    
    \I2.DTO_16_1_IV_0_0_1L0R_1212\ : NOR2
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620__net_1\, 
        B => \I2.DT_TEMPl0r_net_1\, Y => 
        \I2.DTO_16_1_iv_0_0_1l0r_adt_net_35382_\);
    
    \I3.PIPEAl23r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_254_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl23r_net_1\);
    
    \I2.TDCDASl20r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl20r, Q => 
        \I2.TDCDASl20r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_a2_2\ : OR2
      port map(A => \I2.N_128_0_adt_net_55238_\, B => 
        \I2.N_3_0_adt_net_1070__net_1\, Y => \I2.N_128_0\);
    
    \I2.DTE_21_1_IV_0L16R_1268\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855116__net_1\, B => 
        \I2.EVNT_WORDl12r_net_1\, Y => 
        \I2.DTE_21_1l16r_adt_net_37819_\);
    
    \I2.OFFSET_37_20l5r\ : MUX2L
      port map(A => \I2.N_784\, B => \I2.N_776\, S => 
        \I2.PIPE7_DTL26R_357\, Y => \I2.N_792\);
    
    \I3.VDBoffb_54\ : OR3
      port map(A => \I3.VDBoffb_54_adt_net_162790_\, B => 
        \I3.VDBoffb_30l2r_adt_net_162749_\, C => 
        \I3.VDBoffb_30l2r_adt_net_162750_\, Y => 
        \I3.VDBoffb_54_net_1\);
    
    \I2.DTO_16_1_IV_0L4R_1198\ : AND2
      port map(A => \I2.DTO_1l4r\, B => \I2.N_196_52\, Y => 
        \I2.DTO_16_1l4r_adt_net_34374_\);
    
    \I2.DTO_9_ivl24r\ : AO21FTT
      port map(A => \I2.N_4283_i_0_adt_net_854968__net_1\, B => 
        \I2.DT_TEMPl24r_net_1\, C => 
        \I2.DTO_9l24r_adt_net_29802_\, Y => \I2.DTO_9l24r\);
    
    \I1.REG_74_0_IVL181R_2053\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l181r_adt_net_132215_\);
    
    \I3.un29_reg_ads_0_a2_0_a2\ : NAND2
      port map(A => \I3.VASl1r_net_1\, B => \I3.N_550\, Y => 
        \I3.N_562\);
    
    \I2.OFFSET_37_13l5r\ : MUX2L
      port map(A => \I2.N_728\, B => \I2.N_712\, S => 
        \I2.PIPE7_DTL25R_684\, Y => \I2.N_736\);
    
    \I2.TDCDASl12r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl12r, Q => 
        \I2.TDCDASl12r_net_1\);
    
    \I1.RAMDT_SPI_1l5r\ : DFFC
      port map(CLK => CLK_c, D => \FBOUTl5r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.RAMDT_SPI_1l5r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I108_Y\ : AO21
      port map(A => \I2.N321\, B => \I2.N436_adt_net_70670_\, C
         => \I2.N436_adt_net_70753_\, Y => \I2.N436\);
    
    \I3.VDBI_57_IVL4R_2251\ : AO21
      port map(A => \I3.PIPEAl4r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l4r_adt_net_144429_\, Y => 
        \I3.VDBi_57l4r_adt_net_144439_\);
    
    REGl264r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_165_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl264r\);
    
    \I1.REG_74_i_o2_i_0l364r\ : AND2FT
      port map(A => \I1.N_374\, B => \I1.N_273_6_i_0\, Y => 
        \I1.REG_74_i_o2_i_0l364r_net_1\);
    
    \I2.PIPE8_DT_21l13r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl13r_adt_net_854940__net_1\, B
         => \I2.PIPE8_DT_16l13r_net_1\, S => \I2.NWPIPE7_net_1\, 
        Y => \I2.PIPE8_DT_21l13r_net_1\);
    
    \I1.BITCNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BITCNT_316_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BITCNTl1r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I76_Y\ : AO21
      port map(A => \I2.N237_0\, B => \I2.N233\, C => \I2.N236\, 
        Y => \I2.N326_0\);
    
    \I2.PIPE4_DTl14r_1531\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL14R_638\);
    
    REGl235r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_136_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl235r\);
    
    REGl238r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_139_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl238r\);
    
    \I2.PIPE1_DT_730\ : MUX2L
      port map(A => \I2.PIPE1_DTl3r_net_1\, B => 
        \I2.PIPE1_DT_42l3r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854588__net_1\, 
        Y => \I2.PIPE1_DT_730_net_1\);
    
    \I1.ISCK_0_SQMUXA_0_0_A2_0_1761\ : NOR2
      port map(A => \I1.SSTATEL3R_713\, B => \I1.SSTATEL0R_755\, 
        Y => \I1.N_628_adt_net_107115_\);
    
    \I3.REGMAPL7R_2942\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un33_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL7R_459\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__2769\ : NAND3FFT
      port map(A => \I2.ENDF_837\, B => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149__net_1\, C => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_62\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__58\);
    
    \I2.G_EVNT_NUM_n7_i\ : NOR3
      port map(A => EV_RES_C_569, B => \I2.N_281\, C => 
        \I2.N_201_adt_net_855048__net_1\, Y => \I2.N_4639\);
    
    \I2.MIC_REG1l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_302_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1l1r_net_1\);
    
    \I3.VDBil0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_340_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil0r_net_1\);
    
    \I2.INT_ERRS_1022\ : OR2
      port map(A => \I2.TOKENB_TIMOUT_i_i\, B => 
        \I2.TOKENA_TIMOUT_net_1\, Y => 
        \I2.INT_ERRS_adt_net_22801_\);
    
    IACKB_pad : IB33
      port map(PAD => IACKB, Y => IACKB_c);
    
    \I2.ADEl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l14r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl14r);
    
    \I1.REG_3_sqmuxa_0_a2_0_817\ : NAND2FT
      port map(A => \I1.PAGECNTL9R_245\, B => \I1.N_238_RD1__314\, 
        Y => \I1.N_254_195\);
    
    \I3.CYCSF1_60\ : AOI21FTT
      port map(A => \I3.CYCSF1_net_1\, B => 
        \I3.N_306_adt_net_161608_\, C => \I3.ASBS_net_1\, Y => 
        \I3.CYCSF1_60_net_1\);
    
    \I3.REGMAPL21R_3025\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un86_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL21R_779\);
    
    \I1.REG_74_8_0_o4_a0_0l324r\ : OR2
      port map(A => \I1.PAGECNTL5R_308\, B => \I1.PAGECNTL6R_249\, 
        Y => \I1.REG_74_1_a0_0l228r\);
    
    \I2.DTE_21_1_IV_0L10R_1301\ : AND2
      port map(A => \I2.DTE_1l10r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1l10r_adt_net_38517_\);
    
    \I2.PIPE8_DT_21l24r\ : MUX2H
      port map(A => \I2.PIPE7_DTl24r_net_1\, B => 
        \I2.LSRAM_OUTl24r\, S => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l24r_net_1\);
    
    \I2.L2SERVl0r_1500\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_922_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL12R_607\);
    
    \I2.FCNTl2r\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_945_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.FCNTl2r_net_1\);
    
    \I2.OFFSET_37_18l6r\ : MUX2L
      port map(A => \REGl251r\, B => \REGl187r\, S => 
        \I2.PIPE7_DTL27R_77\, Y => \I2.N_777\);
    
    \I2.PIPE6_DT_465\ : MUX2H
      port map(A => \I2.PIPE5_DTl11r_net_1\, B => 
        \I2.PIPE6_DTl11r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_465_net_1\);
    
    \I2.un1_TOKENB_CNT_I_8\ : XOR2
      port map(A => TICKL0R_557, B => \I2.TOKENB_CNTl0r_net_1\, Y
         => \I2.DWACT_ADD_CI_0_partial_suml0r\);
    
    \I2.DTE_21_1_IVL15R_1277\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l15r\, C
         => \I2.DTE_21_1l15r_adt_net_37952_\, Y => 
        \I2.DTE_21_1l15r_adt_net_37953_\);
    
    \I2.DTO_1l9r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l9r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l9r_Rd1__net_1\);
    
    \I2.PIPE9_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_299_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl30r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L0R_2635\ : OR3
      port map(A => \I3.VDBoffa_31l0r_adt_net_164647_\, B => 
        \I3.VDBoffa_31l0r_adt_net_164643_\, C => 
        \I3.VDBoffa_31l0r_adt_net_164644_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164650_\);
    
    TDCDA_padl18r : IB33
      port map(PAD => TDCDA(18), Y => TDCDA_cl18r);
    
    \I3.VDBOFFB_30_IV_0L4R_2413\ : AO21
      port map(A => \REGl329r\, B => \I3.REGMAP_i_0_il38r_net_1\, 
        C => \I3.VDBoffb_30l4r_adt_net_162330_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162362_\);
    
    \I2.un1_PIPE1_DT_1_sqmuxa_2_0_a3\ : AND3FTT
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855240__net_1\, 
        B => \I2.STATE1l7r_net_1\, C => \I2.N_3879\, Y => 
        \I2.N_3902\);
    
    \I3.PIPEB_84\ : AO21
      port map(A => DPR_cl5r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_84_adt_net_160503_\, Y => 
        \I3.PIPEB_84_net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2563\ : OR3
      port map(A => \I3.VDBoffa_31l4r_adt_net_163887_\, B => 
        \I3.VDBoffa_31l4r_adt_net_163883_\, C => 
        \I3.VDBoffa_31l4r_adt_net_163884_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163890_\);
    
    \I2.OFFSET_37_17l6r\ : MUX2L
      port map(A => \I2.N_761\, B => \I2.N_753\, S => 
        \I2.PIPE7_DTL26R_352\, Y => \I2.N_769\);
    
    \I2.TDCGDAi\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TDCGDAi_672_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => TDCGDA_c);
    
    \I2.MIC_REG2_313\ : MUX2L
      port map(A => \I2.MIC_REG2_i_0_il5r_net_1\, B => 
        \I2.MIC_REG2_i_0_il4r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG2_313_net_1\);
    
    \I2.LEAD_FLAG6_7_i_0l4r\ : AOI21
      port map(A => \I2.N_215\, B => \I2.N_483\, C => \I2.N_222\, 
        Y => \I2.N_4531_adt_net_64140_\);
    
    \I1.REG_1_247\ : MUX2H
      port map(A => \REGl346r\, B => \I1.REG_74l346r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_247_net_1\);
    
    SDAA_pad : IOB33PH
      port map(PAD => SDAA, A => \I5.SDAout_net_1\, EN => 
        un1_sdaa_0_a2, Y => SDAA_in);
    
    \I2.MIC_ERR_REGSl34r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_363_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl34r_net_1\);
    
    \I2.DT_TEMP_7l20r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854240__net_1\, B => 
        \I2.DT_SRAMl20r_net_1\, Y => \I2.DT_TEMP_7l20r_net_1\);
    
    \I3.PIPEAl8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_239_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl8r_net_1\);
    
    \I1.N_65_adt_net_1433_\ : OR3
      port map(A => \I1.N_65_12\, B => 
        \I1.N_193_adt_net_118653__net_1\, C => \I1.N_97_6\, Y => 
        \I1.N_65_adt_net_1433__net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2592\ : AO21
      port map(A => \REGl175r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        C => \I3.VDBoffa_31l2r_adt_net_164226_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164261_\);
    
    \I2.DTO_16_1_iv_0_a2_2l21r\ : AND3
      port map(A => \I2.N_223_54\, B => \I2.N_4182\, C => 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_888__net_1\, Y => 
        \I2.N_196\);
    
    \I3.SINGCYC_1775\ : DFFC
      port map(CLK => CLK_c, D => \I3.SINGCYC_115_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.SINGCYC_881\);
    
    \I2.PIPE1_DT_42_1_IVL12R_1451\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl44r_net_1\, C => 
        \I2.PIPE1_DT_42l12r_adt_net_49438_\, Y => 
        \I2.PIPE1_DT_42l12r_adt_net_49456_\);
    
    \I1.PAGECNT_n2_0_0\ : OAI21
      port map(A => \I1.un1_sbyte13_1_i_1_adt_net_854524__net_1\, 
        B => \I1.N_390_i_i_0_i\, C => \I1.N_473_206\, Y => 
        \I1.PAGECNT_n2\);
    
    \I2.STATE1l12r_1540\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl6r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1L12R_647\);
    
    \I2.OFFSET_37_15l2r\ : MUX2L
      port map(A => \REGl231r\, B => \REGl167r\, S => 
        \I2.PIPE7_DTL27R_72\, Y => \I2.N_749\);
    
    \I2.L2TYPE_596\ : MUX2L
      port map(A => \I2.L2TYPEl7r_net_1\, B => \I2.N_4445\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_596_net_1\);
    
    \I2.DTO_16_1_IV_0L24R_1093\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.G_EVNT_NUMl8r_net_1\, Y
         => \I2.DTO_16_1l24r_adt_net_29860_\);
    
    \I2.LEAD_FLAG6l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LEAD_FLAG6_644_net_1\, CLR
         => CLEAR_STAT_i_0, Q => LEAD_FLAGl7r);
    
    \I3.VDBOFFB_30_IV_0L2R_2445\ : AO21
      port map(A => \REGl399r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l2r_adt_net_162694_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162738_\);
    
    \I1.REG_10_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_240\, B => \I1.N_259\, Y => 
        \I1.REG_10_sqmuxa\);
    
    \I5.TEMPDATAl3r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_77_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl3r_net_1\);
    
    \I5.SBYTE_9_il2r\ : MUX2L
      port map(A => \I5.COMMANDl10r_net_1\, B => 
        \I5.SBYTEl1r_net_1\, S => 
        \I5.N_155_0_adt_net_983__adt_net_855864__net_1\, Y => 
        \I5.N_18\);
    
    \I2.PIPE9_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_296_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl27r_net_1\);
    
    \I3.VDBi_57_iv_0_0_m2l0r\ : MUX2L
      port map(A => REGl18r, B => \I3.N_2063_i\, S => 
        \I3.REGMAPl50r_net_1\, Y => \I3.N_1923\);
    
    \I3.PIPEA_8l15r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854468__net_1\, B => 
        \I3.N_224\, Y => \I3.PIPEA_8l15r_net_1\);
    
    \I1.PAGECNTl6r_adt_net_854924_\ : BFR
      port map(A => \I1.PAGECNTl6r_net_1\, Y => 
        \I1.PAGECNTl6r_adt_net_854924__net_1\);
    
    \I2.PIPE8_DT_21l23r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl23r\, B => 
        \I2.PIPE7_DTl23r_net_1\, S => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l23r_net_1\);
    
    \I5.TEMPDATA_76\ : MUX2L
      port map(A => \I5.TEMPDATAl2r_net_1\, B => REGl127r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_76_net_1\);
    
    \I3.un86_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_580\, B => \I3.N_553\, Y => 
        \I3.un86_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.I_1336_G_1\ : XOR2FT
      port map(A => \I2.OFFSETL1R_679\, B => \I2.SUB8L4R_709\, Y
         => \I2.G_1_5\);
    
    \I2.DTE_21_1_ivl11r\ : AO21
      port map(A => \I2.DTE_1l11r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, C => 
        \I2.DTE_21_1l11r_adt_net_38417_\, Y => \I2.DTE_21_1l11r\);
    
    \I1.REG_74_0_ivl284r\ : AO21
      port map(A => \REGl284r\, B => \I1.N_153\, C => 
        \I1.REG_74l284r_adt_net_122377_\, Y => 
        \I1.REG_74l284r_net_1\);
    
    \I5.sstate1se_10_0_0\ : AO21FTT
      port map(A => TICKl0r, B => \I5.sstate1l2r_net_1\, C => 
        \I5.N_73\, Y => \I5.sstate1_ns_el11r\);
    
    \I3.STATE1l9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL9R_11\);
    
    \I2.PIPE5_DT_703\ : MUX2L
      port map(A => \I2.PIPE5_DTl27r_net_1\, B => 
        \I2.PIPE4_DTl27r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_703_net_1\);
    
    \I3.un126_reg_ads_0_a2_1_a2\ : OR2
      port map(A => \I3.VASl5r_net_1\, B => \I3.VASl3r_net_1\, Y
         => \I3.N_553\);
    
    REGl275r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_176_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl275r\);
    
    \I3.VDBi_40_sn_m2_0_750\ : NOR2
      port map(A => \I3.REGMAPL57R_808\, B => 
        \I3.REGMAP_I_0_IL58R_803\, Y => \I3.N_354_0_128\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I31_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl10r\, B => 
        \I2.PIPE7_DTL10R_695\, Y => \I2.N261_0\);
    
    REGl278r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_179_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl278r\);
    
    \I3.REG3l4r_1169\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_129_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3L4R_431\);
    
    \I3.PIPEBl27r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_106_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl27r_net_1\);
    
    \I3.PIPEB_80\ : AO21
      port map(A => DPR_cl1r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_80_adt_net_160671_\, Y => 
        \I3.PIPEB_80_net_1\);
    
    \I2.TDCTRGi_1463\ : DFFC
      port map(CLK => CLK_c, D => \I2.TDCTRGi_266_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => TDCTRG_C_570);
    
    \I1.REG_74_0_IVL354R_1859\ : NOR2FT
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_24_sqmuxa_adt_net_854776__net_1\, Y => 
        \I1.REG_74l354r_adt_net_115773_\);
    
    DTE_padl24r : IOB33PH
      port map(PAD => DTE(24), A => \I2.DTE_1l24r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl24r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I181_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_801\, B => 
        \I2.PIPE4_DTl11r_net_1\, Y => 
        \I2.ADD_21x21_fast_I181_Y_0_0\);
    
    \I2.ADE_4l13r\ : MUX2L
      port map(A => \I2.RPAGEl13r\, B => \I2.WPAGEl13r_net_1\, S
         => NOESRAME_C_243, Y => \I2.ADE_4l13r_net_1\);
    
    \I2.REG_1_c11_i\ : OAI21TTF
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => \I2.N_3856\, C => \I2.N_3840_adt_net_101218_\, Y => 
        \I2.N_3840\);
    
    \I1.REG_74_0_ivl332r\ : AO21
      port map(A => \REGl332r\, B => \I1.N_201\, C => 
        \I1.REG_74l332r_adt_net_117916_\, Y => 
        \I1.REG_74l332r_net_1\);
    
    \I3.un186_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.N_558\, B => \I3.N_580\, Y => 
        \I3.un186_reg_ads_0_a2_1_a3_net_1\);
    
    \I2.STATE2L3R_2921\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl2r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L3R_438\);
    
    DTE_padl30r : IOB33PH
      port map(PAD => DTE(30), A => \I2.DTE_1l30r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl30r);
    
    \I2.N507_adt_net_56246_\ : AND3
      port map(A => \I2.N_107\, B => \I2.N_128\, C => 
        \I2.N507_adt_net_258084__net_1\, Y => 
        \I2.N507_adt_net_56246__net_1\);
    
    \I2.FID_7_0_IVL31R_974\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl79r, C => 
        \I2.FID_7l31r_adt_net_18457_\, Y => 
        \I2.FID_7l31r_adt_net_18465_\);
    
    \I1.N_305_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_305_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_305_Rd1__net_1\);
    
    \I2.TDC_653\ : MUX2H
      port map(A => \I2.TDCl3r_net_1\, B => 
        \I2.RAMAD1_12l16r_net_1\, S => 
        \I2.un1_FIRST_TDC_1_sqmuxa_0_adt_net_1038__net_1\, Y => 
        \I2.TDC_653_net_1\);
    
    \I2.PIPE5_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_696_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl20r_net_1\);
    
    \I2.PIPE5_DT_692\ : MUX2L
      port map(A => \I2.PIPE5_DTl16r_net_1\, B => 
        \I2.PIPE5_DT_6l16r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_692_net_1\);
    
    \I1.COMMAND_1609\ : DFFS
      port map(CLK => CLK_c, D => \I1.COMMAND_52_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.COMMAND_716\);
    
    \I2.ROFFSET_n9\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\, B => 
        \I2.ROFFSET_n9_tz_i\, Y => \I2.ROFFSET_n9_net_1\);
    
    \I2.G_EVNT_NUM_932\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl2r_net_1\, B => \I2.N_4342\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_932_net_1\);
    
    \I5.PULSE_FL_53\ : AO21
      port map(A => \I5.sstate1l13r_net_1\, B => 
        \I5.PULSE_FL_net_1\, C => \I5.PULSE_I2C_net_1\, Y => 
        \I5.PULSE_FL_53_net_1\);
    
    \I3.VDBi_57_0_ivl12r\ : AO21FTT
      port map(A => \I3.N_1905_1_adt_net_855380__net_1\, B => 
        \I3.VDBi_40l12r_net_1\, C => 
        \I3.VDBi_57l12r_adt_net_140998_\, Y => \I3.VDBi_57l12r\);
    
    \I2.EVNT_NUMl4r_1491\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_959_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUML4R_598\);
    
    \I3.UN1_SINGCYC8_I_0_O3_2312\ : NOR3
      port map(A => AMB_cl1r, B => AMB_cl0r, C => \I3.N_2055\, Y
         => \I3.N_80_adt_net_159051_\);
    
    \I2.STATE1_ns_i_o2l9r_967\ : OR3
      port map(A => FLUSH, B => \I2.FCNT_c1\, C => 
        \I2.FCNTL2R_892\, Y => \I2.N_3272_345\);
    
    \I3.REG_1l62r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_163_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl62r);
    
    \I2.RAMDT4L12R_3075\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_829\);
    
    \I2.PIPE9_DTl30r_1561\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_299_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTL30R_668\);
    
    \I2.PIPE10_DT_631\ : MUX2L
      port map(A => \I2.PIPE10_DTl26r_net_1\, B => 
        \I2.PIPE9_DTl26r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_631_net_1\);
    
    \I5.REG_1l421r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_34_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl421r);
    
    \I2.DT_SRAM_0_il27r\ : MUX2L
      port map(A => \I2.PIPE10_DTl27r_net_1\, B => 
        \I2.PIPE5_DTl27r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854204__net_1\, Y => 
        \I2.DT_SRAM_0_il27r_net_1\);
    
    \I2.STATE5_ns_0_a5l3r\ : OR2FT
      port map(A => \I2.STATE5l0r_net_1\, B => 
        \I2.W_ERR_WORDS_net_1\, Y => \I2.N_4332\);
    
    \I3.un7_cycs_i\ : OR2FT
      port map(A => \I3.CYCS_net_1\, B => \I3.ASBS_net_1\, Y => 
        \I3.un7_cycs_i_net_1\);
    
    \I2.DTE_21_1_0_iv_1l30r\ : OAI21FTF
      port map(A => \I2.STATE2L3R_440\, B => 
        \I2.DTO_9_ivl30r_net_1\, C => 
        \I2.DTE_21_1_0_iv_1l30r_adt_net_36511_\, Y => 
        \I2.DTE_21_1_0_iv_1l30r_net_1\);
    
    \I3.REGMAPl33r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un146_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPl33r_net_1\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2272\ : AO21
      port map(A => REGl82r, B => \I3.REGMAPl12r_net_1\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146347_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146304_\);
    
    \I3.REG2l7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG2_148_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l7r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2616\ : OR3
      port map(A => \I3.VDBoffa_31l1r_adt_net_164455_\, B => 
        \I3.VDBoffa_31l1r_adt_net_164449_\, C => 
        \I3.VDBoffa_31l1r_adt_net_164450_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164459_\);
    
    \I2.DT_SRAMl28r\ : MUX2L
      port map(A => \I2.N_896\, B => \I2.PIPE2_DTl28r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672__net_1\, 
        Y => \I2.DT_SRAMl28r_net_1\);
    
    \I2.DTO_9_ivl1r\ : OAI21TTF
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl1r_net_1\, C => 
        \I2.DTO_9_ivl1r_adt_net_35072_\, Y => 
        \I2.DTO_9_ivl1r_net_1\);
    
    \I1.REG_74_0_iv_0_0l259r\ : AO21
      port map(A => \REGl259r\, B => \I1.N_658\, C => 
        \I1.REG_74l259r_adt_net_124884_\, Y => \I1.REG_74l259r\);
    
    TDCDA_padl25r : IB33
      port map(PAD => TDCDA(25), Y => TDCDA_cl25r);
    
    \I3.RAMAD_VMEl5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_29_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl5r);
    
    \I1.REG_74l268r\ : OR3FFT
      port map(A => \I1.REG_74_1l268r\, B => \I1.N_145_12\, C => 
        \I1.REG_14_sqmuxa\, Y => \I1.N_137\);
    
    \I1.REG_5_sqmuxa_0_a2_0_789\ : OR3FTT
      port map(A => \I1.PAGECNTL7R_526\, B => 
        \I1.PAGECNTl8r_net_1\, C => 
        \I1.N_1169_adt_net_854812__net_1\, Y => \I1.N_243_167\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I181_Y\ : XOR2
      port map(A => \I2.N519\, B => \I2.ADD_21x21_fast_I181_Y_0\, 
        Y => \I2.un27_pipe5_dt0l11r\);
    
    \I3.STATE2_ns_0l0r\ : OAI21TTF
      port map(A => \I3.N_1896\, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854456__net_1\, C => 
        \I3.STATE2_nsl0r_adt_net_136048_\, Y => \I3.STATE2_nsl0r\);
    
    \I2.NWPIPE7_1582\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE6_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE7_689\);
    
    \I2.NWPIPE9\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE8_I_0_I_0_0_6\, SET
         => CLEAR_STAT_i_0, Q => \I2.NWPIPE9_0_7\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I140_Y_0_753\ : AO21FTF
      port map(A => \I2.N_74_I_0_I_132\, B => 
        \I2.N519_adt_net_54631_\, C => \I2.N_70\, Y => 
        \I2.N519_131\);
    
    \I1.SSTATEL10R_2911\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_43_i_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL10R_380\);
    
    \I2.N_2826_1_ADT_NET_794__2888\ : OAI21FTF
      port map(A => \I2.N_4261_304\, B => \I2.N_4282\, C => 
        \I2.N_2826_1_adt_net_40744__net_1\, Y => 
        \I2.N_2826_1_ADT_NET_794__329\);
    
    \I2.MIC_ERR_REGSl38r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_367_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl38r_net_1\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2385\ : AND2
      port map(A => \REGl354r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162128_\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854504_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854512__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854504__net_1\);
    
    \I2.LSRAM_IN_392\ : MUX2L
      port map(A => \I2.PIPE5_DTl8r_net_1\, B => 
        \I2.LSRAM_INl8r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_392_net_1\);
    
    \I3.REGMAPl50r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un221_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl50r_net_1\);
    
    \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__2746\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__19\);
    
    \I2.OFFSET_37_23l5r\ : MUX2L
      port map(A => \REGl274r\, B => \REGl210r\, S => 
        \I2.PIPE7_DTL27R_88\, Y => \I2.N_816\);
    
    \I2.DTE_1l8r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l8r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l8r_Rd1__net_1\);
    
    \I2.PIPE5_DT_6_0L28R_1541\ : AND2
      port map(A => \I2.dataout_0_adt_net_855804__net_1\, B => 
        \I2.dataout_1\, Y => \I2.PIPE5_DT_6l28r_adt_net_53820_\);
    
    \I2.OFFSET_37_4l4r\ : MUX2L
      port map(A => \REGl369r\, B => \REGl305r\, S => 
        \I2.PIPE7_DTL27R_70\, Y => \I2.N_663\);
    
    \I2.PIPE1_DT_42_1_IVL17R_1407\ : NOR2FT
      port map(A => REGl421r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, Y => 
        \I2.PIPE1_DT_42l17r_adt_net_47643_\);
    
    \I1.REG_74_0_ivl282r\ : AO21
      port map(A => \REGl282r\, B => \I1.N_153\, C => 
        \I1.REG_74l282r_adt_net_122549_\, Y => \I1.REG_74l282r\);
    
    \I2.PIPE6_DT_482\ : MUX2H
      port map(A => \I2.PIPE5_DTl28r_net_1\, B => 
        \I2.PIPE6_DTl28r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_482_net_1\);
    
    \I3.STBMIC_78\ : MUX2H
      port map(A => STBMIC_c, B => \I3.STATE1_IPL8R_10\, S => 
        \I3.N_1902\, Y => \I3.STBMIC_78_net_1\);
    
    \I2.PIPE6_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_479_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl25r_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl23r\ : OR3
      port map(A => \I2.PIPE1_DT_42l23r_adt_net_46641_\, B => 
        \I2.PIPE1_DT_42l23r_adt_net_46653_\, C => 
        \I2.PIPE1_DT_42l23r_adt_net_46654_\, Y => 
        \I2.PIPE1_DT_42l23r\);
    
    \I3.VDBi_57l2r_adt_net_145285_\ : AND2
      port map(A => REGl408r, B => \I3.REGMAPl55r_net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145285__net_1\);
    
    \I2.ROFFSETl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_908_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl10r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I176_Y\ : XOR2FT
      port map(A => \I2.N_31\, B => \I2.ADD_21x21_fast_I176_Y_0\, 
        Y => \I2.un27_pipe5_dt0l6r\);
    
    \I1.SBYTE_65\ : MUX2L
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.N_1194\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_65_0\);
    
    \I1.REG_74_0_iv_0l273r\ : AO21
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, C => 
        \I1.REG_74l273r_adt_net_123560_\, Y => \I1.REG_74l273r\);
    
    \I2.FID_7_0_IVL26R_984\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl74r, C => 
        \I2.FID_7l26r_adt_net_18927_\, Y => 
        \I2.FID_7l26r_adt_net_18935_\);
    
    \I2.PIPE4_DTl2r_1251\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL2R_513\);
    
    \I2.PIPE2_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl19r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl19r_net_1\);
    
    \I1.REG_74_0_ivl278r\ : AO21
      port map(A => \REGl278r\, B => \I1.N_153\, C => 
        \I1.REG_74l278r_adt_net_122893_\, Y => \I1.REG_74l278r\);
    
    \I1.REG_74_0_ivl398r\ : AO21
      port map(A => \REGl398r\, B => \I1.N_273\, C => 
        \I1.REG_74l398r_adt_net_110272_\, Y => \I1.REG_74l398r\);
    
    \I2.LSRAM_IN_406\ : MUX2L
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => 
        \I2.LSRAM_INl22r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_406_net_1\);
    
    \I2.L2TYPEl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_593_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl4r_net_1\);
    
    MSERCLK_pad : IB33
      port map(PAD => MSERCLK, Y => MSERCLK_c);
    
    \I3.VDBi_57_0_iv_0_a3_9_1l15r\ : NOR3
      port map(A => \I3.N_2015\, B => \I3.N_1905\, C => 
        \I3.N_2033\, Y => \I3.N_403_1\);
    
    \I2.PIPE8_DT_536\ : MUX2L
      port map(A => \I2.PIPE8_DTl8r_net_1\, B => 
        \I2.PIPE8_DT_21l8r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_536_net_1\);
    
    \I3.un7_cycs_0_a3_0_a3\ : NOR2FT
      port map(A => \I3.CYCS_net_1\, B => \I3.ASBS_net_1\, Y => 
        \I3.un7_cycs_0_a3_0_a3_net_1\);
    
    \I2.ROFFSETe_0_adt_net_27185_\ : OAI21FTF
      port map(A => \I2.STATE3l1r_net_1\, B => \I2.N_3015\, C => 
        \I2.ROFFSETe_0_adt_net_27184__net_1\, Y => 
        \I2.ROFFSETe_0_adt_net_27185__net_1\);
    
    \I2.OFFSET_37_28l6r\ : MUX2L
      port map(A => \I2.N_849\, B => \I2.N_801\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_857\);
    
    \I1.REG_74_0_IVL237R_1989\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_10_sqmuxa_adt_net_854720__net_1\, Y => 
        \I1.REG_74l237r_adt_net_126985_\);
    
    \I2.DT_TEMPl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_788_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl27r_net_1\);
    
    \I2.PIPE8_DT_21l19r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl19r\, B => 
        \I2.PIPE8_DT_16l19r_net_1\, S => \I2.NWPIPE7_net_1\, Y
         => \I2.PIPE8_DT_21l19r_net_1\);
    
    \I2.MIC_REG3L1R_2937\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_318_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3L1R_454\);
    
    \I3.VDBoffbl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffb_53_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffbl1r_net_1\);
    
    \I5.sstate1se_7_0_0\ : OR2
      port map(A => \I5.sstate1_ns_el8r_adt_net_8886_\, B => 
        \I5.sstate1_ns_el8r_adt_net_8891_\, Y => 
        \I5.sstate1_ns_el8r\);
    
    \I5.REG_1l117r_1128\ : DFFS
      port map(CLK => CLK_c, D => \I5.REG_1_54_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => REGL117R_390);
    
    TDCDA_padl26r : IB33
      port map(PAD => TDCDA(26), Y => TDCDA_cl26r);
    
    REGl224r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_125_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl224r\);
    
    \I5.SSTATE1SE_13_0_899\ : OAI21FTF
      port map(A => \I5.sstate1l0r_net_1\, B => 
        \I5.COMMANDl2r_net_1\, C => \I5.sstate1l9r_net_1\, Y => 
        \I5.sstate1_ns_el0r_adt_net_7898_\);
    
    \I5.REG_1_18\ : MUX2H
      port map(A => REGl132r, B => REGl435r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\, Y
         => \I5.REG_1_18_net_1\);
    
    \I3.PIPEA_247\ : MUX2L
      port map(A => \I3.PIPEAl16r_net_1\, B => 
        \I3.PIPEA_8l16r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854664__net_1\, Y
         => \I3.PIPEA_247_net_1\);
    
    \I2.OFFSET_37_27l6r\ : MUX2L
      port map(A => \I2.N_841\, B => \I2.N_825\, S => 
        \I2.PIPE7_DTL25R_687\, Y => \I2.N_849\);
    
    \I2.L2TYPE_4_IL2R_1637\ : NAND2
      port map(A => \I2.N_4456\, B => \I2.N_4461\, Y => 
        \I2.N_4450_adt_net_68435_\);
    
    \I2.STATE1l13r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_il5r_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.STATE1l13r_net_1\);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_501\ : MUX2L
      port map(A => \I2.LSRAM_RADDRil2r_net_1\, B => 
        \I2.PIPE4_DTl23r_net_1\, S => \I2.N_4642\, Y => 
        \I2.LSRAM_RADDRi_501\);
    
    \I2.MIC_ERR_REGS_374\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl46r_net_1\, B => 
        \I2.MIC_ERR_REGSl45r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_374_net_1\);
    
    \I3.REGMAPL41R_2983\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un186_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL41R_530\);
    
    \I2.DTE_cl_96_iv_0_i_0l31r\ : OA21FTT
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.N_2838_i_0\, C
         => \I2.N_4293\, Y => \I2.N_2822\);
    
    \I2.BNCID_VECTria_11_0\ : AND2
      port map(A => \I2.BNCID_VECTra15_1_net_1\, B => 
        \I2.BNCID_VECTro_11\, Y => \I2.BNCID_VECTria_11_0_i\);
    
    \I2.RAMDT4L12R_3039\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_793\);
    
    \I2.PIPE9_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_270_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl1r_net_1\);
    
    \I2.PIPE9_DT_281\ : MUX2L
      port map(A => \I2.PIPE9_DTl12r_net_1\, B => 
        \I2.PIPE8_DTl12r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_281_net_1\);
    
    \I2.SUB8_512\ : MUX2H
      port map(A => \I2.SUB8l9r_net_1\, B => \I2.SUB8_2l9r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855144__net_1\, Y => 
        \I2.SUB8_512_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I178_Y_2731\ : AO21
      port map(A => \I2.N479_adt_net_642172_\, B => 
        \I2.N479_adt_net_642225_\, C => \I2.N479_adt_net_642266_\, 
        Y => \I2.N479_adt_net_538261_\);
    
    \I5.BITCNTe_0_a2_0_a2_0\ : OR3FFT
      port map(A => TICKL0R_3, B => \I5.COMMANDl0r_net_1\, C => 
        \I5.N_64_adt_net_855868__net_1\, Y => \I5.N_130\);
    
    \I2.LEAD_FLAG6_1_SQMUXA_I_1598\ : AND3FTT
      port map(A => \I2.NWPIPE5_net_1\, B => 
        \I2.PIPE5_DTl31r_net_1\, C => \I2.N_4551\, Y => 
        \I2.N_4527_adt_net_63801_\);
    
    \I2.DTE_21_1_IV_2L0R_1345\ : OAI21TTF
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855208__net_1\, 
        B => \I2.DT_TEMPl0r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39723_\, Y => 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39732_\);
    
    \I3.RAMAD_VME_33\ : MUX2H
      port map(A => RAMAD_VMEl9r, B => \I3.REGl92r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_33_net_1\);
    
    \I2.OFFSET_37_25l2r\ : MUX2L
      port map(A => \REGl255r\, B => \REGl191r\, S => 
        \I2.PIPE7_DTL27R_91\, Y => \I2.N_829\);
    
    \I2.STATE2l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl3r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2l2r_net_1\);
    
    \I2.PIPE6_DT_471\ : MUX2H
      port map(A => \I2.PIPE5_DTl17r_net_1\, B => 
        \I2.PIPE6_DTl17r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_471_net_1\);
    
    \I2.DTO_16_1_IVL11R_1167\ : AO21
      port map(A => \I2.N_182_adt_net_1007__net_1\, B => 
        \I2.DT_SRAMl11r_net_1\, C => 
        \I2.DTO_16_1l11r_adt_net_32878_\, Y => 
        \I2.DTO_16_1l11r_adt_net_32879_\);
    
    \I2.WOFFSETl2r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.WOFFSETl2r_adt_net_854984__net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl2r_Rd1__net_1\);
    
    \I2.TDCDBSl14r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl14r, Q => 
        \I2.TDCDBSl14r_net_1\);
    
    \I1.REG_74_0_iv_0_0l251r\ : AO21
      port map(A => \REGl251r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l251r_adt_net_125691_\, Y => \I1.REG_74l251r\);
    
    \I2.DTE_21_1_IV_0L27R_1238\ : AO21FTT
      port map(A => \I2.N_4647\, B => 
        \I2.N_199_0_adt_net_1054__net_1\, C => 
        \I2.DTE_21_1l27r_adt_net_36849_\, Y => 
        \I2.DTE_21_1l27r_adt_net_36860_\);
    
    \I2.DTO_16_1_IV_0L5R_1195\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608__net_1\, 
        B => \I2.DT_TEMPl5r_net_1\, C => 
        \I2.DTO_16_1l5r_adt_net_34192_\, Y => 
        \I2.DTO_16_1l5r_adt_net_34198_\);
    
    \I1.sstatel6r_1155\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl4r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL6R_417\);
    
    \I2.ROFFSET_c6\ : NOR2FT
      port map(A => \I2.ROFFSETl6r_net_1\, B => 
        \I2.ROFFSET_c5_net_1\, Y => \I2.ROFFSET_c6_net_1\);
    
    \I3.REGMAPl1r_1617\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un10_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL1R_724\);
    
    \I3.VADm_0_a3l24r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl24r_net_1\, Y => \I3.VADml24r\);
    
    \I2.UN1_REG80_I_1696\ : NOR2
      port map(A => REG_i_0_il42r, B => REGl39r, Y => 
        \I2.N_3824_adt_net_90285_\);
    
    BNC_RESIN_pad : IB33
      port map(PAD => BNC_RESIN, Y => BNC_RESIN_c);
    
    \I2.STATE3l6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_ns_il7r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3l6r_net_1\);
    
    \I1.REG_74l340r\ : NAND2FT
      port map(A => \I1.REG_21_sqmuxa\, B => \I1.REG_74_0l332r\, 
        Y => \I1.N_209\);
    
    \I3.REGMAPl9r_adt_net_854312_\ : BFR
      port map(A => \I3.REGMAPl9r_adt_net_854316__net_1\, Y => 
        \I3.REGMAPl9r_adt_net_854312__net_1\);
    
    \I2.L2RF1\ : DFFC
      port map(CLK => CLK_c, D => L2R_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L2RF1_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I3_G0N_0_o3\ : NAND2
      port map(A => \I2.RAMDT4L10R_442\, B => 
        \I2.PIPE4_DTl3r_net_1\, Y => \I2.N_17_0\);
    
    \I5.DATA_12_ivl1r\ : AO21FTT
      port map(A => TICKl0r, B => REGl118r, C => 
        \I5.DATA_12_ivl1r_adt_net_14302_\, Y => 
        \I5.DATA_12_ivl1r_net_1\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2273\ : NOR3FFT
      port map(A => REGl80r, B => \I3.REGMAPl11r_net_1\, C => 
        \I3.REGMAPl12r_net_1\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146347_\);
    
    \I2.DTE_21_1_IV_0_IL25R_1244\ : AO21
      port map(A => \I2.DT_SRAMl25r_net_1\, B => 
        \I2.N_199_0_ADT_NET_1054__37\, C => 
        \I2.N_4644_adt_net_37053_\, Y => 
        \I2.N_4644_adt_net_37064_\);
    
    \I2.OFFSET_37_14l6r\ : MUX2L
      port map(A => \I2.N_737\, B => \I2.N_689\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_745\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I136_Y_0_o2_m4_e_2\ : AND2
      port map(A => \I2.N_53_0\, B => \I2.N_92_0\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_2_adt_net_56513_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I30_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl9r\, B => \I2.PIPE7_DTL9R_696\, 
        Y => \I2.N258_0\);
    
    \I3.VDBi_23l1r_adt_net_145542_\ : OR2
      port map(A => \I3.VDBi_23l1r_adt_net_145530__net_1\, B => 
        \I3.VDBi_23l1r_adt_net_145532__net_1\, Y => 
        \I3.VDBi_23l1r_adt_net_145542__net_1\);
    
    \I1.un1_sbyte13_1_i_1_adt_net_854524_\ : BFR
      port map(A => \I1.un1_sbyte13_1_i_1\, Y => 
        \I1.un1_sbyte13_1_i_1_adt_net_854524__net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2533\ : AND2
      port map(A => \REGl250r\, B => \I3.REGMAPl28r_net_1\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163664_\);
    
    \I2.DTOSl16r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl16r, Q => 
        \I2.DTOSl16r_net_1\);
    
    \I3.VDBoffa_31_iv_0l0r\ : AND2
      port map(A => \REGl205r\, B => 
        \I3.REGMAPl23r_adt_net_855016__net_1\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164594_\);
    
    \I2.PIPE8_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_543_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl15r_net_1\);
    
    \I1.REG_74_0_IVL327R_1889\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l327r_adt_net_118346_\);
    
    \I1.N_591_1_adt_net_106236_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => 
        \I1.N_591_1_adt_net_106236_Ra1_\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.N_591_1_adt_net_106236_Rd1__net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2547\ : AND2
      port map(A => \REGl241r\, B => \I3.REGMAPl27r_net_1\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163838_\);
    
    \I2.DTO_cl_0_sqmuxa_0_adt_net_855204_\ : BFR
      port map(A => \I2.DTO_cl_0_sqmuxa_0\, Y => 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\);
    
    \I2.DTE_cl_0_sqmuxa_2_adt_net_20061_\ : AO21TTF
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__149\, B => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_19952__net_1\, C => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_160\, Y => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20061__net_1\);
    
    \I1.N_349_RD1__2969\ : DFFC
      port map(CLK => CLK_c, D => \I1.N_349_Ra1_\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.N_349_RD1__486\);
    
    \I3.VDBm_0l17r\ : MUX2L
      port map(A => \I3.PIPEAl17r_net_1\, B => 
        \I3.PIPEBl17r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_159\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I166_Y_1688\ : NAND3FTT
      port map(A => \I2.N356\, B => \I2.N400_adt_net_88380_\, C
         => \I2.N411_adt_net_4092__net_1\, Y => 
        \I2.N501_i_adt_net_88539_\);
    
    \I3.VDBOFFB_58_2384\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl6r_net_1\, Y => 
        \I3.VDBoffb_58_adt_net_162030_\);
    
    \I3.UN10_TCNT2_2108\ : OR3
      port map(A => \I3.TCNT2_i_0_il2r_net_1\, B => 
        \I3.TCNT2l1r_net_1\, C => \I3.un10_tcnt2_adt_net_135288_\, 
        Y => \I3.un10_tcnt2_adt_net_135291_\);
    
    \I2.TOKENTOB_RES_649\ : AO21TTF
      port map(A => \I2.TOKENTOB_RES_net_1\, B => \I2.N_3302\, C
         => \I2.un1_STATE1_27\, Y => \I2.TOKENTOB_RES_649_net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2549\ : AND2
      port map(A => \REGl217r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.VDBoffa_31l4r_adt_net_163846_\);
    
    \I3.REG_1l153r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_201_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl153r\);
    
    \I2.L2SERVl2r_1509\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_920_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL14R_616\);
    
    \I2.DTE_21_1_iv_0l26r\ : AO21
      port map(A => \I2.DTE_1l26r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.DTE_21_1l26r_adt_net_36963_\, Y => \I2.DTE_21_1l26r\);
    
    \I2.PIPE8_DT_21l8r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl8r\, B => \I2.N_574\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l8r_net_1\);
    
    \I2.SUB9_572\ : MUX2H
      port map(A => \I2.SUB9l4r_net_1\, B => \I2.SUB9_1l4r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_572_net_1\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854496_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854512__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854496__net_1\);
    
    \I3.PIPEB_95\ : AO21
      port map(A => DPR_cl16r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_95_adt_net_160041_\, Y => 
        \I3.PIPEB_95_net_1\);
    
    \I2.OFFSET_37_11l1r\ : MUX2L
      port map(A => \REGl374r\, B => \REGl310r\, S => 
        \I2.PIPE7_DTL27R_84\, Y => \I2.N_716\);
    
    \I3.REG_1_290\ : MUX2L
      port map(A => VDB_inl8r, B => REGl109r, S => 
        \I3.N_318_adt_net_855888__net_1\, Y => \I3.REG_1_290_0\);
    
    \I1.REG_1_129\ : MUX2H
      port map(A => \REGl228r\, B => \I1.REG_74l228r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\, Y
         => \I1.REG_1_129_net_1\);
    
    \I3.un1_REGMAP_30_0_a2_997\ : AND3
      port map(A => \I3.un1_REGMAP_30_adt_net_134454_\, B => 
        \I3.un1_REGMAP_30_0_a2_0_net_1\, C => \I3.N_68\, Y => 
        \I3.UN1_REGMAP_30_375\);
    
    \I2.PIPE5_DT_679\ : MUX2L
      port map(A => \I2.PIPE5_DTl3r_net_1\, B => 
        \I2.PIPE5_DT_6l3r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_679_net_1\);
    
    \I2.STATE1l6r_1523\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3875_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1L6R_630\);
    
    \I1.REG_74_0_iv_0l370r\ : AO21
      port map(A => \REGl370r\, B => \I1.N_660\, C => 
        \I1.REG_74l370r_adt_net_113482_\, Y => \I1.REG_74l370r\);
    
    \I2.STATE1_0_sqmuxa_0_a3_0_a3_0\ : OR2
      port map(A => \I2.CHAINA_EN244_i_adt_net_855260__net_1\, B
         => \I2.N_3287_i_0\, Y => \I2.STATE1_ns_0l5r\);
    
    \I2.ADOl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l14r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl14r);
    
    \I2.TDCDBSl17r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl17r, Q => 
        \I2.TDCDBSl17r_net_1\);
    
    SP4_pad : OB33PH
      port map(PAD => SP4, A => \GND\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I136_Y_0_O2_M4_2_2664\ : 
        OR2
      port map(A => \I2.PIPE4_DTL10R_851\, B => 
        \I2.PIPE4_DTL9R_847\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_2_i_adt_net_271662_\);
    
    \I2.DTO_9_iv_0_m2l5r\ : MUX2L
      port map(A => \I2.DTE_2_1l5r_net_1\, B => \I2.N_4266\, S
         => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996__net_1\, 
        Y => \I2.DTO_9l5r\);
    
    \I1.PAGECNTLDE_0_A2_0_1_1756\ : NAND2
      port map(A => \I1.BYTECNT_306_net_1\, B => 
        \I1.sstate_nsl6r\, Y => \I1.N_591_1_adt_net_106236_Ra1_\);
    
    \I1.REG_74_0_ivl182r\ : AO21
      port map(A => \REGl182r\, B => \I1.N_57\, C => 
        \I1.REG_74l182r_adt_net_132129_\, Y => \I1.REG_74l182r\);
    
    \I3.VDBOFFB_30_IV_0L0R_2484\ : AO21
      port map(A => \REGl293r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l0r_adt_net_163086_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163121_\);
    
    \I2.TRGSERV_2_I_15\ : XOR2
      port map(A => \I2.DWACT_ADD_CI_0_TMP_0l0r\, B => 
        \I2.TRGSERVl1r_net_1\, Y => \I2.TRGSERV_2l1r\);
    
    \I2.PIPE5_DT_6l8r\ : MUX2L
      port map(A => 
        \I2.PIPE4_DTl8r_adt_net_854556__adt_net_855024__net_1\, B
         => \I2.N_1077\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855612__net_1\, Y => 
        \I2.PIPE5_DT_6l8r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I183_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_801\, B => 
        \I2.PIPE4_DTl13r_net_1\, Y => 
        \I2.ADD_21x21_fast_I183_Y_0_0\);
    
    \I2.N_4534_adt_net_1171_\ : AO21FTT
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_4673\, C
         => LEAD_FLAGl1r, Y => \I2.N_4534_adt_net_1171__net_1\);
    
    \I3.REG_1l86r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_267_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl86r);
    
    \I2.DTE_21_1_IV_0L27R_1237\ : AND2
      port map(A => \I2.DT_TEMPl27r_net_1\, B => \I2.N_4038_233\, 
        Y => \I2.DTE_21_1l27r_adt_net_36849_\);
    
    \I1.REG_74_0_ivl228r\ : AO21
      port map(A => \REGl228r\, B => \I1.N_97\, C => 
        \I1.REG_74l228r_adt_net_127964_\, Y => 
        \I1.REG_74l228r_net_1\);
    
    \I2.resyn_0_I2_GIROT_452\ : MUX2L
      port map(A => TDCTRG_c, B => \I2.GIROT_net_1\, S => 
        \I2.N_3760\, Y => \I2.GIROT_452\);
    
    \I2.FID_7_0_IVL21R_993\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl21r_net_1\, 
        Y => \I2.FID_7l21r_adt_net_19397_\);
    
    \I3.un47_reg_ads_0_a2_0_a3_1\ : OR3
      port map(A => \I3.VASl12r_net_1\, B => \I3.VASl2r_net_1\, C
         => \I3.N_555\, Y => \I3.un47_reg_ads_1\);
    
    \I2.WOFFSETl3r_adt_net_854988_\ : BFR
      port map(A => \I2.WOFFSETl3r\, Y => 
        \I2.WOFFSETl3r_adt_net_854988__net_1\);
    
    \I2.LSRAM_IN_388\ : MUX2L
      port map(A => \I2.PIPE5_DTl4r_net_1\, B => 
        \I2.LSRAM_INl4r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_388_net_1\);
    
    \I2.PIPE10_DT_632\ : MUX2L
      port map(A => \I2.PIPE10_DTl27r_net_1\, B => 
        \I2.PIPE9_DTl27r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_632_net_1\);
    
    \I2.DTE_21_1_IVL15R_1275\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, 
        B => \I2.DT_TEMPl15r_net_1\, C => 
        \I2.DTE_21_1l15r_adt_net_37935_\, Y => 
        \I2.DTE_21_1l15r_adt_net_37950_\);
    
    \I3.PIPEA_8l25r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854460__net_1\, B => 
        \I3.N_234\, Y => \I3.PIPEA_8l25r_net_1\);
    
    \I2.un1_STATE1_39_6\ : OR2
      port map(A => \I2.un1_STATE1_39_6_i_adt_net_52472_\, B => 
        \I2.un1_STATE1_39_6_i_adt_net_52473_\, Y => 
        \I2.un1_STATE1_39_6_i\);
    
    \I2.sram_empty_3\ : XOR2
      port map(A => \I2.RPAGEL15R_522\, B => \I2.WPAGEL15R_749\, 
        Y => \I2.sram_empty_3_i_0_i\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I183_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl13r_net_1\, Y => 
        \I2.ADD_21x21_fast_I183_Y_0\);
    
    \I3.VDBOFFB_30_IV_0L4R_2408\ : AND2
      port map(A => \REGl305r\, B => \I3.REGMAPl35r_net_1\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162338_\);
    
    \I1.REG_74_0_ivl391r\ : AO21
      port map(A => \REGl391r\, B => \I1.N_265\, C => 
        \I1.REG_74l391r_adt_net_110956_\, Y => \I1.REG_74l391r\);
    
    \I3.REG_1_160\ : MUX2L
      port map(A => VDB_inl11r, B => REGl59r, S => 
        \I3.N_1935_adt_net_855328__net_1\, Y => \I3.REG_1_160_0\);
    
    \I3.VDBm_0l8r\ : MUX2L
      port map(A => \I3.PIPEAl8r_net_1\, B => \I3.PIPEBl8r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_150\);
    
    \I2.SUB8l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_506_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l3r_net_1\);
    
    \I2.STATE3l11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_i_il12r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE3l11r_net_1\);
    
    \I2.EVNT_NUM_c9\ : AND2
      port map(A => \I2.EVNT_NUMl9r_net_1\, B => 
        \I2.EVNT_NUM_c8_net_1\, Y => \I2.EVNT_NUM_c9_net_1\);
    
    \I3.un224_reg_ads_0_a2_3_a2_2\ : AND2
      port map(A => \I3.N_544\, B => \I3.N_545_adt_net_165682_\, 
        Y => \I3.N_545\);
    
    \I3.PIPEA1_12l27r\ : AND2
      port map(A => DPR_cl27r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854488__net_1\, Y => 
        \I3.PIPEA1_12l27r_net_1\);
    
    \I5.REG_1_37\ : MUX2L
      port map(A => \I5.TEMPDATAl4r_net_1\, B => REGl424r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_37_net_1\);
    
    \I3.REG_1_i_s_i_il4r\ : OR2
      port map(A => \I3.N_203_adt_net_24459_\, B => 
        \I3.N_203_adt_net_24461_\, Y => \I3.N_203\);
    
    \I2.RAMAD1_12l4r\ : MUX2L
      port map(A => \I2.TDCDASl2r_net_1\, B => 
        \I2.TDCDBSl2r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855184__net_1\, Y => 
        \I2.RAMAD1_12l4r_net_1\);
    
    \I2.PIPE7_DTL27R_2779\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_72\);
    
    \I2.N_4249_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4249\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4249_Rd1__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I178_Y_2729\ : AO21
      port map(A => \I2.N305_0\, B => \I2.N308_0\, C => 
        \I2.N304_0\, Y => \I2.N479_adt_net_642225_\);
    
    \I2.LSRAM_IN_395\ : MUX2L
      port map(A => \I2.PIPE5_DTl11r_net_1\, B => 
        \I2.LSRAM_INl11r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_395_net_1\);
    
    \I2.PIPE8_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_550_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl22r_net_1\);
    
    \I3.PIPEA_8_0l29r\ : MUX2L
      port map(A => DPR_cl29r, B => \I3.PIPEA1l29r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855356__net_1\, Y => \I3.N_238\);
    
    \I2.ROFFSET_n11_tz\ : XOR2FT
      port map(A => \I2.ROFFSETl11r_net_1\, B => 
        \I2.ROFFSET_c10_net_1\, Y => \I2.ROFFSET_n11_tz_i\);
    
    \I1.PAGECNT_324\ : MUX2H
      port map(A => \I1.PAGECNTl3r_adt_net_835116_Rd1__net_1\, B
         => \I1.PAGECNT_n3\, S => 
        \I1.PAGECNTe_adt_net_854896__net_1\, Y => 
        \I1.PAGECNT_324_net_1\);
    
    \I2.ADEl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l13r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl13r);
    
    \I1.PAGECNT_320_adt_net_854868_\ : BFR
      port map(A => \I1.PAGECNT_320_net_1\, Y => 
        \I1.PAGECNT_320_adt_net_854868__net_1\);
    
    \I3.PIPEA_8_0l22r\ : MUX2L
      port map(A => DPR_cl22r, B => \I3.PIPEA1l22r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855360__net_1\, Y => \I3.N_231\);
    
    \I2.TRGARR_3_I_19\ : AND2
      port map(A => \I2.DWACT_ADD_CI_0_TMPl0r\, B => 
        \I2.TRGARRl1r_net_1\, Y => 
        \I2.DWACT_ADD_CI_0_g_array_1l0r\);
    
    \I1.REG_1_305\ : MUX2H
      port map(A => \REGl404r\, B => \I1.REG_74l404r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\, Y
         => \I1.REG_1_305_net_1\);
    
    \I2.BNCID_VECTwa14_1\ : AND2FT
      port map(A => \I2.TRGARRl0r_net_1\, B => 
        \I2.TRGARRl1r_net_1\, Y => \I2.BNCID_VECTwa14_1_net_1\);
    
    \I2.END_EVNT8\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT7_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT8_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I12_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L5R_138\, B => 
        \I2.PIPE4_DTL12R_858\, Y => \I2.N_53\);
    
    \I2.OFFSET_37_17l7r\ : MUX2L
      port map(A => \I2.N_762\, B => \I2.N_754\, S => 
        \I2.PIPE7_DTL26R_351\, Y => \I2.N_770\);
    
    \I2.un2_evnt_word_I_23\ : AND3
      port map(A => \I2.WOFFSETl3r\, B => 
        \I2.DWACT_FINC_E_0L0R_337\, C => \I2.WOFFSETl4r\, Y => 
        \I2.N_39\);
    
    \I4.bcntl3r\ : DFFC
      port map(CLK => CLK_c, D => \I4.bcnt_8_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I4.bcntl3r_net_1\);
    
    \I3.REG_1l87r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_268_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl87r);
    
    \I2.un1_STATE3_8_0\ : OR2
      port map(A => \I2.STATE3_nsl12r_adt_net_24672_\, B => 
        \I2.un1_STATE3\, Y => \I2.un1_STATE3_8\);
    
    \I2.PIPE7_DTL26R_2898\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_352\);
    
    \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_1_1_net_1\, Y => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\);
    
    \I1.REG_74_0_IV_0L394R_1796\ : AND2
      port map(A => \REGl394r\, B => \I1.N_265\, Y => 
        \I1.REG_74l394r_adt_net_110698_\);
    
    \I2.LSRAM_IN_414_0_0\ : OR2
      port map(A => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, B => 
        \I2.LSRAM_INl31r_net_1\, Y => \I2.LSRAM_IN_414_0_0_net_1\);
    
    \I3.RAMAD_VMEl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_27_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl3r);
    
    \I2.OFFSET_37_10l7r\ : MUX2L
      port map(A => \I2.N_706\, B => \I2.N_698\, S => 
        \I2.PIPE7_DTL26R_350\, Y => \I2.N_714\);
    
    \I2.PIPE4_DTl12r_1249\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL12R_511\);
    
    \I2.CRC32_12_0_0_m2l28r\ : MUX2L
      port map(A => \I2.DT_TEMPl28r_net_1\, B => 
        \I2.DT_SRAMl28r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854192__net_1\, Y => 
        \I2.N_4156_i_i\);
    
    \I3.un1_vdb_0_a3_0\ : NOR2
      port map(A => NOE16R_c, B => \I3.REGMAPl10r_net_1\, Y => 
        \I3.un1_vdb_0\);
    
    \I2.STATE1l12r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl6r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1l12r_net_1\);
    
    \I1.REG_74_0_ivl185r\ : AO21
      port map(A => \REGl185r\, B => \I1.N_57_268\, C => 
        \I1.REG_74l185r_adt_net_131871_\, Y => \I1.REG_74l185r\);
    
    \I3.REG_44_i_a2_0l86r\ : NOR2
      port map(A => VDB_inl3r, B => \I3.N_98\, Y => \I3.N_1667\);
    
    \I3.N_1645_i_i_o3\ : NAND2FT
      port map(A => \I3.REGMAPl0r_net_1\, B => 
        \I3.STATE1_IPL9R_877\, Y => \I3.N_1905\);
    
    \I0.TDC_RESi\ : DFFC
      port map(CLK => CLK_c, D => \I0.TDC_RESi_1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TDC_RES_c_c);
    
    \I2.PIPE9_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_294_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl25r_net_1\);
    
    \I2.TEMPF_adt_net_855740_\ : BFR
      port map(A => \I2.TEMPF_net_1\, Y => 
        \I2.TEMPF_adt_net_855740__net_1\);
    
    \I1.REG_74_0_ivl307r\ : AO21
      port map(A => \REGl307r\, B => \I1.N_177\, C => 
        \I1.REG_74l307r_adt_net_120266_\, Y => \I1.REG_74l307r\);
    
    \I2.PIPE1_DT_12l19r\ : MUX2L
      port map(A => \I2.TDCDASl19r_net_1\, B => 
        \I2.TDCDASl17r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092__net_1\, Y
         => \I2.PIPE1_DT_12l19r_net_1\);
    
    DTO_padl11r : IOB33PH
      port map(PAD => DTO(11), A => \I2.DTO_1l11r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl11r);
    
    \I2.SUB8l10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_513_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l10r_net_1\);
    
    \I2.PIPE4_DTL9R_3082\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL9R_846\);
    
    \I5.sstate2se_4\ : AO21
      port map(A => \I5.N_464\, B => \I5.sstate2l4r_net_1\, C => 
        \I5.sstate2_5_sqmuxa\, Y => \I5.sstate2_ns_el0r\);
    
    \I2.OFFSET_37_24l6r\ : MUX2L
      port map(A => \I2.N_817\, B => \I2.N_809\, S => 
        \I2.PIPE7_DTL26R_357\, Y => \I2.N_825\);
    
    \I2.FIDl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_438\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl22r);
    
    \I1.BYTECNT_307\ : MUX2H
      port map(A => \I1.BYTECNTl7r_net_1\, B => \I1.N_79\, S => 
        \I1.N_1383_225\, Y => \I1.BYTECNT_307_net_1\);
    
    \I2.STATE2_NS_0L1R_1051\ : AND2
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.N_4282\, Y => 
        \I2.STATE2_nsl1r_adt_net_24963_\);
    
    \I1.REG_74L220R_2012\ : OR2FT
      port map(A => \I1.N_347_adt_net_854788__net_1\, B => 
        \I1.N_12233_I_166\, Y => \I1.N_89_adt_net_128733_\);
    
    \I4.STATE1_tr5\ : OR2FT
      port map(A => \I4.STATE1l1r_net_1\, B => \I4.N_48_3\, Y => 
        \I4.FLUSH_1_sqmuxa\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_o2\ : OAI21TTF
      port map(A => \I2.N_72_0_107\, B => 
        \I2.N_108_0_adt_net_55153_\, C => 
        \I2.N_107_0_adt_net_320362_\, Y => 
        \I2.N_45_1_adt_net_271427_\);
    
    \I2.BNC_IDl5r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_24_0\, CLR => 
        \I2.N_4625_i_0\, SET => \I2.N_4611_i_0\, Q => 
        \I2.BNC_IDl5r_net_1\);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854656_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854656__net_1\);
    
    \I2.MIC_ERR_REGS_354\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl26r_net_1\, B => 
        \I2.MIC_ERR_REGSl25r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_354_net_1\);
    
    TDCDA_padl19r : IB33
      port map(PAD => TDCDA(19), Y => TDCDA_cl19r);
    
    \I2.ADO_3l14r\ : MUX2H
      port map(A => \I2.RPAGEl14r\, B => \I2.WPAGEl14r_net_1\, S
         => NOESRAME_c, Y => \I2.ADO_3l14r_net_1\);
    
    \I2.DT_SRAM_il27r\ : OAI21TTF
      port map(A => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, B => 
        \I2.PIPE2_DTl27r_net_1\, C => \I2.N_4647_adt_net_29104_\, 
        Y => \I2.N_4647\);
    
    \I3.PIPEA_8_0l5r\ : MUX2L
      port map(A => DPR_cl5r, B => \I3.PIPEA1l5r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855364__net_1\, Y => \I3.N_214\);
    
    \I3.REG3_0_sqmuxa_adt_net_855624_\ : BFR
      port map(A => \I3.REG3_0_sqmuxa\, Y => 
        \I3.REG3_0_sqmuxa_adt_net_855624__net_1\);
    
    \I2.DTE_21_1_IV_0_0L4R_1332\ : AND2
      port map(A => \I2.DTE_1l4r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\, Y => 
        \I2.DTE_21_1l4r_adt_net_39201_\);
    
    \I2.N_2864_0_adt_net_854268_\ : BFR
      port map(A => \I2.N_2864_0\, Y => 
        \I2.N_2864_0_adt_net_854268__net_1\);
    
    \I2.PIPE1_DT_42_1_IVL2R_1508\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl18r_net_1\, Y => 
        \I2.PIPE1_DT_42l2r_adt_net_51819_\);
    
    \I3.TCNTlde_0_o2_0\ : NOR2
      port map(A => \I3.REGMAPL13R_726\, B => \I3.REGMAPL51R_723\, 
        Y => \I3.N_1641\);
    
    \I3.REG_0_sqmuxa_2_adt_net_855296_\ : BFR
      port map(A => \I3.REG_0_sqmuxa_2\, Y => 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\);
    
    \I2.MIC_REG1l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_301_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1l0r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L6R_2382\ : OR3
      port map(A => \I3.VDBoffb_30l6r_adt_net_161985_\, B => 
        \I3.VDBoffb_30l6r_adt_net_161979_\, C => 
        \I3.VDBoffb_30l6r_adt_net_161980_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161989_\);
    
    \I2.L2TYPE_603\ : MUX2L
      port map(A => \I2.L2TYPEl14r_net_1\, B => \I2.N_4438\, S
         => \I2.N_4482_0\, Y => \I2.L2TYPE_603_net_1\);
    
    \I2.STATE1_ns_i_a2l8r\ : NAND2FT
      port map(A => \I2.END_CHAINA1_1_sqmuxa_3\, B => 
        \I2.un1_STATE1_23_net_1\, Y => \I2.N_3344_i\);
    
    \I2.BNCID_VECT_tile_0_DOUTl0r\ : MUX2L
      port map(A => \I2.DIN_REG1l0r\, B => \I2.DOUT_TMPl0r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl8r\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_682\ : AO21
      port map(A => 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855220__net_1\, B
         => 
        \I2.DTE_0_sqmuxa_i_o2_m6_i_a5_2_i_adt_net_2404__net_1\, C
         => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__182\, 
        Y => \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_60\);
    
    \I3.REGMAPl1r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un10_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl1r_net_1\);
    
    \I2.EVNT_NUM_n9\ : NOR2
      port map(A => EV_RES_c, B => \I2.EVNT_NUM_n9_tz_i\, Y => 
        \I2.EVNT_NUM_n9_net_1\);
    
    \I2.DTE_2_1l4r\ : XOR2
      port map(A => \I2.CRC32l24r_net_1\, B => 
        \I2.DTE_2_1_0l4r_net_1\, Y => \I2.DTE_2_1l4r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I14_P0N\ : OR2FT
      port map(A => \I2.N_3562_i\, B => \I2.N_3560_i_net_1\, Y
         => \I2.N268\);
    
    \I2.PIPE9_DT_295\ : MUX2L
      port map(A => \I2.PIPE9_DTl26r_net_1\, B => 
        \I2.PIPE8_DTl26r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_295_net_1\);
    
    \I1.LUT\ : DFFC
      port map(CLK => CLK_c, D => \I1.LUT_55_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.LUT_net_1\);
    
    \I2.dataout_0_adt_net_855808_\ : BFR
      port map(A => \I2.dataout_0\, Y => 
        \I2.dataout_0_adt_net_855808__net_1\);
    
    \I2.OFFSET_37_21l1r\ : MUX2L
      port map(A => \I2.N_788\, B => \I2.N_764\, S => 
        \I2.PIPE7_DTL25R_686\, Y => \I2.N_796\);
    
    \I2.NWPIPE7_1581\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE6_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE7_688\);
    
    \I1.REG_74_0_IVL322R_1894\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l322r_adt_net_118873_\);
    
    \I2.DTE_21_1_iv_0l28r\ : AO21
      port map(A => \I2.DTE_1l28r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.DTE_21_1l28r_adt_net_36759_\, Y => \I2.DTE_21_1l28r\);
    
    \I2.ROFFSETl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_907_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl11r_net_1\);
    
    \I2.WOFFSET_828\ : MUX2L
      port map(A => \I2.WOFFSETl1r_Rd1__net_1\, B => 
        \I2.N_4244_Rd1__net_1\, S => 
        \I2.N_2828_ADT_NET_1062__ADT_NET_835312_RD1__379\, Y => 
        \I2.WOFFSETl1r\);
    
    \I2.PIPE1_DT_42_1_ivl24r\ : NOR3
      port map(A => \I2.EVNT_NUM_i_m_il8r\, B => 
        \I2.PIPE1_DT_42_1_iv_1_il24r\, C => 
        \I2.PIPE1_DT_42_1_iv_0_il24r\, Y => 
        \I2.PIPE1_DT_42_1_iv_i_0l24r\);
    
    \I2.un17_tokoutas_i_a3\ : NOR2
      port map(A => \I2.TOKOUTAS_net_1\, B => \I2.TDCDRYAS_net_1\, 
        Y => \I2.N_3899\);
    
    \I3.TCNT1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT1_n5_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT1l5r_net_1\);
    
    \I2.PIPE5_DT_707\ : MUX2H
      port map(A => \I2.PIPE4_DTl31r_net_1\, B => 
        \I2.PIPE5_DTl31r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_707_net_1\);
    
    \I1.REG_74_0_IV_0L357R_1850\ : AND2
      port map(A => \FBOUTl0r\, B => \I1.REG_25_sqmuxa\, Y => 
        \I1.REG_74l357r_adt_net_115127_\);
    
    \I2.WPAGEe_adt_net_855060_\ : BFR
      port map(A => \I2.WPAGEe\, Y => 
        \I2.WPAGEe_adt_net_855060__net_1\);
    
    \I2.DTE_21_1_IV_0L10R_1300\ : AND2
      port map(A => \I2.DT_SRAMl10r_net_1\, B => 
        \I2.N_199_0_ADT_NET_1054__36\, Y => 
        \I2.DTE_21_1l10r_adt_net_38515_\);
    
    \I3.REG_1l407r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_214_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl407r);
    
    \I2.L2TYPE_4_IL12R_1621\ : AND2
      port map(A => \I2.L2TYPEl12r_net_1\, B => 
        \I2.N_4440_adt_net_67210_\, Y => 
        \I2.N_4440_adt_net_67253_\);
    
    \I3.VAS_72\ : MUX2L
      port map(A => VAD_inl10r, B => \I3.VAS_i_0_il10r\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_72_net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2531\ : AND2
      port map(A => \REGl218r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.VDBoffa_31l5r_adt_net_163656_\);
    
    \I3.VDBI_57_0_IV_0L18R_2178\ : AO21
      port map(A => \I3.VDBil18r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l18r_adt_net_139485_\, Y => 
        \I3.VDBi_57l18r_adt_net_139495_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I186_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L5R_139\, B => 
        \I2.PIPE4_DTl16r_net_1\, Y => 
        \I2.ADD_21x21_fast_I186_Y_0\);
    
    \I2.L2TYPEl7r_1556\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_596_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL7R_663\);
    
    \I1.REG_74_0_IVL379R_1820\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_27_sqmuxa_adt_net_854808__net_1\, Y => 
        \I1.REG_74l379r_adt_net_112571_\);
    
    \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852_\ : BFR
      port map(A => \I2.MIC_REG1_1_sqmuxa_0\, Y => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__2765\ : NAND3FFT
      port map(A => \I2.ENDF_838\, B => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149__net_1\, C => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_net_1\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__48\);
    
    \I2.PIPE7_DTL26R_2905\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_359\);
    
    \I2.DTE_1_869\ : MUX2L
      port map(A => \I2.DTE_1l31r_net_1\, B => \I2.DTE_21_1l31r\, 
        S => \I2.N_2868_1\, Y => \I2.DTE_1_869_net_1\);
    
    \I1.REG_74_9_i_a2l380r\ : NOR2
      port map(A => \I1.N_374\, B => \I1.N_1370\, Y => \I1.N_179\);
    
    \I3.SINGCYC_1774\ : DFFC
      port map(CLK => CLK_c, D => \I3.SINGCYC_115_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.SINGCYC_880\);
    
    \I1.N_238_Rd1__adt_net_854888_\ : BFR
      port map(A => \I1.N_238_Rd1__net_1\, Y => 
        \I1.N_238_Rd1__adt_net_854888__net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I139_Y_I_A4_2690\ : 
        AO21FTT
      port map(A => \I2.N_70_adt_net_54406__net_1\, B => 
        \I2.N525_383\, C => \I2.N_96_adt_net_481750_\, Y => 
        \I2.N_96\);
    
    \I2.PIPE10_DTl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_620_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl15r_net_1\);
    
    \I3.VDBil10r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_350_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil10r_net_1\);
    
    \I2.PIPE8_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_545_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl17r_net_1\);
    
    \I5.SDAout_12_iv_0\ : OR3
      port map(A => \I5.SDAnoe_8_adt_net_991__net_1\, B => 
        \I5.SDAout_12_adt_net_9916_\, C => 
        \I5.SDAout_12_adt_net_9915_\, Y => \I5.SDAout_12\);
    
    TOKOUTA_pad : IB33
      port map(PAD => TOKOUTA, Y => TOKOUTA_c);
    
    \I1.REG_74_0_IV_I_A2L198R_2036\ : AND2
      port map(A => \REGl198r\, B => \I1.N_182_i\, Y => 
        \I1.N_1337_adt_net_130705_\);
    
    \I2.OFFSET_37_12l1r\ : MUX2L
      port map(A => \REGl342r\, B => \I2.N_716\, S => 
        \I2.PIPE7_DTL26R_359\, Y => \I2.N_724\);
    
    \I3.PIPEA_243\ : MUX2L
      port map(A => \I3.PIPEAl12r_net_1\, B => 
        \I3.PIPEA_8l12r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854668__net_1\, Y
         => \I3.PIPEA_243_net_1\);
    
    \PULSE_0l0r_adt_net_834380_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854736__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0l0r_adt_net_834380_Rd1__net_1\);
    
    \I3.un136_reg_ads_0_a2_2_a3\ : NOR2
      port map(A => \I3.N_584\, B => \I3.N_551\, Y => 
        \I3.un136_reg_ads_0_a2_2_a3_net_1\);
    
    \I3.VDBOFFB_30_IV_0L4R_2417\ : OR2
      port map(A => \I3.VDBoffb_30l4r_adt_net_162361_\, B => 
        \I3.VDBoffb_30l4r_adt_net_162362_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162367_\);
    
    \I3.VDBi_16_m_i_o3l3r_886\ : OR2
      port map(A => \I3.REGMAPL8R_739\, B => \I3.REGMAPL9R_784\, 
        Y => \I3.N_1907_264\);
    
    \I1.REG_74L396R_1793\ : OA21FTT
      port map(A => \I1.PAGECNT_0l7r_adt_net_835112_Rd1__net_1\, 
        B => \I1.REG_74_1_396_m7_i_a5_0\, C => 
        \I1.REG_74_1_396_N_12\, Y => \I1.N_265_adt_net_110486_\);
    
    \I2.REG_1_C3_I_1743\ : OR2
      port map(A => \I2.un8_evread_1_adt_net_855780__net_1\, B
         => \I2.N_3845\, Y => \I2.N_3832_adt_net_101495_\);
    
    \I2.DTO_1l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_877_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l3r_net_1\);
    
    \I4.UN2_END_TDC_0_929\ : OR2
      port map(A => LEAD_FLAGl3r, B => LEAD_FLAGl2r, Y => 
        \I4.un2_end_tdc_0_adt_net_15179_\);
    
    \I0.TDC_RESi_1\ : AO21
      port map(A => \I0.CLEARF1_net_1\, B => \I0.CLEARF2_i\, C
         => \I0.TDC_RESi_1_adt_net_15858_\, Y => 
        \I0.TDC_RESi_1_net_1\);
    
    \I1.REG_74l404r\ : AO21FTF
      port map(A => 
        \I1.REG_74_1_396_m7_i_3_adt_net_854840__net_1\, B => 
        \I1.N_273_adt_net_109616_\, C => \I1.REG_74_13_388_N_11\, 
        Y => \I1.N_273\);
    
    \I3.un221_reg_ads_0_a2_0_a3\ : AND2FT
      port map(A => \I3.N_632\, B => 
        \I3.un221_reg_ads_0_a2_0_a3_adt_net_165933_\, Y => 
        \I3.un221_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.PIPE8_DT_16_0l8r\ : MUX2H
      port map(A => \I2.PIPE8_DTl8r_net_1\, B => 
        \I2.PIPE7_DTl8r_net_1\, S => 
        \I2.N_565_0_adt_net_855732__net_1\, Y => \I2.N_574\);
    
    \I2.N_4532_adt_net_1157_\ : AO21
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_4673\, C
         => LEAD_FLAGl3r, Y => \I2.N_4532_adt_net_1157__net_1\);
    
    \I1.REG_74_0_iv_0l368r\ : AO21
      port map(A => \REGl368r\, B => \I1.N_660\, C => 
        \I1.REG_74l368r_adt_net_113654_\, Y => \I1.REG_74l368r\);
    
    \I1.REG_1_285\ : MUX2H
      port map(A => \REGl384r\, B => \I1.REG_74l384r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y => 
        \I1.REG_1_285_net_1\);
    
    \I3.REG_1l113r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_294_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl113r);
    
    \I2.SUB9_587\ : MUX2H
      port map(A => \I2.SUB9_i_0_il19r\, B => \I2.SUB9_1l19r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_587_net_1\);
    
    \I3.TCNT_381\ : MUX2H
      port map(A => \I3.TCNTl3r_net_1\, B => \I3.TCNT_n3\, S => 
        \I3.TCNTe\, Y => \I3.TCNT_381_net_1\);
    
    \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_adt_net_803__net_1\, Y
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\);
    
    \I3.REG3_0_sqmuxa_0_a2_0_a3\ : AND2
      port map(A => \I3.REGMAPL1R_725\, B => \I3.N_1906_i_0_0\, Y
         => \I3.REG3_0_sqmuxa\);
    
    \I4.un1_FLUSH_1_sqmuxa_1\ : AND2
      port map(A => \I4.FLUSH_0_sqmuxa_net_1\, B => 
        \I4.FLUSH_1_sqmuxa\, Y => \I4.un1_FLUSH_1_sqmuxa_1_net_1\);
    
    \I1.BYTECNTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_312_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTl2r_net_1\);
    
    \I2.DTESl22r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl22r, Q => 
        \I2.DTESl22r_net_1\);
    
    \I2.G_EVNT_NUM_I_0_IL0R_2880\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_934_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUM_I_0_IL0R_312\);
    
    \I2.DTE_21_1_ivl0r\ : AOI21FTT
      port map(A => \I2.DTE_1l0r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, C => 
        \I2.DTE_21_1_iv_2_il0r\, Y => \I2.DTE_21_1_iv_i_0l0r\);
    
    \I3.VASl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_63_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl1r_net_1\);
    
    \I3.VDBI_57_IVL1R_2267\ : AO21
      port map(A => \I3.PIPEAl1r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l1r_adt_net_145935_\, Y => 
        \I3.VDBi_57l1r_adt_net_145945_\);
    
    \I2.PIPE9_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_290_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl21r_net_1\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_685\ : AO21
      port map(A => 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855220__net_1\, B
         => \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__870\, 
        C => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_adt_net_19813_\, Y
         => \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_63\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I153_Y_I_O4_1566\ : AO21
      port map(A => \I2.PIPE4_DTl15r_net_1\, B => 
        \I2.PIPE4_DTl16r_net_1\, C => \I2.RAMDT4L12R_796\, Y => 
        \I2.N_33_0_adt_net_55958_\);
    
    \I2.INT_ERRBS\ : DFFC
      port map(CLK => CLK_c, D => \I2.INT_ERRBS_527_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.INT_ERRBS_i_i\);
    
    \I2.un1_END_CHAINA1_0_sqmuxa_i_a2_1\ : OAI21TTF
      port map(A => \I2.STATE1l7r_net_1\, B => 
        \I2.END_CHAINB1_709_adt_net_2397__net_1\, C => 
        \I2.N_3347_1_adt_net_21905_\, Y => \I2.N_3347_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I109_UN1_Y_1661\ : AND2
      port map(A => \I2.N288\, B => \I2.N292\, Y => 
        \I2.I109_un1_Y_adt_net_70914_\);
    
    \I1.REG_74_0_IVL272R_1951\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, Y => 
        \I1.REG_74l272r_adt_net_123646_\);
    
    \I2.DTO_16_1_iv_0_a2_4_18_m7_0_m5\ : MUX2H
      port map(A => \I2.END_EVNT5_net_1\, B => 
        \I2.END_EVNT10_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854216__net_1\, Y => 
        \I2.DTO_16_1_iv_0_a2_4_18_N_11\);
    
    \I3.VAS_68\ : MUX2L
      port map(A => VAD_inl6r, B => \I3.VASl6r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_68_net_1\);
    
    \I2.L2SERV_n3\ : XOR2FT
      port map(A => \I2.RPAGEL15R_522\, B => \I2.L2SERV_c2_net_1\, 
        Y => \I2.L2SERV_n3_net_1\);
    
    \I2.OFFSET_37_27l7r\ : MUX2L
      port map(A => \I2.N_842\, B => \I2.N_826\, S => 
        \I2.PIPE7_DTL25R_686\, Y => \I2.N_850\);
    
    \I2.SUB9_1_ADD_18x18_fast_I156_Y\ : XOR2
      port map(A => \I2.N436\, B => \I2.ADD_18x18_fast_I156_Y_0\, 
        Y => \I2.SUB9_1l19r\);
    
    \I5.un1_AIR_PULSE_0_sqmuxa_i\ : AND2
      port map(A => REGl117r, B => \I5.N_479\, Y => \I5.N_459\);
    
    DTO_padl28r : IOB33PH
      port map(PAD => DTO(28), A => \I2.DTO_1l28r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl28r);
    
    \I3.REG_1_195\ : MUX2L
      port map(A => VDB_inl14r, B => \I3.REGl147r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\, Y => 
        \I3.REG_1_195_0\);
    
    \I2.DTO_16_1l24r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l24r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l24r_Rd1__net_1\);
    
    \I1.LUT_55_2072\ : NOR2FT
      port map(A => \I1.LUT_net_1\, B => \I1.N_56\, Y => 
        \I1.LUT_55_adt_net_133935_\);
    
    \I3.VDBi_40_sn_m2_0_752\ : NOR2
      port map(A => \I3.REGMAPL57R_539\, B => 
        \I3.REGMAP_I_0_IL58R_537\, Y => \I3.N_354_0_130\);
    
    \I3.VDBOFFA_31_IV_0L2R_2584\ : AND2
      port map(A => \REGl231r\, B => \I3.REGMAPl26r_net_1\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164222_\);
    
    \I2.OFFSET_37_20l7r\ : MUX2L
      port map(A => \I2.N_786\, B => \I2.N_778\, S => 
        \I2.PIPE7_DTL26R_355\, Y => \I2.N_794\);
    
    \I1.PAGECNTL8R_2939\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_319_adt_net_854860__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL8R_456\);
    
    \I2.OFFSET_562\ : MUX2L
      port map(A => \I2.OFFSETl2r_net_1\, B => \I2.OFFSET_37l2r\, 
        S => \I2.UN1_NWPIPE7_2_298\, Y => \I2.OFFSET_562_net_1\);
    
    FID_padl15r : OB33PH
      port map(PAD => FID(15), A => FID_cl15r);
    
    \I5.AIR_CHAIN\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_CHAIN_15_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_CHAIN_net_1\);
    
    \I4.STATE1_ns_0l2r\ : AO21FTF
      port map(A => \I4.FLUSH_0_sqmuxa_net_1\, B => 
        \I4.STATE1_nsl2r_adt_net_15265_\, C => 
        \I4.FLUSH_1_sqmuxa\, Y => \I4.STATE1_nsl2r\);
    
    \I3.VDBOFFB_30_IV_0L0R_2478\ : AND2
      port map(A => \REGl357r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        Y => \I3.VDBoffb_30l0r_adt_net_163090_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I149_Y\ : XOR2
      port map(A => \I2.N457\, B => \I2.ADD_18x18_fast_I149_Y_0\, 
        Y => \I2.SUB9_1l12r\);
    
    REGl259r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_160_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl259r\);
    
    \I5.AIR_WDATA_9l11r\ : AND2
      port map(A => \I5.sstate2l3r_net_1\, B => 
        \I5.SENS_ADDRl2r_net_1\, Y => \I5.AIR_WDATA_9l11r_net_1\);
    
    \I2.OFFSET_37_11l2r\ : MUX2L
      port map(A => \REGl375r\, B => \REGl311r\, S => 
        \I2.PIPE7_DTL27R_83\, Y => \I2.N_717\);
    
    \I3.VDBI_57_IVL3R_2258\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => 
        \I3.VDBi_55l3r_net_1\, C => 
        \I3.VDBi_57l3r_adt_net_145072_\, Y => 
        \I3.VDBi_57l3r_adt_net_145073_\);
    
    \I3.PIPEAl25r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_256_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl25r_net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__3076\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854736__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__830\);
    
    \I2.L2TYPE_4_il13r\ : OAI21TTF
      port map(A => \I2.L2AS_adt_net_855716__net_1\, B => 
        \I2.N_4439_adt_net_67071_\, C => 
        \I2.N_4439_adt_net_67114_\, Y => \I2.N_4439\);
    
    \I2.FID_7_0_IVL20R_952\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl68r, C => 
        \I2.FID_7l20r_adt_net_17380_\, Y => 
        \I2.FID_7l20r_adt_net_17388_\);
    
    \I2.PIPE5_DT_701\ : MUX2L
      port map(A => \I2.PIPE5_DTl25r_net_1\, B => 
        \I2.PIPE4_DTl25r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_701_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I178_Y_2733\ : AO21
      port map(A => \I2.N479_adt_net_538167_\, B => 
        \I2.N479_adt_net_538220_\, C => \I2.N479_adt_net_649015_\, 
        Y => \I2.N479\);
    
    \I3.VDBoff_117\ : MUX2L
      port map(A => \I3.VDBoffl1r_net_1\, B => \I3.N_2065\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_117_net_1\);
    
    \I1.REG_74_0_ivl184r\ : AO21
      port map(A => \REGl184r\, B => \I1.N_57_269\, C => 
        \I1.REG_74l184r_adt_net_131957_\, Y => \I1.REG_74l184r\);
    
    \I2.SUB8_519\ : MUX2H
      port map(A => \I2.N_3558_i_adt_net_855584__net_1\, B => 
        \I2.SUB8_2_i_i_0l16r\, S => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855140__net_1\, Y => 
        \I2.SUB8_519_net_1\);
    
    DPR_padl8r : IB33
      port map(PAD => DPR(8), Y => DPR_cl8r);
    
    \I3.un15_anycyc\ : OR2
      port map(A => \I3.un15_anycyc_adt_net_147611_\, B => 
        \I3.un15_anycyc_adt_net_147613_\, Y => 
        \I3.un15_anycyc_net_1\);
    
    \I2.G_EVNT_NUM_N9_0_1055\ : XOR2
      port map(A => \I2.N_207\, B => \I2.G_EVNT_NUMl9r_net_1\, Y
         => \I2.G_EVNT_NUM_n9_adt_net_26657_\);
    
    STBMIC_pad : OB33PH
      port map(PAD => STBMIC, A => STBMIC_c);
    
    \I3.un131_reg_ads_0_a2_1_a3\ : NOR2
      port map(A => \I3.N_586\, B => \I3.N_551\, Y => 
        \I3.un131_reg_ads_0_a2_1_a3_net_1\);
    
    \I2.N_182_ADT_NET_1007__2822\ : OR2
      port map(A => \I2.STATE2L0R_588\, B => 
        \I2.STATE2_nsl2r_adt_net_24911_\, Y => 
        \I2.N_182_ADT_NET_1007__155\);
    
    \I5.AIR_WDATA_55\ : MUX2H
      port map(A => \I5.N_480\, B => \I5.AIR_WDATAl0r_net_1\, S
         => \I5.N_461\, Y => \I5.AIR_WDATA_55_net_1\);
    
    \I3.REG_1_213\ : MUX2L
      port map(A => VDB_inl0r, B => REGl406r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_213_0\);
    
    \I2.FIDl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_440\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl24r);
    
    VDB_padl17r : IOB33PH
      port map(PAD => VDB(17), A => \I3.VDBml17r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl17r);
    
    \I2.un1_ERR_WORDS_RDY_0_sqmuxa_0_0_a5\ : AND2
      port map(A => \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23154_\, 
        B => \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23155_\, Y => 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1\);
    
    \I2.L2TYPE_4_IL5R_1633\ : AND2
      port map(A => \I2.L2TYPE_i_0_il5r\, B => 
        \I2.N_4447_adt_net_68073_\, Y => 
        \I2.N_4447_adt_net_68116_\);
    
    \I2.L2TYPE_4_IL14R_1617\ : AND2
      port map(A => \I2.L2TYPEl14r_net_1\, B => 
        \I2.N_4438_adt_net_66932_\, Y => 
        \I2.N_4438_adt_net_66975_\);
    
    \I2.REG_1_n8_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855788__net_1\, B
         => REGl40r, Y => \I2.REG_1_n8_0_net_1\);
    
    \I3.VDBI_57_IVL1R_2266\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854360__net_1\, B
         => \I3.VDBoffl1r_net_1\, Y => 
        \I3.VDBi_57l1r_adt_net_145935_\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854616_\ : BFR
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620__net_1\, 
        Y => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854616__net_1\);
    
    \I4.STATE1_NS_0L2R_931\ : NOR2
      port map(A => \I4.un2_end_tdc_0_net_1\, B => 
        \I4.un2_end_tdc_1_net_1\, Y => 
        \I4.STATE1_nsl2r_adt_net_15265_\);
    
    \I2.TDCDASl21r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl21r, Q => 
        \I2.TDCDASl21r_net_1\);
    
    \I1.LUT_0_sqmuxa_i_0_a2\ : NOR3FTT
      port map(A => \I1.sstate_nsl4r\, B => \I1.N_317_Ra1_\, C
         => \I1.N_333_Ra1_\, Y => \I1.N_606_Ra1_\);
    
    \I3.TCNTlde_0_a2_1_i_o3\ : NAND2
      port map(A => \I3.SINGCYC_334\, B => \I3.STATE1_IPL9R_877\, 
        Y => \I3.N_276\);
    
    \I2.PIPE4_DTL4R_2961\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL4R_478\);
    
    \I1.REG_74_0_iv_0_0l248r\ : AO21
      port map(A => \REGl248r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l248r_adt_net_125949_\, Y => \I1.REG_74l248r\);
    
    \I5.SCL_1_i\ : MUX2L
      port map(A => \I5.SCL_net_1\, B => 
        \I5.SCL_1_i_a2_0_1_net_1\, S => \I5.N_82\, Y => 
        \I5.N_484\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_a2_4\ : AND2
      port map(A => \I2.RAMDT4L12R_822\, B => 
        \I2.N_140_0_adt_net_947__net_1\, Y => \I2.N_140_0\);
    
    \I3.REGMAPL20R_3026\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un81_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL20R_780\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I138_Y_0_0\ : AO21FTT
      port map(A => \I2.N_74_104\, B => 
        \I2.ADD_21x21_fast_I138_Y_0_0_0_adt_net_58684_\, C => 
        \I2.N_112_1\, Y => \I2.ADD_21x21_fast_I138_Y_0_0_0\);
    
    VAD_padl28r : IOB33PH
      port map(PAD => VAD(28), A => \I3.VADml28r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl28r);
    
    \I1.REG_74_1_I_A2_A0L404R_1814\ : OR2
      port map(A => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__198\, 
        B => \I1.N_237\, Y => \I1.N_1367_i_adt_net_112072_\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l6r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl6r_net_1\, Q => 
        \I2.DIN_REG1l6r\);
    
    \I2.PIPE1_DT_749\ : MUX2L
      port map(A => \I2.PIPE1_DTl22r_net_1\, B => 
        \I2.PIPE1_DT_42l22r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854568__net_1\, 
        Y => \I2.PIPE1_DT_749_net_1\);
    
    \I1.REG_0_sqmuxa_i_0_a2_645_944\ : AND3
      port map(A => \I1.SSTATEL0R_307\, B => \I1.N_324_25\, C => 
        \I1.BITCNTL2R_753\, Y => \I1.N_598_322\);
    
    \I2.PIPE8_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_544_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl16r_net_1\);
    
    \I2.SUB8l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_505_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l2r_net_1\);
    
    REGl351r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_252_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl351r\);
    
    \I3.un6_asb_0_0_x2\ : XOR2FT
      port map(A => VAD_inl28r, B => GA_cl0r, Y => \I3.N_260_i_0\);
    
    \I2.DTO_16_1_IV_0L4R_1200\ : AO21
      port map(A => \I2.N_457\, B => \I2.DTE_2_1l4r_net_1\, C => 
        \I2.DTO_16_1l4r_adt_net_34376_\, Y => 
        \I2.DTO_16_1l4r_adt_net_34385_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I138_Y_0_A2_1580\ : AND3
      port map(A => \I2.N357_0\, B => \I2.N_53_0\, C => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_i_1\, Y => 
        \I2.N_100_0_adt_net_58633_\);
    
    \I2.LSRAM_WR\ : DFFS
      port map(CLK => CLK_c, D => \I2.LSRAM_WR_380_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_WR_net_1\);
    
    \I2.PIPE6_DT_474\ : MUX2H
      port map(A => \I2.PIPE5_DTl20r_net_1\, B => 
        \I2.PIPE6_DTl20r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_474_net_1\);
    
    \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__2839\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__197\);
    
    \I4.un1_lead_flag_1_6_0\ : MUX2L
      port map(A => \I4.N_5\, B => \I4.N_4\, S => 
        \I4.bcntl1r_net_1\, Y => \I4.N_6\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_684\ : AO21
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__26\, B => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__871\, C
         => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_adt_net_19813_\, Y
         => \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_62\);
    
    \I2.CRC32_12_i_0_x2l27r\ : XOR2FT
      port map(A => \I2.CRC32l27r_net_1\, B => \I2.N_230_i_i\, Y
         => \I2.N_246_i_i_0\);
    
    \I2.PIPE10_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_618_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl13r_net_1\);
    
    \I1.N_1169_adt_net_854828_\ : BFR
      port map(A => \I1.N_1169\, Y => 
        \I1.N_1169_adt_net_854828__net_1\);
    
    \I2.DTE_21_1_iv_2l0r\ : AO21
      port map(A => \I2.STATE2L3R_440\, B => \I2.DTO_9_ivl0r\, C
         => \I2.DTE_21_1_iv_2_il0r_adt_net_39733_\, Y => 
        \I2.DTE_21_1_iv_2_il0r\);
    
    \I5.TEMPDATAl5r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_79_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl5r_net_1\);
    
    \I3.NOEDTKi_636\ : DFFS
      port map(CLK => CLK_c, D => \I3.NOEDTKi_111_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => NOEDTK_C_14);
    
    \I2.ROFFSET_912\ : MUX2H
      port map(A => \I2.ROFFSETl6r_net_1\, B => 
        \I2.ROFFSET_n6_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_912_net_1\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854428_\ : BFR
      port map(A => \I2.N_4667_1_adt_net_1046__net_1\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854428__net_1\);
    
    \I3.PIPEA_8_0l1r\ : MUX2L
      port map(A => DPR_cl1r, B => \I3.PIPEA1l1r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855364__net_1\, Y => \I3.N_210\);
    
    \I2.CRC32_12_il25r\ : NOR2
      port map(A => \I2.N_2867_1_adt_net_854964__net_1\, B => 
        \I2.N_42_i_0_i_0\, Y => \I2.N_3942\);
    
    \I2.OFFSET_37_15l3r\ : MUX2L
      port map(A => \REGl232r\, B => \REGl168r\, S => 
        \I2.PIPE7_DTL27R_71\, Y => \I2.N_750\);
    
    \I3.PIPEA1_12l30r\ : NAND2FT
      port map(A => DPR_cl30r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, Y => 
        \I3.PIPEA1_12l30r_net_1\);
    
    \I2.DTE_21_1_IV_0L13R_1283\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855116__net_1\, B => 
        \I2.EVNT_WORDl9r_net_1\, Y => 
        \I2.DTE_21_1l13r_adt_net_38165_\);
    
    \I3.REG_1l142r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_190_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl142r\);
    
    \I2.PIPE6_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_477_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl23r_net_1\);
    
    \I1.PAGECNTe_adt_net_854900_\ : BFR
      port map(A => \I1.PAGECNTe\, Y => 
        \I1.PAGECNTe_adt_net_854900__net_1\);
    
    \I1.BITCNT_n2_i_i_x2\ : XOR2
      port map(A => \I1.N_324\, B => \I1.BITCNTl2r_net_1\, Y => 
        \I1.N_389_i_i_0\);
    
    \I2.MIC_ERR_REGSl32r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_361_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl32r_net_1\);
    
    \I3.REG_1l146r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_194_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl146r\);
    
    \I2.TRGSERVL0R_2949\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.DWACT_ADD_CI_0_partial_sum_1l0r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGSERVL0R_466\);
    
    \I3.VDBOFFA_31_IV_0L4R_2558\ : AO21
      port map(A => \REGl265r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        C => \I3.VDBoffa_31l4r_adt_net_163854_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163883_\);
    
    \I1.LUT_0_sqmuxa_i_0_o2_i_0_834_1236\ : NOR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__186\, B
         => \I1.N_325_501\, Y => \I1.N_328_I_0_498\);
    
    \I3.PULSE_337\ : MUX2L
      port map(A => PULSEl7r, B => \I3.N_1897\, S => 
        \I3.N_1409_adt_net_854740__net_1\, Y => 
        \I3.PULSE_337_net_1\);
    
    MYBERR_pad : OB33PH
      port map(PAD => MYBERR, A => MYBERR_c);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I138_Y_0_A2_2_2665\ : 
        NOR3FFT
      port map(A => \I2.N_128\, B => \I2.N_114_adt_net_275711_\, 
        C => \I2.N_70_adt_net_255802__net_1\, Y => 
        \I2.N_114_adt_net_275800_\);
    
    \I2.ADOl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l13r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl13r);
    
    \I1.REG_15_sqmuxa_0_a2\ : OR2
      port map(A => 
        \I1.REG_15_sqmuxa_adt_net_1457__adt_net_854380__net_1\, B
         => \I1.N_254_276\, Y => \I1.REG_15_sqmuxa\);
    
    \I2.OFFSET_37_22l1r\ : MUX2L
      port map(A => \REGl238r\, B => \REGl174r\, S => 
        \I2.PIPE7_DTL27R_85\, Y => \I2.N_804\);
    
    \I2.EVNT_WORD_718\ : MUX2H
      port map(A => \I2.EVNT_WORDl5r_net_1\, B => \I2.I_24\, S
         => \I2.N_2864_0_adt_net_854276__net_1\, Y => 
        \I2.EVNT_WORD_718_net_1\);
    
    \I1.REG_74_0_ivl293r\ : AO21
      port map(A => \REGl293r\, B => \I1.N_169\, C => 
        \I1.REG_74l293r_adt_net_121470_\, Y => \I1.REG_74l293r\);
    
    \I1.PAGECNTLDE_0_O4_1757\ : NOR2FT
      port map(A => \I1.SSTATEL10R_380\, B => \I1.N_349_RD1__486\, 
        Y => \I1.N_370_adt_net_106310_\);
    
    \I2.BNCID_VECTror_adt_net_48230_\ : AO21
      port map(A => \I2.BNCID_VECTra15_1_net_1\, B => 
        \I2.BNCID_VECTro_3\, C => 
        \I2.BNCID_VECTror_adt_net_48219__net_1\, Y => 
        \I2.BNCID_VECTror_adt_net_48230__net_1\);
    
    \I2.PIPE9_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_269_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl0r_net_1\);
    
    \I1.REG_74_0_IV_0L275R_1948\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, Y => 
        \I1.REG_74l275r_adt_net_123388_\);
    
    \I5.COMMAND_45\ : MUX2H
      port map(A => \I5.COMMANDl8r_net_1\, B => 
        \I5.COMMAND_4l8r_net_1\, S => \I5.SSTATE1L13R_4\, Y => 
        \I5.COMMAND_45_net_1\);
    
    \I3.PIPEA1_12l11r\ : AND2
      port map(A => DPR_cl11r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854504__net_1\, Y => 
        \I3.PIPEA1_12l11r_net_1\);
    
    \I2.SUB8_522_2738\ : OR3
      port map(A => \I2.SUB8_522_adt_net_659164_\, B => 
        \I2.SUB8_522_adt_net_659169_\, C => 
        \I2.SUB8_522_adt_net_659160_\, Y => \I2.SUB8_522_net_1\);
    
    \I2.MIC_ERR_REGS_330\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl2r_net_1\, B => 
        \I2.MIC_ERR_REGSl1r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_330_net_1\);
    
    \I1.UN1_SBYTE13_I_I_I_1_1772\ : MUX2L
      port map(A => PULSEl6r, B => \I1.N_349_Rd1__net_1\, S => 
        \I1.sstatel3r_net_1\, Y => 
        \I1.un1_sbyte13_i_i_i_1_adt_net_108180_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I66_Y_1682\ : AND2FT
      port map(A => \I2.LSRAM_OUTl6r\, B => 
        \I2.PIPE7_DTl6r_net_1\, Y => \I2.N316_i_i_adt_net_86582_\);
    
    REGl350r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_251_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl350r\);
    
    \I2.DTO_1l18r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l18r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l18r_Rd1__net_1\);
    
    \I3.TCNT_n2_0_0_o2\ : OR2
      port map(A => \I3.TCNTL0R_428\, B => \I3.TCNTL1R_429\, Y
         => \I3.N_1911\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_o2\ : NAND3
      port map(A => \I2.N_128\, B => \I2.N_95\, C => \I2.N_108\, 
        Y => \I2.N_45_0\);
    
    \I2.EVNT_WORDl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_718_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl5r_net_1\);
    
    \I2.SRAM_EVNT_c2_i\ : OAI21TTF
      port map(A => \I2.SRAM_EVNTl2r_net_1\, B => \I2.N_135\, C
         => \I2.N_3827_adt_net_101792_\, Y => \I2.N_3827\);
    
    \I3.un106_reg_ads_0_a2_0_a2_0_989\ : NOR2FT
      port map(A => \I3.VASl12r_net_1\, B => \I3.N_547_371\, Y
         => \I3.N_548_367\);
    
    NWRSRAM_TST_pad : OB33PH
      port map(PAD => NWRSRAM_TST, A => NWRSRAM_TST_c);
    
    \I2.CHA_DATA8_2_i\ : OAI21FTF
      port map(A => \I2.CHA_DATA8_net_1\, B => \I2.N_4403\, C => 
        \I2.N_4398_adt_net_90118_\, Y => \I2.N_4398\);
    
    \I1.PAGECNT_n0_0_0\ : OAI21
      port map(A => \I1.PAGECNTl0r_adt_net_833884_Rd1__net_1\, B
         => \I1.un1_sbyte13_1_i_1\, C => \I1.N_473_204\, Y => 
        \I1.PAGECNT_n0\);
    
    \I2.SUB9l8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_576_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l8r_net_1\);
    
    \I2.STATE4_ns_il2r\ : AOI21FTT
      port map(A => \I2.STATE4l2r_net_1\, B => \I2.N_3376_1\, C
         => \I2.STATE4l1r_net_1\, Y => \I2.STATE4_ns_il2r_net_1\);
    
    \I2.DTO_1_900\ : MUX2L
      port map(A => \I2.DTO_1l26r_Rd1__net_1\, B => 
        \I2.DTO_16_1l26r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834756_Rd1__net_1\, Y
         => \I2.DTO_1l26r\);
    
    \I1.REG_1_170\ : MUX2H
      port map(A => \REGl269r\, B => \I1.REG_74l269r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y => 
        \I1.REG_1_170_net_1\);
    
    \I3.REG3l4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_129_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l4r_net_1\);
    
    \I0.EV_RESi_1460\ : DFFC
      port map(CLK => CLK_c, D => \I0.EV_RESi_1_net_1\, CLR => 
        \I0.un4_hwresi_i\, Q => EV_RES_C_567);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I179_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_800\, B => 
        \I2.PIPE4_DTl9r_net_1\, Y => 
        \I2.ADD_21x21_fast_I179_Y_0_0\);
    
    \I1.REG_5_sqmuxa_adt_net_854704_\ : BFR
      port map(A => \I1.REG_5_sqmuxa\, Y => 
        \I1.REG_5_sqmuxa_adt_net_854704__net_1\);
    
    \I2.DT_SRAM_i_ml30r\ : NOR2
      port map(A => \I2.CRC32_1_SQMUXA_0_38\, B => 
        \I2.DT_SRAMl30r_net_1\, Y => \I2.DT_SRAM_i_ml30r_net_1\);
    
    \I3.N_127_adt_net_855312_\ : BFR
      port map(A => \I3.N_127\, Y => 
        \I3.N_127_adt_net_855312__net_1\);
    
    \I2.FID_7_0_IVL14R_964\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl62r, C => 
        \I2.FID_7l14r_adt_net_17987_\, Y => 
        \I2.FID_7l14r_adt_net_17995_\);
    
    VDB_padl12r : IOB33PH
      port map(PAD => VDB(12), A => \I3.VDBml12r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl12r);
    
    \I3.VDBi_40l3r\ : MUX2L
      port map(A => \I3.N_341\, B => \I3.N_135\, S => 
        \I3.N_354_0_adt_net_855368__net_1\, Y => 
        \I3.VDBi_40l3r_net_1\);
    
    \I3.VDBi_365\ : MUX2L
      port map(A => \I3.VDBil25r_net_1\, B => \I3.VDBi_57l25r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_365_net_1\);
    
    \I3.VDBi_359\ : MUX2L
      port map(A => \I3.VDBil19r_net_1\, B => \I3.VDBi_57l19r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_359_net_1\);
    
    VAD_padl9r : IOB33PH
      port map(PAD => VAD(9), A => \I3.VADml9r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl9r);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I136_Y_0_o2\ : AO21
      port map(A => \I2.N_92\, B => \I2.N_147_0_adt_net_604832_\, 
        C => \I2.N_163_adt_net_1241__net_1\, Y => \I2.N507\);
    
    \I3.un76_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_585\, B => \I3.N_553\, Y => 
        \I3.un76_reg_ads_0_a2_0_a3_net_1\);
    
    \I4.un2_end_tdc_0\ : OR3
      port map(A => LEAD_FLAGl1r, B => LEAD_FLAGl0r, C => 
        \I4.un2_end_tdc_0_adt_net_15179_\, Y => 
        \I4.un2_end_tdc_0_net_1\);
    
    \I2.DTO_16_1l23r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l23r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l23r_Rd1__net_1\);
    
    \I2.CRC32_12_i_0l11r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_248_i_i_0\, Y => 
        \I2.N_3928\);
    
    \I2.ROFFSET_c10\ : AND2
      port map(A => \I2.ROFFSETl10r_net_1\, B => 
        \I2.ROFFSET_c9_net_1\, Y => \I2.ROFFSET_c10_net_1\);
    
    \I5.REG_1_32\ : MUX2L
      port map(A => REGl132r, B => REGl419r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_32_net_1\);
    
    \I2.DTE_21_1_iv_0l6r\ : OR3
      port map(A => \I2.DTE_21_1l6r_adt_net_38973_\, B => 
        \I2.DTE_21_1l6r_adt_net_38981_\, C => 
        \I2.DTE_21_1l6r_adt_net_38982_\, Y => \I2.DTE_21_1l6r\);
    
    \I2.BNCID_VECT_tile_0_DIN_REG1l0r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl8r_net_1\, Q => 
        \I2.DIN_REG1l0r\);
    
    VDB_padl16r : IOB33PH
      port map(PAD => VDB(16), A => \I3.VDBml16r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl16r);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I153_Y_i_o4\ : AND3
      port map(A => \I2.N_33_0_adt_net_55958_\, B => \I2.N_57_0\, 
        C => \I2.N_33_0_adt_net_55957_\, Y => \I2.N_33_0\);
    
    \I2.TRGSERVL1R_2951\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l1r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVL1R_468\);
    
    \I2.FIDl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_426\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl10r);
    
    VAD_padl3r : IOB33PH
      port map(PAD => VAD(3), A => \I3.VADml3r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl3r);
    
    \I1.REG_74l292r\ : OR2FT
      port map(A => \I1.REG_15_sqmuxa\, B => 
        \I1.N_161_adt_net_1449__net_1\, Y => \I1.N_161\);
    
    \I3.VADm_0_a3l19r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl19r_net_1\, Y => \I3.VADml19r\);
    
    \I5.BITCNT_86\ : MUX2H
      port map(A => \I5.BITCNT_c0\, B => \I5.N_50\, S => 
        \I5.BITCNTe\, Y => \I5.BITCNT_86_net_1\);
    
    \I3.REGMAPl17r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un68_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPl17r_net_1\);
    
    \I2.PIPE6_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_485_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl31r_net_1\);
    
    \I3.STATE1_TR24_I_0_O2_1_0_2109\ : NOR2
      port map(A => \I3.REGMAPl33r_net_1\, B => 
        \I3.REGMAPl51r_net_1\, Y => 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135383_\);
    
    TDCDA_padl1r : IB33
      port map(PAD => TDCDA(1), Y => TDCDA_cl1r);
    
    \I2.OFFSET_37_21l2r\ : MUX2L
      port map(A => \I2.N_789\, B => \I2.N_765\, S => 
        \I2.PIPE7_DTL25R_685\, Y => \I2.N_797\);
    
    \I2.PIPE7_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl11r_net_1\);
    
    \I2.un28_sram_empty_8_0\ : MUX2L
      port map(A => \I2.L2TYPE_I_0_IL9R_658\, B => 
        \I2.L2TYPE_I_0_IL1R_657\, S => \I2.RPAGEL15R_517\, Y => 
        \I2.N_627\);
    
    \I2.BNCID_VECTrff_0\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_0_265_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_0\);
    
    \I1.PAGECNT_322\ : MUX2H
      port map(A => \I1.PAGECNTl5r_adt_net_855548__net_1\, B => 
        \I1.PAGECNT_n5\, S => \I1.PAGECNTe_adt_net_854896__net_1\, 
        Y => \I1.PAGECNT_322_net_1\);
    
    \I2.PIPE7_DTL26R_2904\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_358\);
    
    \I3.PIPEA1l11r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_309_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l11r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I57_Y_0_O2_1560\ : OA21TTF
      port map(A => \I2.RAMDT4L8R_527\, B => 
        \I2.PIPE4_DT_I_IL1R_473\, C => \I2.N_85_0\, Y => 
        \I2.N357_0_adt_net_55523_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I180_UN1_Y_2661\ : AO21
      port map(A => \I2.I180_un1_Y_adt_net_240062_\, B => 
        \I2.I180_un1_Y_adt_net_240115_\, C => 
        \I2.I180_un1_Y_adt_net_252355_\, Y => \I2.I180_un1_Y\);
    
    \I2.RAMDT4L12R_3068\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_822\);
    
    \I1.UN1_SBYTE13_1_I_0_S_1759\ : AO21FTT
      port map(A => \I1.SSTATEL10R_759\, B => 
        \I1.N_606_Rd1__net_1\, C => \I1.N_328_I_0_211\, Y => 
        \I1.un1_sbyte13_1_i_1_adt_net_106369_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I190_Y\ : XOR2FT
      port map(A => \I2.N_1_1\, B => \I2.ADD_21x21_fast_I190_Y_0\, 
        Y => \I2.un27_pipe5_dt0l20r\);
    
    \I2.DTE_21_1_ivl3r\ : AOI21FTT
      port map(A => \I2.DTE_1l3r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, C => 
        \I2.DTE_21_1_iv_2_il3r\, Y => \I2.DTE_21_1_iv_i_0l3r\);
    
    \I5.SENS_ADDRl2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SENS_ADDR_6l2r_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.SENS_ADDRl2r_net_1\);
    
    \I2.un21_sram_empty_1\ : XOR2
      port map(A => \I2.RPAGEL13R_610\, B => \I2.L2ARRL1R_603\, Y
         => \I2.un21_sram_empty_1_net_1\);
    
    \I2.STATE2_ns_4_0l2r\ : OR3
      port map(A => \I2.STATE2_nsl2r_adt_net_24907_\, B => 
        \I2.STATE2_nsl2r_adt_net_24911_\, C => 
        \I2.STATE2_nsl2r_adt_net_24916_\, Y => \I2.STATE2_nsl2r\);
    
    \I2.PIPE6_DT_475\ : MUX2H
      port map(A => \I2.PIPE5_DTl21r_net_1\, B => 
        \I2.PIPE6_DTl21r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_475_net_1\);
    
    \I2.L2TYPE_598\ : MUX2L
      port map(A => \I2.L2TYPE_i_0_il9r\, B => \I2.N_4443\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_598_net_1\);
    
    \I3.REG_44_IL87R_2304\ : AOI21FTT
      port map(A => REGl87r, B => \I3.N_98_0\, C => \I3.N_1669\, 
        Y => \I3.N_1633_adt_net_150293_\);
    
    N_1_I3_TCNT3_372 : MUX2H
      port map(A => \I3.TCNT3l7r_net_1\, B => \N_1.I3.TCNT3_n7\, 
        S => \TICKl1r\, Y => TCNT3_372);
    
    \I2.un8_evread_1_adt_net_855796_\ : BFR
      port map(A => \I2.un8_evread_1\, Y => 
        \I2.un8_evread_1_adt_net_855796__net_1\);
    
    \I2.TOKOUTAS_3_i\ : MUX2H
      port map(A => TOKOUTA_BP_c, B => TOKOUTA_c, S => 
        \I2.N_4424\, Y => \I2.TOKOUTAS_3_i_net_1\);
    
    \I1.REG_74l220r_786\ : OR3
      port map(A => \I1.N_89_adt_net_128732_\, B => 
        \I1.N_97_6_adt_net_854712__net_1\, C => 
        \I1.N_89_adt_net_128736_\, Y => \I1.N_89_164\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__2821\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__149\);
    
    \I3.RAMAD_VME_39\ : MUX2H
      port map(A => RAMAD_VMEl15r, B => \I3.REGl98r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_39_net_1\);
    
    \I2.OFFSET_37_18l2r\ : MUX2L
      port map(A => \REGl247r\, B => \REGl183r\, S => 
        \I2.PIPE7_DTL27R_83\, Y => \I2.N_773\);
    
    \I2.L2TYPEl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_601_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl12r_net_1\);
    
    \I3.REG_1l76r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_177_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl76r);
    
    \I3.EVREAD_DS_1622\ : DFFC
      port map(CLK => CLK_c, D => \I3.EVREAD_DS_124_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I3.EVREAD_DS_729\);
    
    \I2.un28_sram_empty_4_0\ : MUX2L
      port map(A => \I2.L2TYPEL10R_654\, B => \I2.L2TYPEL2R_653\, 
        S => \I2.RPAGEL15R_516\, Y => \I2.N_623\);
    
    \I3.VDBI_57_0_IV_0_0L24R_2158\ : AO21
      port map(A => \I3.VDBil24r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l24r_adt_net_138805_\, Y => 
        \I3.VDBi_57l24r_adt_net_138815_\);
    
    \I2.STATE2l2r_adt_net_855212_\ : BFR
      port map(A => \I2.STATE2L2R_589\, Y => 
        \I2.STATE2l2r_adt_net_855212__net_1\);
    
    \I2.PIPE7_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl16r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl16r_net_1\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620_\ : BFR
      port map(A => \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\, Y
         => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620__net_1\);
    
    \I3.VDBi_16_m_i_o3l3r_884\ : OR2
      port map(A => \I3.REGMAPL8R_741\, B => 
        \I3.REGMAPl9r_adt_net_854320__net_1\, Y => 
        \I3.N_1907_262\);
    
    \I3.VDBI_57_0_IVL12R_2205\ : AND2
      port map(A => \I3.VDBil12r_net_1\, B => 
        \I3.N_1764_adt_net_854352__net_1\, Y => 
        \I3.VDBi_57l12r_adt_net_140988_\);
    
    \I3.VADm_0_a3l11r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl11r_net_1\, Y => \I3.VADml11r\);
    
    \I2.G_EVNT_NUM_n10_0_o2_1286\ : NAND2
      port map(A => \I2.N_207_550\, B => \I2.G_EVNT_NUMl9r_net_1\, 
        Y => \I2.N_218_548\);
    
    \I2.PIPE4_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl3r_net_1\);
    
    \I2.N_3234_adt_net_855648_\ : BFR
      port map(A => \I2.N_3234\, Y => 
        \I2.N_3234_adt_net_855648__net_1\);
    
    \I2.PIPE5_DT_702\ : MUX2L
      port map(A => \I2.PIPE5_DTl26r_net_1\, B => 
        \I2.PIPE4_DTl26r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_702_net_1\);
    
    \I2.PIPE10_DT_613\ : MUX2L
      port map(A => \I2.PIPE10_DTl8r_net_1\, B => 
        \I2.PIPE9_DTl8r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_613_net_1\);
    
    \I5.SDAout_82\ : MUX2H
      port map(A => \I5.SDAout_net_1\, B => \I5.SDAout_12\, S => 
        TICKL0R_3, Y => \I5.SDAout_82_net_1\);
    
    \I3.un1_noe16wi_0_a2_i\ : OR2FT
      port map(A => \I3.N_268\, B => \I3.WRITES_8\, Y => NOE16W_c);
    
    \I1.REG_74_12L268R_1946\ : NOR2
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__761\, B
         => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854404__net_1\, 
        Y => \I1.N_145_12_adt_net_123179_\);
    
    \I1.REG_74_0_IVL350R_1863\ : NOR2FT
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_24_sqmuxa_adt_net_854780__net_1\, Y => 
        \I1.REG_74l350r_adt_net_116117_\);
    
    \I2.L2TYPEl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_603_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl14r_net_1\);
    
    \I3.PIPEBl28r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEB_107_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl28r_net_1\);
    
    \I2.ROFFSET_907\ : MUX2H
      port map(A => \I2.ROFFSETl11r_net_1\, B => 
        \I2.ROFFSET_n11_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_907_net_1\);
    
    \I2.PIPE6_DT_454\ : MUX2H
      port map(A => \I2.PIPE5_DTl0r_net_1\, B => 
        \I2.PIPE6_DTl0r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_454_net_1\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l3r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl3r_net_1\, Q => 
        \I2.DIN_REG1_0l3r\);
    
    \I3.PIPEA_246\ : MUX2L
      port map(A => \I3.PIPEAl15r_net_1\, B => 
        \I3.PIPEA_8l15r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854668__net_1\, Y
         => \I3.PIPEA_246_net_1\);
    
    \I2.DTO_1l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_874_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l0r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I187_Y\ : XOR2FT
      port map(A => \I2.N502_i_0\, B => 
        \I2.ADD_21x21_fast_I187_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l17r\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I98_Y_1656\ : AND3FTT
      port map(A => \I2.N344\, B => \I2.N302\, C => \I2.N306\, Y
         => \I2.N460_adt_net_70355_\);
    
    \I3.STATE2l4r\ : DFFS
      port map(CLK => CLK_c, D => \I3.STATE2_nsl0r\, SET => 
        CLEAR_STAT_i_0, Q => \I3.STATE2l4r_net_1\);
    
    N_1_I3_TCNT3_c4 : AND2
      port map(A => \I3.TCNT3_i_0_il4r_net_1\, B => \I3.TCNT3_c3\, 
        Y => \I3.TCNT3_c4\);
    
    \I2.PIPE1_DT_42_1_IVL0R_1520\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl16r_net_1\, Y => 
        \I2.PIPE1_DT_42l0r_adt_net_52231_\);
    
    \I5.REG_1_27\ : MUX2H
      port map(A => \I5.SENS_ADDRl0r_net_1\, B => REGl444r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_27_net_1\);
    
    \I2.PIPE4_DTL7R_2964\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL7R_481\);
    
    \I5.SSTATE1SE_12_I_903\ : AND2
      port map(A => TICKL0R_557, B => \I5.sstate1l1r_net_1\, Y
         => \I5.sstate1se_12_i_adt_net_8689_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I111_Y\ : AOI21TTF
      port map(A => \I2.N469\, B => 
        \I2.I111_un1_Y_adt_net_71419_\, C => 
        \I2.N445_i_adt_net_71447_\, Y => \I2.N445_i\);
    
    \I2.MIC_REG2l7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_316_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2l7r_net_1\);
    
    \I3.REG_1_217\ : MUX2L
      port map(A => VDB_inl4r, B => REGl410r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_217_0\);
    
    \I2.PIPE8_DT_16l19r\ : AND2
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855164__net_1\, B => 
        \I2.N_585\, Y => \I2.PIPE8_DT_16l19r_net_1\);
    
    \I2.DTO_9_iv_0l20r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl20r_net_1\, 
        C => \I2.DTO_9l20r_adt_net_30726_\, Y => \I2.DTO_9l20r\);
    
    \I2.OFFSET_37_25l3r\ : MUX2L
      port map(A => \REGl256r\, B => \REGl192r\, S => 
        \I2.PIPE7_DTL27R_90\, Y => \I2.N_830\);
    
    \I3.PIPEA1l14r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_312_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l14r_net_1\);
    
    \I1.REG_1_178\ : MUX2H
      port map(A => \REGl277r\, B => \I1.REG_74l277r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\, Y => 
        \I1.REG_1_178_net_1\);
    
    \I3.REG_1l77r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_178_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl77r);
    
    \I3.PIPEB_87_2336\ : NOR2FT
      port map(A => \I3.PIPEBl8r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_87_adt_net_160377_\);
    
    \I2.WOFFSETl4r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.WOFFSETl4r_adt_net_854980__net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl4r_Rd1__net_1\);
    
    \I2.un1_tdc_res_41_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl408r, Y => 
        \I2.N_4622_i_0\);
    
    REGl292r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_193_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl292r\);
    
    \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854396_\ : BFR
      port map(A => \I1.PAGECNT_0l8r_adt_net_834720_Rd1__net_1\, 
        Y => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854396__net_1\);
    
    \I2.REG_1_C14_I_1736\ : OA21FTF
      port map(A => REGl46r, B => \I2.N_3859\, C => 
        \I2.un8_evread_1_adt_net_855784__net_1\, Y => 
        \I2.N_3843_adt_net_101094_\);
    
    \I3.VDBi_57_0_iv_0_o3l13r\ : OR2
      port map(A => \I3.N_1764_adt_net_854352__net_1\, B => 
        \I3.STATE1_nsl8r_adt_net_136092_\, Y => \I3.N_56\);
    
    \I3.STATE1l9r_1624\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL9R_731\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l7r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl7r_net_1\, Q => 
        \I2.DIN_REG1l7r\);
    
    \I3.VDBI_57_IV_0_0_O2_0_8_TZL0R_2270\ : NOR2
      port map(A => GA_cl0r, B => \I3.N_2042\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_adt_net_146105_\);
    
    \I3.VDBi_23_0_a2_0l1r\ : NAND2FT
      port map(A => \I3.REGMAPL7R_459\, B => \I3.REGMAPL3R_738\, 
        Y => \I3.N_2042\);
    
    \I3.VASl11r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_73_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl11r_net_1\);
    
    \I2.resyn_0_I2_BITCNT_937\ : MUX2H
      port map(A => \I2.BITCNTl3r_net_1\, B => \I2.N_4324\, S => 
        \I2.BITCNTe\, Y => \I2.BITCNT_937\);
    
    \I2.LSRAM_INl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_401_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl17r_net_1\);
    
    \I2.PIPE6_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_460_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl6r_net_1\);
    
    \I2.PIPE2_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl10r_net_1\);
    
    \I3.VDBi_52l3r\ : MUX2H
      port map(A => \I3.VDBil3r_net_1\, B => \FBOUTl3r\, S => 
        \I3.N_57_i_0_0_adt_net_854696__net_1\, Y => 
        \I3.VDBi_52l3r_net_1\);
    
    \I2.WROi\ : DFFS
      port map(CLK => CLK_c, D => \I2.WROi_793_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.WROi_net_1\);
    
    DTO_padl22r : IOB33PH
      port map(PAD => DTO(22), A => \I2.DTO_1l22r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl22r);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2281\ : AO21
      port map(A => \I3.N_2014\, B => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146446_\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146424_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146448_\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2195\ : AND2
      port map(A => \I3.PIPEAl13r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l13r_adt_net_140578_\);
    
    \I3.VDBOFFB_30_IV_0L4R_2419\ : OR3
      port map(A => \I3.VDBoffb_30l4r_adt_net_162367_\, B => 
        \I3.VDBoffb_30l4r_adt_net_162363_\, C => 
        \I3.VDBoffb_30l4r_adt_net_162364_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162370_\);
    
    \I3.END_PK\ : DFFC
      port map(CLK => CLK_c, D => \I3.END_PK_229_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.END_PK_net_1\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l5r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl5r_net_1\, Q => 
        \I2.DIN_REG1l5r\);
    
    \I1.REG_1_195\ : MUX2H
      port map(A => \REGl294r\, B => \I1.REG_74l294r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\, Y => 
        \I1.REG_1_195_net_1\);
    
    \I3.VDBi_357\ : MUX2L
      port map(A => \I3.VDBil17r_net_1\, B => \I3.VDBi_57l17r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_357_net_1\);
    
    \I2.DTO_16_1_IV_0_0L18R_1126\ : AND2
      port map(A => \I2.DTO_1l18r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l18r_adt_net_31333_\);
    
    \I3.PIPEA_261\ : MUX2L
      port map(A => \I3.PIPEAl30r_net_1\, B => 
        \I3.PIPEA_8l30r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854652__net_1\, Y
         => \I3.PIPEA_261_net_1\);
    
    \I2.N_2867_1_adt_net_854964_\ : BFR
      port map(A => \I2.N_2867_1_338\, Y => 
        \I2.N_2867_1_adt_net_854964__net_1\);
    
    \I2.L2TYPEl14r_1549\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_603_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL14R_656\);
    
    \I2.PIPE7_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl12r_net_1\);
    
    \I3.VASl8r_969\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_70_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASL8R_347\);
    
    \I1.REG_74_1_396_m7_i_1\ : NOR3FTT
      port map(A => \I1.PAGECNT_0l9r_adt_net_835132_Rd1__net_1\, 
        B => \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_1_RD1__458\, C => 
        \PULSEl0r\, Y => \I1.REG_74_8_308_m9_i_1\);
    
    \I3.REG_1_ml64r\ : AND2
      port map(A => REGl64r, B => 
        \I3.REGMAPl9r_adt_net_854312__net_1\, Y => 
        \I3.VDBi_20l16r\);
    
    \I1.REG_74_0_IVL333R_1883\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l333r_adt_net_117830_\);
    
    \I2.LEAD_FLAG6_7_i_0l0r\ : AOI21
      port map(A => \I2.N_217\, B => \I2.N_483\, C => \I2.N_222\, 
        Y => \I2.N_4535_adt_net_64588_\);
    
    \I3.REG_1_263\ : MUX2H
      port map(A => REGl82r, B => VDB_inl0r, S => \I3.N_2277_i\, 
        Y => \I3.REG_1_263_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I137_Y_i\ : AO21TTF
      port map(A => \I2.N_40_adt_net_1100__net_1\, B => 
        \I2.N_40_adt_net_57971_\, C => \I2.N_92\, Y => \I2.N_40\);
    
    \I2.PIPE5_DT_6_0l5r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l5r\, B => 
        \I2.un27_pipe5_dt0l5r\, S => 
        \I2.dataout_0_adt_net_855808__net_1\, Y => \I2.N_1074\);
    
    \I2.N_3834_i_0_adt_net_1384_\ : NAND2FT
      port map(A => \I2.un8_evread_1_adt_net_855792__net_1\, B
         => \I2.N_3847\, Y => \I2.N_3834_i_0_adt_net_1384__net_1\);
    
    \I1.REG_1_197\ : MUX2H
      port map(A => \REGl296r\, B => \I1.REG_74l296r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\, Y => 
        \I1.REG_1_197_net_1\);
    
    \I2.PIPE7_DTl5r_1593\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl5r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL5R_700\);
    
    \I2.DTE_21_1l11r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l11r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l11r_Rd1__net_1\);
    
    \I1.PAGECNT_0L9R_ADT_NET_835132_RD1__3098\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854852__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0L9R_ADT_NET_835132_RD1__884\);
    
    \I3.REGMAPL9R_3032\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un41_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL9R_786\);
    
    \I2.PIPE1_DT_2_SQMUXA_ADT_NET_803__2874\ : OR2FT
      port map(A => \I2.TDCGDA1_net_1\, B => 
        \I2.NWPIPE1_4_SQMUXA_1_0_301\, Y => 
        \I2.PIPE1_DT_2_SQMUXA_ADT_NET_803__299\);
    
    \I2.L2TYPEl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_596_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEl7r_net_1\);
    
    \I2.PIPE7_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl6r_net_1\);
    
    \I2.WOFFSETl3r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.WOFFSETl3r_adt_net_854988__net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl3r_Rd1__net_1\);
    
    REGl399r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_300_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl399r\);
    
    \I2.PIPE7_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl25r_net_1\);
    
    \I2.L2AS_adt_net_855716_\ : BFR
      port map(A => \I2.L2AS_adt_net_855720__net_1\, Y => 
        \I2.L2AS_adt_net_855716__net_1\);
    
    \I2.PIPE8_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_539_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl11r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I56_Y\ : AO21
      port map(A => \I2.N267_0\, B => \I2.N308_0_adt_net_86492_\, 
        C => \I2.N304_0_adt_net_87004_\, Y => \I2.N306_i_i\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2201\ : AO21
      port map(A => \I3.VDBil13r_net_1\, B => \I3.N_56\, C => 
        \I3.VDBi_57l13r_adt_net_140594_\, Y => 
        \I3.VDBi_57l13r_adt_net_140596_\);
    
    \I3.VDBm_0l22r\ : MUX2L
      port map(A => \I3.PIPEAl22r_net_1\, B => 
        \I3.PIPEBl22r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_164\);
    
    \I2.DTE_21_1_IV_0L28R_1234\ : AO21FTF
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, 
        B => \I2.DT_TEMPl28r_net_1\, C => \I2.N_223\, Y => 
        \I2.DTE_21_1l28r_adt_net_36757_\);
    
    \I3.PIPEA_8l19r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854468__net_1\, B => 
        \I3.N_228\, Y => \I3.PIPEA_8l19r_net_1\);
    
    \I2.CRC32_12_0_0_x2l5r\ : XOR2FT
      port map(A => \I2.CRC32l5r_net_1\, B => \I2.N_4267_i_i\, Y
         => \I2.N_131_i_0_i_0\);
    
    \I2.DTE_21_1_IV_0L13R_1286\ : AO21
      port map(A => \I2.DT_TEMPl13r_net_1\, B => \I2.N_4038\, C
         => \I2.DTE_21_1l13r_adt_net_38165_\, Y => 
        \I2.DTE_21_1l13r_adt_net_38179_\);
    
    TDCDA_padl31r : IB33
      port map(PAD => TDCDA(31), Y => TDCDA_cl31r);
    
    \I3.STATE1_tr24_i_0\ : OA21TTF
      port map(A => \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135633_\, 
        B => \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135642_\, C => 
        \I3.un1_REGMAP_34\, Y => \I3.STATE1_tr24_i_0_net_1\);
    
    \I2.DT_TEMP_7l11r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, B => 
        \I2.DT_SRAMl11r_net_1\, Y => \I2.DT_TEMP_7l11r_net_1\);
    
    \I1.PAGECNTlde_0_a2_0_1\ : OR2FT
      port map(A => \I1.N_341_RD1__487\, B => 
        \I1.N_591_1_adt_net_106236_Rd1__net_1\, Y => \I1.N_591_1\);
    
    \I3.VDBm_0l4r\ : MUX2L
      port map(A => \I3.PIPEAl4r_net_1\, B => \I3.PIPEBl4r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_146\);
    
    \I2.un1_sram_evnt12_i_a2_0\ : NOR2
      port map(A => \I2.START_GIRO_net_1\, B => \I2.N_3850\, Y
         => \I2.N_132\);
    
    \I2.WPAGEL15R_2995\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_948_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEL15R_749\);
    
    \I2.DTE_1l21r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l21r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l21r_Rd1__net_1\);
    
    \I2.MIC_ERR_REGS_329\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl1r_net_1\, B => 
        \I2.MIC_ERR_REGSl0r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_329_net_1\);
    
    \I3.REG_1l163r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_211_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl163r\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I162_Y_1691\ : OA21TTF
      port map(A => \I2.N348\, B => \I2.N355_0\, C => 
        \I2.N479_adt_net_642225_\, Y => 
        \I2.N489_i_adt_net_89351_\);
    
    \I1.REG_74_0_ivl384r\ : AO21
      port map(A => \REGl384r\, B => \I1.N_257\, C => 
        \I1.REG_74l384r_adt_net_111663_\, Y => \I1.REG_74l384r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I27_Y\ : AO21
      port map(A => \I2.SUB8l15r_net_1\, B => \I2.SUB8l14r_net_1\, 
        C => \I2.N292_adt_net_68955_\, Y => \I2.N292\);
    
    \I2.PIPE4_DTL6R_2962\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL6R_479\);
    
    \I1.REG_74_0_iv_0l357r\ : AO21
      port map(A => \REGl357r\, B => \I1.N_661\, C => 
        \I1.REG_74l357r_adt_net_115127_\, Y => \I1.REG_74l357r\);
    
    \I5.PULSE_I2C\ : MUX2L
      port map(A => \I5.AIR_PULSE_net_1\, B => PULSEl7r, S => 
        REGl7r, Y => \I5.PULSE_I2C_net_1\);
    
    \I2.OFFSET_37_1l2r\ : MUX2L
      port map(A => \REGl351r\, B => \REGl287r\, S => 
        \I2.PIPE7_DTL27R_66\, Y => \I2.N_637\);
    
    \I2.RAMDT4L2R_3013\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl2r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L2R_767\);
    
    \I1.BYTECNT_311\ : MUX2H
      port map(A => \I1.BYTECNTl3r_net_1\, B => \I1.BYTECNT_n3\, 
        S => \I1.N_1383\, Y => \I1.BYTECNT_311_net_1\);
    
    \I1.REG_74_0_IVL238R_1988\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_10_sqmuxa_adt_net_854720__net_1\, Y => 
        \I1.REG_74l238r_adt_net_126899_\);
    
    \I2.MIC_ERR_REGSl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_346_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl17r_net_1\);
    
    \I2.PIPE8_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_536_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl8r_net_1\);
    
    \I2.REG_1_c12_i_a2_0\ : AND3FFT
      port map(A => REGl43r, B => REGl44r, C => \I2.N_131\, Y => 
        \I2.N_136_1\);
    
    \I2.PIPE6_DT_455\ : MUX2H
      port map(A => \I2.PIPE5_DTl1r_net_1\, B => 
        \I2.PIPE6_DTl1r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_455_net_1\);
    
    \I2.PIPE7_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl17r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl17r_net_1\);
    
    \I3.VDBml28r\ : MUX2L
      port map(A => \I3.VDBil28r_net_1\, B => \I3.N_170\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml28r_net_1\);
    
    \I2.G_EVNT_NUM_n6_i_o2_1290\ : AND2FT
      port map(A => \I2.N_4669_adt_net_855052__net_1\, B => 
        \I2.G_EVNT_NUMl5r_net_1\, Y => \I2.N_4672_552\);
    
    FID_padl12r : OB33PH
      port map(PAD => FID(12), A => FID_cl12r);
    
    \I2.DTE_2_1l8r\ : XOR2
      port map(A => \I2.CRC32l28r_net_1\, B => 
        \I2.DTE_2_1_0l8r_net_1\, Y => \I2.DTE_2_1l8r_net_1\);
    
    \I3.VDBi_40_0_i_m2l1r\ : MUX2L
      port map(A => REGl419r, B => REGl435r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_133\);
    
    \I3.PURGED\ : DFFS
      port map(CLK => CLK_c, D => \I3.PURGED_43_net_1\, SET => 
        \I3.N_2137_i_0\, Q => \I3.PURGED_net_1\);
    
    \I3.REGMAPl14r_1627\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un57_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL14R_734\);
    
    \I3.TCNT2l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT2_391_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT2l5r_net_1\);
    
    \I1.REG_1_71\ : MUX2H
      port map(A => \REGl170r\, B => \I1.REG_74l170r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, Y => 
        \I1.REG_1_71_net_1\);
    
    \I2.SUB9_580\ : MUX2H
      port map(A => \I2.SUB9l12r_net_1\, B => \I2.SUB9_1l12r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_580_net_1\);
    
    \I2.LEAD_FLAG6_637\ : AO21
      port map(A => \I2.N_4535_adt_net_1178__net_1\, B => 
        \I2.N_4535_adt_net_64588_\, C => 
        \I2.LEAD_FLAG6_637_adt_net_64628_\, Y => 
        \I2.LEAD_FLAG6_637_net_1\);
    
    \I2.FIFO_FULL_1485\ : DFFC
      port map(CLK => CLK_c, D => PAF_c_i_0, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.FIFO_FULL_592\);
    
    RAMDT_padl8r : IOB33PH
      port map(PAD => RAMDT(8), A => \I1.RAMDT_SPI_1l1r_net_1\, 
        EN => \I1.RAMDT_SPI_e_net_1\, Y => RAMDT_inl8r);
    
    \I1.REG_74_0_IV_0_0L256R_1969\ : AND2
      port map(A => \FBOUTl3r\, B => \I1.N_596\, Y => 
        \I1.REG_74l256r_adt_net_125142_\);
    
    \I2.OFFSET_37_28l2r\ : MUX2L
      port map(A => \I2.N_845\, B => \I2.N_797\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_853\);
    
    VDB_padl15r : IOB33PH
      port map(PAD => VDB(15), A => \I3.VDBml15r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl15r);
    
    \I3.PULSEl4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_334_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl4r);
    
    \I3.VDBoffl7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_123_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl7r_net_1\);
    
    \I2.SUB9_575\ : MUX2H
      port map(A => \I2.SUB9l7r_net_1\, B => \I2.SUB9_1l7r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_575_net_1\);
    
    \I2.L2SERV_c2\ : NAND2
      port map(A => \I2.RPAGEL14R_616\, B => \I2.L2SERV_c1_net_1\, 
        Y => \I2.L2SERV_c2_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I190_Y\ : XOR2FT
      port map(A => \I2.N_1_1_0\, B => 
        \I2.ADD_21x21_fast_I190_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l20r\);
    
    N_1_I3_TCNT3_c6 : NAND2
      port map(A => \I3.TCNT3_i_0_il6r_net_1\, B => 
        \N_1.I3.TCNT3_c5\, Y => \N_1.I3.TCNT3_c6\);
    
    \I3.VDBOFFB_30_IV_0_0L5R_2400\ : OR3
      port map(A => \I3.VDBoffb_30l5r_adt_net_162175_\, B => 
        \I3.VDBoffb_30l5r_adt_net_162169_\, C => 
        \I3.VDBoffb_30l5r_adt_net_162170_\, Y => 
        \I3.VDBoffb_30l5r_adt_net_162179_\);
    
    \I1.REG_1_193\ : MUX2H
      port map(A => \REGl292r\, B => \I1.REG_74l292r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\, Y
         => \I1.REG_1_193_net_1\);
    
    \I2.STATE1_ns_a3_il12r\ : NOR3FFT
      port map(A => TDCDRYB_c, B => 
        \I2.N_3887_adt_net_855068__net_1\, C => \I2.N_3889\, Y
         => \I2.N_3875_i_0\);
    
    TOKOUTA_BP_pad : IB33
      port map(PAD => TOKOUTA_BP, Y => TOKOUTA_BP_c);
    
    \I2.DTO_cl_29l31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_cl_64_il31r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.DTO_cll31r\);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_1_sqmuxa_0_a4_i_o2\ : AO21FTT
      port map(A => \I2.PIPE4_DTl23r_net_1\, B => 
        \I2.N_4524_adt_net_16701_\, C => 
        \I2.N_4524_adt_net_16804_\, Y => \I2.N_4524\);
    
    \I2.OFFSET_37_6l1r\ : MUX2L
      port map(A => \I2.N_668\, B => \I2.N_660\, S => 
        \I2.PIPE7_DTL26R_354\, Y => \I2.N_676\);
    
    \I2.PIPE9_DT_288\ : MUX2L
      port map(A => \I2.PIPE9_DTl19r_net_1\, B => 
        \I2.PIPE8_DTl19r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_288_net_1\);
    
    VAD_padl25r : OTB33PH
      port map(PAD => VAD(25), A => \I3.VADml25r\, EN => 
        NOEAD_c_i_0);
    
    \I3.PIPEA1l9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_307_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l9r_net_1\);
    
    \I1.REG_1_94\ : MUX2H
      port map(A => \REGl193r\, B => \I1.REG_74l193r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855416__net_1\, Y => 
        \I1.REG_1_94_net_1\);
    
    \I2.DT_SRAMl31r\ : MUX2L
      port map(A => \I2.N_899\, B => \I2.PIPE2_DTl31r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl31r_net_1\);
    
    \I2.MIC_REG2L2R_2946\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_311_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2L2R_463\);
    
    \I2.PIPE10_DT_619\ : MUX2L
      port map(A => \I2.PIPE10_DTl14r_net_1\, B => \I2.N_3800\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_619_net_1\);
    
    \I2.BNCID_VECTrff_6\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_6_259_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_6\);
    
    \I2.L2TYPE_4_IL1R_1639\ : NAND2FT
      port map(A => \I2.N_4457\, B => \I2.N_4461\, Y => 
        \I2.N_4451_adt_net_68574_\);
    
    \I1.N_370_adt_net_854904_\ : BFR
      port map(A => \I1.N_370\, Y => 
        \I1.N_370_adt_net_854904__net_1\);
    
    \I2.ADO_3l2r\ : MUX2L
      port map(A => \I2.WOFFSETl3r_adt_net_854988__net_1\, B => 
        \I2.ROFFSETl3r_net_1\, S => NOESRAME_C_243, Y => 
        \I2.ADO_3l2r_net_1\);
    
    \I3.STATE2_ns_0l4r\ : AO21
      port map(A => \I3.N_1465\, B => \I3.STATE2l1r_net_1\, C => 
        \I3.N_1879\, Y => \I3.STATE2_nsl4r\);
    
    \I5.SDAout\ : DFFS
      port map(CLK => CLK_c, D => \I5.SDAout_82_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SDAout_net_1\);
    
    \I2.CRC32l9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_804_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l9r_net_1\);
    
    \I3.PIPEBl12r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_91_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl12r_net_1\);
    
    \I2.OFFSETl4r_1568\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_564_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL4R_675\);
    
    \I2.STATE3_NS_O3_0L8R_1039\ : NAND3FFT
      port map(A => REGl2r, B => \I2.N_3015\, C => 
        \I2.N_118_i_1_adt_net_1122__net_1\, Y => 
        \I2.N_3012_adt_net_24327_\);
    
    \I2.STATE1_ns_i_o2l8r\ : AOI21FTF
      port map(A => \I2.STATE1l12r_adt_net_855184__net_1\, B => 
        \I2.N_3273\, C => \I2.N_3344_i\, Y => \I2.N_3275\);
    
    \I2.SUB9_1_ADD_18x18_fast_I151_Y\ : XOR2FT
      port map(A => \I2.N451_i\, B => 
        \I2.ADD_18x18_fast_I151_Y_0\, Y => \I2.SUB9_1l14r\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__2971\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__488\);
    
    \I2.DTE_21_1_IV_0_0L17R_1222\ : AND2
      port map(A => \I2.DTE_1l17r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\, Y => 
        \I2.DTE_21_1l17r_adt_net_36142_\);
    
    \I2.PIPE8_DTl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_533_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl5r_net_1\);
    
    \I2.L2TYPE_4_IL9R_1625\ : OR2
      port map(A => \I2.N_4457\, B => \I2.N_4459\, Y => 
        \I2.N_4443_adt_net_67572_\);
    
    \I2.OFFSET_37_4l7r\ : MUX2L
      port map(A => \REGl372r\, B => \REGl308r\, S => 
        \I2.PIPE7_DTL27R_67\, Y => \I2.N_666\);
    
    \I2.L2AF1\ : DFFC
      port map(CLK => CLK_c, D => L2A_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.L2AF1_net_1\);
    
    \I1.REG_74_0_iv_0l173r\ : AO21
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, C => 
        \I1.REG_74l173r_adt_net_132940_\, Y => \I1.REG_74l173r\);
    
    \I5.REG_1l440r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_23_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl440r);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I24_G0N\ : AND2FT
      port map(A => \I2.LSRAM_OUTl3r\, B => \I2.PIPE7_DTL3R_701\, 
        Y => \I2.N239\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I136_Y_0_o2_m2_e\ : AO21
      port map(A => \I2.PIPE4_DTL13R_641\, B => 
        \I2.PIPE4_DTL14R_638\, C => \I2.RAMDT4L12R_145\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_N_6_i_adt_net_56543_\);
    
    \I2.G_EVNT_NUM_925\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl9r_net_1\, B => 
        \I2.G_EVNT_NUM_n9\, S => \I2.N_3769\, Y => 
        \I2.G_EVNT_NUM_925_net_1\);
    
    \I2.OFFSET_37_14l2r\ : MUX2L
      port map(A => \I2.N_733\, B => \I2.N_685\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_741\);
    
    \I1.REG_74_0_IVL171R_2063\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l171r_adt_net_133149_\);
    
    \I2.DTE_21_1_iv_0_il25r\ : AO21
      port map(A => \I2.DTE_1l25r\, B => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, C => 
        \I2.N_4644_adt_net_37065_\, Y => \I2.N_4644\);
    
    \I1.REG_74_0_ivl231r\ : AO21
      port map(A => \REGl231r\, B => \I1.N_105\, C => 
        \I1.REG_74l231r_adt_net_127538_\, Y => \I1.REG_74l231r\);
    
    \I2.SUB8_522_2734\ : AND3
      port map(A => \I2.N477_adt_net_371248_\, B => 
        \I2.N477_adt_net_371301_\, C => 
        \I2.SUB8_522_adt_net_551987_\, Y => 
        \I2.SUB8_522_adt_net_659160_\);
    
    \I3.VDBi_364\ : MUX2L
      port map(A => \I3.VDBil24r_net_1\, B => \I3.VDBi_57l24r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_364_net_1\);
    
    \I3.REG_1_284\ : MUX2L
      port map(A => VDB_inl2r, B => REGl103r, S => 
        \I3.N_318_adt_net_855888__net_1\, Y => \I3.REG_1_284_0\);
    
    \I3.VDBml24r\ : MUX2L
      port map(A => \I3.VDBil24r_net_1\, B => \I3.N_166\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml24r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L3R_2576\ : AO21
      port map(A => \REGl264r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        C => \I3.VDBoffa_31l3r_adt_net_164044_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164073_\);
    
    \I3.REG1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG1_138_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l5r_net_1\);
    
    \I2.I_1342_ca_0_and2\ : NOR2FT
      port map(A => \I2.SUB8l10r_net_1\, B => \I2.OFFSETL7R_670\, 
        Y => \I2.N_3547_i_i\);
    
    \I3.TCNT4_i_0_il0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT4_388_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT4_i_0_il0r_net_1\);
    
    \I2.PIPE6_DT_0_SQMUXA_I_O4_1596\ : AO21
      port map(A => \I2.N_215\, B => \I2.N_4544\, C => 
        \I2.N_4551_adt_net_63747_\, Y => 
        \I2.N_4551_adt_net_63758_\);
    
    \I2.N507_adt_net_347771_\ : AO21FTT
      port map(A => \I2.N_70_adt_net_255802__net_1\, B => 
        \I2.N507_adt_net_347769__net_1\, C => 
        \I2.N507_adt_net_347770__net_1\, Y => 
        \I2.N507_adt_net_347771__net_1\);
    
    \I2.LEAD_FLAG6_643_1600\ : NOR2FT
      port map(A => LEAD_FLAGl6r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_643_adt_net_63956_\);
    
    \I2.SUB8l12r_adt_net_855576_\ : BFR
      port map(A => \I2.SUB8l12r_net_1\, Y => 
        \I2.SUB8l12r_adt_net_855576__net_1\);
    
    \I2.DTO_16_1_ivl3r\ : OA21FTF
      port map(A => \I2.N_182_ADT_NET_1007__386\, B => 
        \I2.DT_SRAMl3r_net_1\, C => \I2.DTO_16_1_iv_1l3r_net_1\, 
        Y => \I2.DTO_16_1_ivl3r_net_1\);
    
    \I1.REG_1_196\ : MUX2H
      port map(A => \REGl295r\, B => \I1.REG_74l295r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\, Y => 
        \I1.REG_1_196_net_1\);
    
    \I1.BITCNTL2R_2999\ : DFFC
      port map(CLK => CLK_c, D => \I1.BITCNT_315_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BITCNTL2R_753\);
    
    \I3.PULSE_46_0_iv_i_i_a3_0l7r\ : AND2
      port map(A => \I3.REGMAP_i_0_il15r\, B => 
        \I3.N_1906_i_0_0_adt_net_855636__net_1\, Y => \I3.N_318\);
    
    \I3.VDBOFFB_30_IV_0L7R_2349\ : AND2
      port map(A => \REGl356r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161748_\);
    
    \I1.REG_74_8_0_324_m6_e\ : NAND2
      port map(A => \I1.PAGECNTL7R_526\, B => 
        \I1.REG_74_1_a0_0l228r\, Y => 
        \I1.REG_74_8_0_324_m6_e_net_1\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2196\ : AND3FFT
      port map(A => \I3.N_2014\, B => \I3.N_1917\, C => 
        \I3.REGl146r\, Y => \I3.VDBi_57l13r_adt_net_140582_\);
    
    \I2.RAMAD1_12l6r\ : MUX2L
      port map(A => \I2.TDCDASl4r_net_1\, B => 
        \I2.TDCDBSl4r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855180__net_1\, Y => 
        \I2.RAMAD1_12l6r_net_1\);
    
    \I1.REG_74_0_IVL239R_1987\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_10_sqmuxa_adt_net_854720__net_1\, Y => 
        \I1.REG_74l239r_adt_net_126813_\);
    
    \I2.L2TYPE_4_IL0R_1641\ : NAND2
      port map(A => \I2.N_4458\, B => \I2.N_4461\, Y => 
        \I2.N_4452_adt_net_68713_\);
    
    \I1.REG_74_0_ivl358r\ : AO21
      port map(A => \REGl358r\, B => \I1.N_661\, C => 
        \I1.REG_74l358r_adt_net_115041_\, Y => \I1.REG_74l358r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I151_Y_0\ : XOR2FT
      port map(A => \I2.SUB8l15r_adt_net_855572__net_1\, B => 
        \I2.SUB8l14r_adt_net_855568__net_1\, Y => 
        \I2.ADD_18x18_fast_I151_Y_0\);
    
    \I1.RAMDT_SPI_1l2r\ : DFFC
      port map(CLK => CLK_c, D => \FBOUTl2r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.RAMDT_SPI_1l2r_net_1\);
    
    \I1.NWRLUTi_57\ : MUX2L
      port map(A => \I1.N_1207\, B => \I1.NWRLUTi_net_1\, S => 
        \I1.N_1192\, Y => \I1.NWRLUTi_57_net_1\);
    
    \I3.TCNT_0_sqmuxa_0_a2_0_a3_0\ : NOR3FFT
      port map(A => \I3.WRITES_8\, B => \I3.REGMAPl51r_net_1\, C
         => \I3.N_276\, Y => \I3.TCNT_0_sqmuxa_0\);
    
    \I3.PIPEB_79\ : AO21
      port map(A => DPR_cl0r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855280__net_1\, 
        C => \I3.PIPEB_79_adt_net_160713_\, Y => 
        \I3.PIPEB_79_net_1\);
    
    \I2.PIPE1_DT_740\ : MUX2L
      port map(A => \I2.PIPE1_DTl13r_net_1\, B => 
        \I2.PIPE1_DT_42l13r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854576__net_1\, 
        Y => \I2.PIPE1_DT_740_net_1\);
    
    \I2.CRC32_12_0_0_m3l18r\ : MUX2L
      port map(A => \I2.DT_TEMPl18r_net_1\, B => 
        \I2.DTO_16_1l18r_adt_net_756__net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854196__net_1\, Y => 
        \I2.N_4096_i_i\);
    
    \I3.VDBI_57_IV_0_0L6R_2235\ : OA21TTF
      port map(A => \I3.VDBi_57l6r_adt_net_143327__net_1\, B => 
        \I3.VDBi_57l6r_adt_net_143328__net_1\, C => 
        \I3.N_1905_1_adt_net_855384__net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143394_\);
    
    \I2.FIDl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_420_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl4r);
    
    \I2.STATE2_ns_a6_2_a2_0l4r\ : AO21TTF
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996__net_1\, 
        B => \I2.N_4261_304\, C => \I2.N_223_156\, Y => 
        \I2.N_2864_0\);
    
    DPR_padl4r : IB33
      port map(PAD => DPR(4), Y => DPR_cl4r);
    
    \I2.L2TYPE_4_i_o2_0l12r\ : NOR2
      port map(A => \I2.L2ARRl1r_net_1\, B => \I2.L2ARRl0r_net_1\, 
        Y => \I2.N_4458\);
    
    \I3.REG_0_sqmuxa_2_adt_net_855292_\ : BFR
      port map(A => \I3.REG_0_sqmuxa_2\, Y => 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\);
    
    \I3.PIPEB_83_2340\ : NOR2FT
      port map(A => \I3.PIPEBl4r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_83_adt_net_160545_\);
    
    \I2.PIPE9_DT_291\ : MUX2L
      port map(A => \I2.PIPE9_DTl22r_net_1\, B => 
        \I2.PIPE8_DTl22r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_291_net_1\);
    
    \I2.REG_1_c2_i_o2\ : AND2
      port map(A => REGL34R_872, B => \I2.N_3844\, Y => 
        \I2.N_3845\);
    
    \I2.EVNT_NUMl2r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_961_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl2r_net_1\);
    
    \I1.REG_74_0_IVL232R_1994\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_9_sqmuxa_adt_net_854728__net_1\, Y => 
        \I1.REG_74l232r_adt_net_127452_\);
    
    \I2.un7_bnc_id_1_I_13\ : XOR2
      port map(A => \I2.BNC_IDl3r_net_1\, B => 
        \I2.DWACT_FINC_El0r\, Y => \I2.I_13_2\);
    
    \I2.RAMAD_4l16r\ : MUX2L
      port map(A => \I2.N_543\, B => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854392__net_1\, 
        S => LOAD_RES_1, Y => \I2.RAMAD_4l16r_net_1\);
    
    \I3.VDBm_0l20r\ : MUX2L
      port map(A => \I3.PIPEAl20r_net_1\, B => 
        \I3.PIPEBl20r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_162\);
    
    \I3.VASl13r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_75_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VAS_i_0_il13r\);
    
    \I2.RAMDT4l11r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl11r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l11r_net_1\);
    
    FID_padl0r : OB33PH
      port map(PAD => FID(0), A => FID_cl0r);
    
    \I3.un7_ronly_0_a2_0_a3\ : AND2
      port map(A => \I3.N_544\, B => 
        \I3.un7_ronly_0_a2_0_a3_adt_net_165588_\, Y => 
        \I3.un7_ronly_0_a2_0_a3_net_1\);
    
    DTO_padl26r : IOB33PH
      port map(PAD => DTO(26), A => \I2.DTO_1l26r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl26r);
    
    \I2.ROFFSET_n4_tz\ : XOR2
      port map(A => \I2.ROFFSETl4r_net_1\, B => 
        \I2.ROFFSET_c3_net_1\, Y => \I2.ROFFSET_n4_tz_i\);
    
    CHAINB_ERR_pad : IB33
      port map(PAD => CHAINB_ERR, Y => CHAINB_ERR_c);
    
    \I3.STATE2_ns_0_a3l4r\ : AND2FT
      port map(A => \I3.DSS_718\, B => \I3.STATE2l0r_net_1\, Y
         => \I3.N_1879\);
    
    \I2.TDCDASl15r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl15r, Q => 
        \I2.TDCDASl15r_net_1\);
    
    \I2.NWPIPE4_1468\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE3_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE4_575\);
    
    \I3.VDBoffl1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_117_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl1r_net_1\);
    
    \I3.STATE1_NS_1_IV_0L3R_2124\ : AND2FT
      port map(A => \I3.DSS_net_1\, B => \I3.STATE1_ipl7r\, Y => 
        \I3.STATE1_nsl3r_adt_net_136439_\);
    
    \I3.PIPEA_8l11r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854476__net_1\, B => 
        \I3.N_220\, Y => \I3.PIPEA_8l11r_net_1\);
    
    \I1.SSTATE_NS_1_IV_0_I_A4_2L8R_1764\ : AND2
      port map(A => \I1.sstatel3r_net_1\, B => PULSEl6r, Y => 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r_adt_net_107356_\);
    
    \I5.sstate1se_12_i\ : MUX2H
      port map(A => \I5.sstate1l0r_net_1\, B => 
        \I5.sstate1l1r_net_1\, S => TICKl0r, Y => 
        \I5.sstate1se_12_i_net_1\);
    
    \I2.resyn_0_I2_FID_429\ : MUX2H
      port map(A => FID_cl13r, B => \I2.FID_7l13r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\, 
        Y => \I2.FID_429\);
    
    \I1.REG_74_0_IV_I_A2L203R_2031\ : AND2
      port map(A => \REGl203r\, B => \I1.N_182_i\, Y => 
        \I1.N_1342_adt_net_130275_\);
    
    \I2.REG_1l36r_1458\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL36R_565);
    
    \I2.PIPE9_DT_287\ : MUX2L
      port map(A => \I2.PIPE9_DTl18r_net_1\, B => 
        \I2.PIPE8_DTl18r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_287_net_1\);
    
    \I2.EVNT_WORDl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_717_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl4r_net_1\);
    
    \I2.PIPE8_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_556_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl28r_net_1\);
    
    \I3.REG_1_267\ : MUX2H
      port map(A => REGl86r, B => \I3.N_1632\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_267_0\);
    
    \I2.RAMAD1l2r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_656_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l2r_net_1\);
    
    \I2.PIPE10_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_626_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl21r_net_1\);
    
    \I3.REG1_140\ : MUX2L
      port map(A => VDB_inl7r, B => \I3.REG1l7r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855628__net_1\, Y => 
        \I3.REG1_140_net_1\);
    
    \I2.TRGARR_3_I_15\ : XOR2
      port map(A => \I2.DWACT_ADD_CI_0_TMPl0r\, B => 
        \I2.TRGARRl1r_net_1\, Y => \I2.TRGARR_3l1r\);
    
    \I1.REG_1_120\ : MUX2H
      port map(A => \REGl219r\, B => \I1.REG_74l219r\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_120_net_1\);
    
    \I2.DTE_21_1_IV_0_0_18_M7_1217\ : AND3FTT
      port map(A => 
        \I2.REG_0l3r_adt_net_848__adt_net_854216__net_1\, B => 
        \I2.STATE2l1r_adt_net_855124__net_1\, C => REGl29r, Y => 
        \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35897_\);
    
    \I5.REG_1l425r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_38_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl425r);
    
    \I3.VDBi_57l8r_adt_net_1606_\ : AO21
      port map(A => \I3.N_2016\, B => \I3.VDBi_29l8r_net_1\, C
         => \I3.VDBi_57l8r_adt_net_142596__net_1\, Y => 
        \I3.VDBi_57l8r_adt_net_1606__net_1\);
    
    \I1.RAMDT_SPI_1l6r\ : DFFC
      port map(CLK => CLK_c, D => \FBOUTl6r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.RAMDT_SPI_1l6r_net_1\);
    
    \I3.TCNT_n1_0_0\ : AO21FTF
      port map(A => \I3.un1_STATE1_10_i_0\, B => 
        \I3.TCNT_n1_adt_net_137059_\, C => \I3.N_1966_1\, Y => 
        \I3.TCNT_n1\);
    
    \I3.un201_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_639\, Y => 
        \I3.un201_reg_ads_0_a2_0_a3_net_1\);
    
    \I3.PULSE_46_0_iv_0_il0r\ : AO21
      port map(A => \I3.REGMAPl4r_net_1\, B => 
        \I3.N_1906_i_0_0_adt_net_855640__net_1\, C => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854912__net_1\, Y
         => \I3.N_116_adt_net_134828_\);
    
    \I2.DTO_16_1_IV_0_0L29R_1071\ : AND2
      port map(A => \I2.N_182_ADT_NET_1007__385\, B => 
        \I2.DT_SRAMl29r_net_1\, Y => 
        \I2.DTO_16_1l29r_adt_net_28730_\);
    
    \I1.SSTATEL0R_3001\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_ns_il10r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL0R_755\);
    
    \I2.FCNTl0r_1136\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_947_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.FCNT_C0_398\);
    
    \I1.REG_74_0_IVL165R_2069\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l165r_adt_net_133665_\);
    
    \I2.TDCl3r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TDC_653_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TDCl3r_net_1\);
    
    \I2.DTE_1l23r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l23r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l23r_Rd1__net_1\);
    
    \I2.RAMAD1l15r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_669_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l15r_net_1\);
    
    \I2.G_EVNT_NUMl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_930_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl4r_net_1\);
    
    \I1.ISCK_0_sqmuxa_0_0_a2_1234\ : NAND3FFT
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__861\, B => 
        \I1.N_359\, C => \I1.sstatel4r_net_1\, Y => 
        \I1.N_656_496\);
    
    \I2.L1AF2_i\ : INV
      port map(A => \I2.L1AF2_net_1\, Y => \I2.L1AF2_i_net_1\);
    
    \I2.CRC32_12_0_0_x2l22r\ : XOR2FT
      port map(A => \I2.CRC32l22r_net_1\, B => \I2.N_4268_i_i\, Y
         => \I2.N_130_i_0_i_0\);
    
    \I2.CRC32_12_i_m2l16r\ : MUX2L
      port map(A => \I2.DT_TEMPl16r_net_1\, B => 
        \I2.DT_SRAMl16r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854196__net_1\, Y => 
        \I2.N_3961_i_i\);
    
    \I2.MSERCLKF1\ : DFFC
      port map(CLK => CLK_c, D => MSERCLK_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.MSERCLKF1_net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_45406_\ : OR3
      port map(A => \I2.STATE1_i_0_il16r\, B => 
        \I2.STATE1l2r_net_1\, C => 
        \I2.un1_STATE1_40_1_adt_net_45405__net_1\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45406__net_1\);
    
    \I2.ROFFSET_909\ : MUX2H
      port map(A => \I2.ROFFSETl9r_net_1\, B => 
        \I2.ROFFSET_n9_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_909_net_1\);
    
    \I3.STATE1_tr24_i_0_a3_28_tz\ : OR3FFT
      port map(A => \I3.N_58_i_0\, B => 
        \I3.un1_REGMAP_30_0_a2_0_net_1\, C => 
        \I3.N_178_adt_net_134608__net_1\, Y => 
        \I3.STATE1_tr24_i_0_a3_28_tz_i\);
    
    \I1.SSTATE_NS_1_IV_0_IL8R_1766\ : AO21
      port map(A => \I1.sstatel4r_net_1\, B => \I1.N_359\, C => 
        \I1.sstate_ns_1_iv_0_i_a4_2_il8r\, Y => 
        \I1.N_289_adt_net_107403_\);
    
    \I2.PIPE1_DT_12l5r\ : MUX2L
      port map(A => \I2.TDCDASl5r_net_1\, B => 
        \I2.TDCDASl3r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, Y
         => \I2.PIPE1_DT_12l5r_net_1\);
    
    \I3.REGMAPl51r\ : DFF
      port map(CLK => CLK_c, D => \I3.un7_ronly_0_a2_0_a3_net_1\, 
        Q => \I3.REGMAPl51r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I181_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl11r_net_1\, Y => 
        \I2.ADD_21x21_fast_I181_Y_0\);
    
    \I1.REG_1_211\ : MUX2H
      port map(A => \REGl310r\, B => \I1.REG_74l310r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_211_net_1\);
    
    \I2.PIPE10_DT_618\ : MUX2L
      port map(A => \I2.PIPE10_DTl13r_net_1\, B => \I2.N_3799\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_618_net_1\);
    
    \I2.L2TYPE_4_i_o2_1l14r\ : NOR2FT
      port map(A => \I2.L2ARRl1r_net_1\, B => \I2.L2ARRl0r_net_1\, 
        Y => \I2.N_4456\);
    
    \I3.VDBOFFB_30_IV_0L2R_2441\ : AND2
      port map(A => \REGl287r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162706_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I187_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_800\, B => 
        \I2.PIPE4_DTl17r_net_1\, Y => 
        \I2.ADD_21x21_fast_I187_Y_0_0\);
    
    \I2.PIPE4_DTL6R_3089\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL6R_853\);
    
    \I3.VDBOFFA_31_IV_0L0R_2632\ : AO21
      port map(A => \REGl181r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.VDBoffa_31l0r_adt_net_164638_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164645_\);
    
    \I2.TOKINBi\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKINBi_326_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => TOKINB_c);
    
    \I3.VDBi_29_0_a2l9r\ : OR2FT
      port map(A => \I3.REGMAPL7R_460\, B => \I3.N_1907_265\, Y
         => \I3.N_2033\);
    
    \I3.VDBoffal1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_45_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal1r_net_1\);
    
    \I1.REG_74_0_IVL346R_1867\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l346r_adt_net_116498_\);
    
    \I3.REG_1l98r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_279_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl98r\);
    
    \I2.STATE2_NS_I_0_O2_0_0_M7_I_1004\ : AO21FTT
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__890\, B => 
        \I2.END_EVNT2_619\, C => \I2.N_4273_adt_net_20927_\, Y
         => \I2.N_4273_adt_net_20928_\);
    
    \I2.PIPE8_DT_21_I_1L28R_1674\ : NOR3
      port map(A => \I2.NWPIPE7_689\, B => 
        \I2.N_565_0_adt_net_855728__net_1\, C => 
        \I2.PIPE8_DTl28r_net_1\, Y => 
        \I2.PIPE8_DT_21_i_1l28r_adt_net_82871_\);
    
    \I2.SUB8l19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_522_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l19r_net_1\);
    
    \I1.REG_74_0_ivl385r\ : AO21
      port map(A => \REGl385r\, B => \I1.N_257\, C => 
        \I1.REG_74l385r_adt_net_111577_\, Y => \I1.REG_74l385r\);
    
    \I1.REG_23_SQMUXA_0_A2_M2_E_2_1815\ : AND2FT
      port map(A => \I1.PAGECNT_319_net_1\, B => 
        \I1.PAGECNT_320_adt_net_854872__net_1\, Y => 
        \I1.REG_74_9_0_o4_a0_2l372r_adt_net_112100_Ra1_\);
    
    \I5.COMMAND_4l9r\ : MUX2L
      port map(A => \I5.AIR_WDATAl9r_net_1\, B => REGl110r, S => 
        REGl7r, Y => \I5.COMMAND_4l9r_net_1\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854624_\ : BFR
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854628__net_1\, 
        Y => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854624__net_1\);
    
    \I2.DT_TEMP_761\ : MUX2H
      port map(A => \I2.DT_TEMPl0r_net_1\, B => 
        \I2.DT_TEMP_7l0r_net_1\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.DT_TEMP_761_net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2430\ : AO21
      port map(A => \REGl296r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l3r_adt_net_162516_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162551_\);
    
    \I2.PIPE10_DT_614\ : MUX2L
      port map(A => \I2.PIPE10_DTl9r_net_1\, B => 
        \I2.PIPE9_DTl9r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_614_net_1\);
    
    \I2.DTE_cl_0_sqmuxa_2_adt_net_20059_\ : OR3FTT
      port map(A => \I2.STATE2L5R_507\, B => \I2.ENDF_401\, C => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20049__net_1\, Y => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20059__net_1\);
    
    \I2.PIPE5_DT_6_dl19r\ : MUX2L
      port map(A => \I2.PIPE4_DTl19r_net_1\, B => 
        \I2.un27_pipe5_dt1l19r\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855616__net_1\, Y => 
        \I2.PIPE5_DT_6_dl19r_net_1\);
    
    \I1.REG_21_sqmuxa_adt_net_855496_\ : BFR
      port map(A => \I1.REG_21_sqmuxa\, Y => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\);
    
    \I3.un2_vsel_2_i_0\ : OR2
      port map(A => \I3.ASBS_net_1\, B => 
        \I3.N_1510_adt_net_135035_\, Y => \I3.N_1510\);
    
    \I3.REG_1_150\ : MUX2L
      port map(A => VDB_inl1r, B => REGl49r, S => 
        \I3.N_1935_adt_net_855332__net_1\, Y => \I3.REG_1_150_0\);
    
    \I2.STATE1l11r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl7r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE1l11r_net_1\);
    
    \I2.PIPE4_DTL6R_3090\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL6R_854\);
    
    \I1.sstatel3r_1606\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl7r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL3R_713\);
    
    \I2.RAMAD_4l9r\ : MUX2L
      port map(A => \I2.N_536\, B => 
        \I1.PAGECNTl1r_adt_net_834904_Rd1__net_1\, S => LOAD_RES, 
        Y => \I2.RAMAD_4l9r_net_1\);
    
    \I2.NWPIPE2\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE1_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE2_net_1\);
    
    \I3.VDBOFFB_30_IV_0L6R_2370\ : AND2
      port map(A => \REGl379r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161950_\);
    
    \I1.REG_1_135\ : MUX2H
      port map(A => \REGl234r\, B => \I1.REG_74l234r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\, Y => 
        \I1.REG_1_135_net_1\);
    
    \I3.REG_44_i_0_m3l83r\ : MUX2H
      port map(A => VDB_inl0r, B => REGl83r, S => \I3.N_98\, Y
         => \I3.N_327\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I4_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L11R_441\, B => 
        \I2.PIPE4_DTL4R_477\, Y => \I2.N_64_0\);
    
    \I2.ADE_4l14r\ : MUX2L
      port map(A => \I2.RPAGEl14r\, B => \I2.WPAGEl14r_net_1\, S
         => NOESRAME_c, Y => \I2.ADE_4l14r_net_1\);
    
    \I1.N_268_Rd1__adt_net_854800_\ : BFR
      port map(A => \I1.N_268_Rd1__net_1\, Y => 
        \I1.N_268_Rd1__adt_net_854800__net_1\);
    
    \I3.TCNT_384\ : MUX2H
      port map(A => \I3.TCNTl0r_net_1\, B => \I3.TCNT_n0\, S => 
        \I3.TCNTe\, Y => \I3.TCNT_384_net_1\);
    
    \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854912_\ : BFR
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__831\, Y => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854912__net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_45413_\ : OR3
      port map(A => \I2.un1_STATE1_40_1_adt_net_45410__net_1\, B
         => \I2.un1_STATE1_40_1_adt_net_45389__net_1\, C => 
        \I2.un1_STATE1_40_1_adt_net_45408__net_1\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45413__net_1\);
    
    \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__2908\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_320_adt_net_854876__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__362\);
    
    \I2.N477_adt_net_302171_\ : NOR3FFT
      port map(A => \I2.N299_0\, B => \I2.N346_0_542\, C => 
        \I2.N353\, Y => \I2.N477_adt_net_302171__net_1\);
    
    \I2.L2TYPE_4_IL10R_1624\ : AND2
      port map(A => \I2.L2TYPEl10r_net_1\, B => 
        \I2.N_4442_adt_net_67433_\, Y => 
        \I2.N_4442_adt_net_67476_\);
    
    \I2.PIPE7_DTL27R_2789\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_82\);
    
    \I2.UN1_REG80_I_1701\ : NOR3FTT
      port map(A => \I2.N_3824_adt_net_90285_\, B => REGl46r, C
         => REGl35r, Y => \I2.N_3824_adt_net_90293_\);
    
    \I2.PIPE1_DT_42_1_IVL22R_1380\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855032__net_1\, 
        B => \I2.TDCDASl22r_net_1\, Y => 
        \I2.PIPE1_DT_42l22r_adt_net_46749_\);
    
    \I2.DTE_21_1_IV_0_0_18_M7_1216\ : AND2
      port map(A => \I2.DT_TEMPl18r_net_1\, B => \I2.N_4038_233\, 
        Y => \I2.DTE_21_1_iv_0_18_N_8_i_0_adt_net_35893_\);
    
    \I3.PULSE_332\ : AO21
      port map(A => \I3.N_311_adt_net_854748__net_1\, B => 
        \I3.N_122_adt_net_147352_\, C => 
        \I3.PULSE_332_adt_net_147433_\, Y => \I3.PULSE_332_net_1\);
    
    \I2.OFFSET_37_24l2r\ : MUX2L
      port map(A => \I2.N_813\, B => \I2.N_805\, S => 
        \I2.PIPE7_DTL26R_359\, Y => \I2.N_821\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854432_\ : BFR
      port map(A => \I2.N_4667_1_adt_net_1046__net_1\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854432__net_1\);
    
    \I1.REG_1_137\ : MUX2H
      port map(A => \REGl236r\, B => \I1.REG_74l236r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\, Y
         => \I1.REG_1_137_net_1\);
    
    \I3.TCNT_n3_0_0\ : AO21FTF
      port map(A => \I3.un1_STATE1_10_i_0\, B => 
        \I3.TCNT_n3_adt_net_137329_\, C => \I3.N_1966_1\, Y => 
        \I3.TCNT_n3\);
    
    \I2.L2AS_adt_net_855720_\ : BFR
      port map(A => \I2.L2AS_net_1\, Y => 
        \I2.L2AS_adt_net_855720__net_1\);
    
    \I2.REG_1_c0_i_a2_0\ : NAND2FT
      port map(A => REGL32R_388, B => \I2.N_119\, Y => \I2.N_121\);
    
    \I3.PIPEA_8l29r\ : OR2FT
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854484__net_1\, B => 
        \I3.N_238\, Y => \I3.PIPEA_8l29r_net_1\);
    
    \I2.un1_END_CHAINA1_0_sqmuxa_i_o3\ : AO21FTT
      port map(A => \I2.N_3870\, B => \I2.N_3347_1\, C => 
        \I2.N_3281_adt_net_53327_\, Y => \I2.N_3281\);
    
    \I1.REG_1_111\ : MUX2H
      port map(A => \REGl210r\, B => \I1.N_1349\, S => 
        \I1.N_50_0_ADT_NET_1409__320\, Y => \I1.REG_1_111_net_1\);
    
    \I2.DT_SRAMl11r\ : MUX2L
      port map(A => \I2.N_879\, B => \I2.PIPE2_DTl11r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672__net_1\, 
        Y => \I2.DT_SRAMl11r_net_1\);
    
    \I2.PIPE1_DT_12l3r\ : MUX2L
      port map(A => \I2.TDCDASl3r_net_1\, B => 
        \I2.TDCDASl1r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092__net_1\, Y
         => \I2.PIPE1_DT_12l3r_net_1\);
    
    \I3.DSS_0\ : DFFS
      port map(CLK => CLK_c, D => \I3.DSSF1_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.DSS_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I154_Y_0_O2_2694\ : AO21
      port map(A => \I2.N_33_adt_net_55020_\, B => 
        \I2.N_147_0_adt_net_604832_\, C => 
        \I2.N_82_adt_net_496796_\, Y => \I2.N_82\);
    
    \I2.DTE_21_1_IV_0_0L17R_1223\ : AND3FTT
      port map(A => 
        \I2.REG_0l3r_adt_net_848__adt_net_854216__net_1\, B => 
        \I2.STATE2l1r_adt_net_855124__net_1\, C => REGl28r, Y => 
        \I2.DTE_21_1l17r_adt_net_36146_\);
    
    \I2.PIPE1_DT_738\ : MUX2L
      port map(A => \I2.PIPE1_DTl11r_net_1\, B => 
        \I2.PIPE1_DT_42l11r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854580__net_1\, 
        Y => \I2.PIPE1_DT_738_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I188_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl18r_net_1\, Y => 
        \I2.ADD_21x21_fast_I188_Y_0\);
    
    AMB_padl3r : IB33
      port map(PAD => AMB(3), Y => AMB_cl3r);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I13_P0N_i_a4\ : OR2
      port map(A => \I2.RAMDT4L5R_821\, B => 
        \I2.PIPE4_DTl13r_net_1\, Y => \I2.N_92\);
    
    \I5.REG_1_22\ : MUX2H
      port map(A => \I5.TEMPDATAl3r_net_1\, B => REGl439r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855876__net_1\, Y
         => \I5.REG_1_22_net_1\);
    
    \I2.ROFFSETe_0_adt_net_1030_\ : AO21FTT
      port map(A => \I2.N_3012\, B => 
        \I2.N_12254_i_adt_net_24491_\, C => 
        \I2.ROFFSETe_0_adt_net_27187__net_1\, Y => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\);
    
    \I2.FID_416\ : MUX2H
      port map(A => FID_cl0r, B => \I2.FID_7l0r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        Y => \I2.FID_416_net_1\);
    
    \I1.REG_1_76\ : MUX2H
      port map(A => \REGl175r\, B => \I1.REG_74l175r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\, Y => 
        \I1.REG_1_76_net_1\);
    
    \I1.REG_74_0_ivl351r\ : AO21
      port map(A => \REGl351r\, B => \I1.N_225\, C => 
        \I1.REG_74l351r_adt_net_116031_\, Y => \I1.REG_74l351r\);
    
    REGl394r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_295_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl394r\);
    
    \I2.CRC32_12_i_0_m2l7r\ : MUX2H
      port map(A => \I2.DT_SRAMl7r_net_1\, B => 
        \I2.DT_TEMPl7r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854436__net_1\, Y => 
        \I2.N_226_i_i\);
    
    \I3.RAMAD_VMEl9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_33_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl9r);
    
    \I2.END_TDC1_1_sqmuxa_i_o2\ : OR2
      port map(A => \I2.N_3887_adt_net_21857_\, B => 
        \I2.N_3887_adt_net_21865_\, Y => \I2.N_3887\);
    
    \I3.VDBi_358\ : MUX2L
      port map(A => \I3.VDBil18r_net_1\, B => \I3.VDBi_57l18r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_358_net_1\);
    
    ADE_padl1r : OB33PH
      port map(PAD => ADE(1), A => ADE_cl1r);
    
    \I2.DTO_16_1l22r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l22r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l22r_Rd1__net_1\);
    
    \I2.PIPE1_DT_753\ : MUX2L
      port map(A => \I2.PIPE1_DTl26r_net_1\, B => 
        \I2.PIPE1_DT_42_1_iv_i_0l26r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854564__net_1\, 
        Y => \I2.PIPE1_DT_753_net_1\);
    
    \I2.SRAM_EVNT_n2_0\ : XOR2FT
      port map(A => \I2.SRAM_EVNTl2r_net_1\, B => \I2.N_128_1\, Y
         => \I2.SRAM_EVNT_n2_0_net_1\);
    
    \I2.G_EVNT_NUM_n6_i_o2_0_1289\ : AND2
      port map(A => \I2.N_4672_553\, B => 
        \I2.G_EVNT_NUMl6r_net_1\, Y => \I2.N_198_551\);
    
    \I1.REG_1_128\ : MUX2H
      port map(A => \REGl227r\, B => \I1.REG_74l227r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855432__net_1\, Y => 
        \I1.REG_1_128_net_1\);
    
    \I3.STATE2_0_sqmuxa_2_i_o3\ : NAND2FT
      port map(A => \I3.DSS_net_1\, B => \I3.N_258\, Y => 
        \I3.N_281\);
    
    \I2.SUB8_522\ : AND2
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855160__net_1\, B
         => \I2.SUB_21x21_fast_I215_Y_0\, Y => 
        \I2.SUB8_522_adt_net_551987_\);
    
    REGl249r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_150_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl249r\);
    
    \I1.REG_1_289\ : MUX2H
      port map(A => \REGl388r\, B => \I1.REG_74l388r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y
         => \I1.REG_1_289_net_1\);
    
    \I2.PIPE4_DTL9R_2954\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL9R_471\);
    
    \I2.EVNT_REJ_2_SQMUXA_1059\ : NOR3FFT
      port map(A => REGl1r, B => 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26947_\, C => REGl2r, Y => 
        \I2.EVNT_REJ_2_sqmuxa_adt_net_26950_\);
    
    \I2.FIDl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_446\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl30r);
    
    \I2.TRGSERV_2_I_1\ : AND2
      port map(A => \I2.TRGSERVl0r_net_1\, B => 
        \I2.STATE1_i_0_il15r\, Y => \I2.DWACT_ADD_CI_0_TMP_0l0r\);
    
    \I2.STATE1_ns_il8r\ : OA21
      port map(A => \I2.N_3272\, B => \I2.N_3870\, C => 
        \I2.N_3316\, Y => \I2.N_3206_i_0\);
    
    \I3.REG_1_161\ : MUX2L
      port map(A => VDB_inl12r, B => REGl60r, S => 
        \I3.N_1935_adt_net_855328__net_1\, Y => \I3.REG_1_161_0\);
    
    \I2.PIPE4_DTl7r_adt_net_854552__adt_net_854948_\ : BFR
      port map(A => \I2.PIPE4_DTL7R_481\, Y => 
        \I2.PIPE4_DTl7r_adt_net_854552__adt_net_854948__net_1\);
    
    \I1.PAGECNTl8r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_319_adt_net_854860__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTl8r_net_1\);
    
    \I2.N_182_ADT_NET_1007__2914\ : OR2
      port map(A => \I2.STATE2L0R_588\, B => 
        \I2.STATE2_nsl2r_adt_net_24911_\, Y => 
        \I2.N_182_ADT_NET_1007__385\);
    
    \I4.bcnt_5\ : MUX2H
      port map(A => \I4.bcntl0r_net_1\, B => \I4.bcnt_3l0r_net_1\, 
        S => \I4.STATE1l1r_net_1\, Y => \I4.bcnt_5_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I146_Y\ : AO21
      port map(A => \I2.N323_0\, B => \I2.N510_adt_net_220925_\, 
        C => \I2.N322\, Y => \I2.N516\);
    
    \I2.FIRST_TDC\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.FIRST_TDC_675_net_1\, 
        SET => CLEAR_STAT_i_0, Q => \I2.FIRST_TDC_i_0_i\);
    
    \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855088_\ : BFR
      port map(A => \I2.un2_tdcgdb1_0_adt_net_830__net_1\, Y => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855088__net_1\);
    
    \I2.un1_tdc_res_46_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl410r, Y => 
        \I2.N_4627_i_0\);
    
    \I2.PIPE5_DT_686\ : MUX2L
      port map(A => \I2.PIPE5_DTl10r_net_1\, B => 
        \I2.PIPE5_DT_6l10r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_686_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I165_Y_1687\ : AND2FT
      port map(A => \I2.N311_0\, B => \I2.N315\, Y => 
        \I2.N498_1_adt_net_88035_\);
    
    \I1.REG_74_0_IV_0L262R_1961\ : AND2
      port map(A => \REGl262r\, B => 
        \I1.N_137_adt_net_854764__net_1\, Y => 
        \I1.REG_74l262r_adt_net_124543_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I140_Y_0_o2\ : OA21FTT
      port map(A => \I2.N_128_135\, B => 
        \I2.N_70_adt_net_255802__net_1\, C => \I2.N_112_2\, Y => 
        \I2.N_70\);
    
    \I1.BYTECNTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_306_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BYTECNTl8r_net_1\);
    
    \I2.ROFFSET_913\ : MUX2H
      port map(A => \I2.ROFFSETl5r_net_1\, B => 
        \I2.ROFFSET_n5_net_1\, S => 
        \I2.ROFFSETe_0_adt_net_1030__net_1\, Y => 
        \I2.ROFFSET_913_net_1\);
    
    \I2.ERR_WORDS_RDY\ : DFFC
      port map(CLK => CLK_c, D => \I2.ERR_WORDS_RDY_415_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.ERR_WORDS_RDY_net_1\);
    
    \I1.REG_3_sqmuxa_0_a2_0_816\ : NAND2FT
      port map(A => \I1.PAGECNTL9R_245\, B => \I1.N_238_RD1__313\, 
        Y => \I1.N_254_194\);
    
    \I1.REG_74_0_IVL266R_1957\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, Y => 
        \I1.REG_74l266r_adt_net_124199_\);
    
    \I2.SUB8l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_507_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l4r_net_1\);
    
    \I3.VDBi_361\ : MUX2L
      port map(A => \I3.VDBil21r_net_1\, B => \I3.VDBi_57l21r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__115\, Y => 
        \I3.VDBi_361_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL11R_1456\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl7r\, Y => 
        \I2.PIPE1_DT_42l11r_adt_net_49695_\);
    
    \I2.N_4244_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4244\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4244_Rd1__net_1\);
    
    \I2.TRGCNT_c1_i_o2\ : AND2
      port map(A => \I2.TRGCNTl0r_net_1\, B => 
        \I2.TRGCNT_i_0_il1r\, Y => \I2.N_3765\);
    
    \I2.LSRAM_INl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_411_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl27r_net_1\);
    
    \I1.REG_74_0_ivl168r\ : AO21
      port map(A => \REGl168r\, B => \I1.N_41\, C => 
        \I1.REG_74l168r_adt_net_133407_\, Y => \I1.REG_74l168r\);
    
    \I2.FID_7_IVL2R_1731\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl2r_net_1\, 
        C => \I2.FID_7l2r_adt_net_93351_\, Y => 
        \I2.FID_7l2r_adt_net_93359_\);
    
    \I2.EVNT_REJ_646\ : MUX2L
      port map(A => \I2.EVNT_REJ_2_sqmuxa_net_1\, B => 
        \I2.EVNT_REJ_net_1\, S => \I2.STATE3l5r_net_1\, Y => 
        \I2.EVNT_REJ_646_net_1\);
    
    \I2.OFFSET_37_8l7r\ : MUX2L
      port map(A => \REGl364r\, B => \REGl300r\, S => 
        \I2.PIPE7_DTL27R_67\, Y => \I2.N_698\);
    
    \I2.ADOl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl0r);
    
    \I3.un231_reg_ads_0_a2_4_a3_1\ : NAND3FFT
      port map(A => \I3.VASl12r_net_1\, B => \I3.N_555\, C => 
        \I3.VASl2r_net_1\, Y => \I3.un231_reg_ads_1\);
    
    \I1.REG_1_133\ : MUX2H
      port map(A => \REGl232r\, B => \I1.REG_74l232r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\, Y => 
        \I1.REG_1_133_net_1\);
    
    \I2.SUB8l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_504_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l1r_net_1\);
    
    \I3.REG_1l84r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_265_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl84r);
    
    \I2.PIPE1_DTl8r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_735_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl8r_net_1\);
    
    \I2.LEAD_FLAG6_639_1604\ : NOR2FT
      port map(A => LEAD_FLAGl2r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_639_adt_net_64404_\);
    
    \I2.OFFSET_37_16l0r\ : MUX2L
      port map(A => \REGl261r\, B => \REGl197r\, S => 
        \I2.PIPE7_DTL27R_86\, Y => \I2.N_755\);
    
    REGl341r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_242_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl341r\);
    
    \I3.REG_1l134r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_182_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl134r\);
    
    \I2.DT_TEMP_769\ : MUX2H
      port map(A => \I2.DT_TEMPl8r_net_1\, B => 
        \I2.DT_TEMP_7l8r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_769_net_1\);
    
    \I1.PAGECNT_n6_i_i_a2_852\ : AND2FT
      port map(A => \I1.PAGECNTL6R_836\, B => \I1.PAGECNTL5R_310\, 
        Y => \I1.N_590_230\);
    
    \I3.TCNT3l1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT3_378_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT3l1r_net_1\);
    
    \I2.RAMADl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l14r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl14r);
    
    \I1.REG_74_0_iv_0l225r\ : AO21
      port map(A => \FBOUTl4r\, B => \I1.N_12233_i\, C => 
        \I1.REG_74l225r_adt_net_128222_\, Y => \I1.REG_74l225r\);
    
    DTE_padl19r : IOB33PH
      port map(PAD => DTE(19), A => \I2.DTE_1l19r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl19r);
    
    \I3.STATE1_illegalpipe2\ : DFFLS
      port map(CLK => CLK_c, D => \I3.N_1309_i_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.N_1310_i_0\);
    
    \I3.un224_reg_ads_0_a2_3_a2\ : NAND2
      port map(A => \I3.LWORDS_788\, B => \I3.N_545\, Y => 
        \I3.N_546\);
    
    \I3.PIPEAl11r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_242_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl11r_net_1\);
    
    \I3.un91_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_583\, B => \I3.N_551\, Y => 
        \I3.un91_reg_ads_0_a2_0_a3_net_1\);
    
    ADO_padl8r : OB33PH
      port map(PAD => ADO(8), A => ADO_cl8r);
    
    \I1.REG_74_0_IVL189R_2045\ : AND2
      port map(A => \FBOUTl0r\, B => \I1.REG_4_sqmuxa\, Y => 
        \I1.REG_74l189r_adt_net_131527_\);
    
    \I1.REG_1_286\ : MUX2H
      port map(A => \REGl385r\, B => \I1.REG_74l385r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y => 
        \I1.REG_1_286_net_1\);
    
    \I2.PIPE5_DTl30r_1514\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_706_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTL30R_621\);
    
    \I1.sstate_ns_0_iv_0_0_o2l2r_854\ : OR2
      port map(A => \I1.N_317_Rd1__net_1\, B => 
        \I1.N_321_adt_net_105403_\, Y => \I1.N_321_232\);
    
    \I2.REG_1_C11_I_1738\ : AND2FT
      port map(A => REGl43r, B => \I2.N_131\, Y => 
        \I2.N_3840_adt_net_101218_\);
    
    \I1.REG_74_0_IV_0L362R_1845\ : AND2
      port map(A => \FBOUTl5r\, B => \I1.REG_25_sqmuxa\, Y => 
        \I1.REG_74l362r_adt_net_114697_\);
    
    \I2.SRAM_FULL_1486\ : DFFC
      port map(CLK => CLK_c, D => \I2.SRAM_FULL_488_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.SRAM_FULL_593\);
    
    \I1.REG_1_89\ : MUX2H
      port map(A => \REGl188r\, B => \I1.REG_74l188r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, Y
         => \I1.REG_1_89_net_1\);
    
    \I2.DTE_1_854\ : MUX2L
      port map(A => \I2.DTE_1l14r_Rd1__net_1\, B => 
        \I2.DTE_21_1l14r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\, Y => 
        \I2.DTE_1l14r\);
    
    \I3.VDBOFFA_31_IV_0L0R_2633\ : OR2
      port map(A => \I3.VDBoffa_31l0r_adt_net_164641_\, B => 
        \I3.VDBoffa_31l0r_adt_net_164642_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164647_\);
    
    \I2.FIDl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_424_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl8r);
    
    \I3.VDBml26r\ : MUX2L
      port map(A => \I3.VDBil26r_net_1\, B => \I3.N_168\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml26r_net_1\);
    
    \I3.REG1_134\ : MUX2L
      port map(A => VDB_inl1r, B => \I3.REG1l1r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG1_134_net_1\);
    
    \I2.OFFSET_37_7l3r\ : MUX2L
      port map(A => \I2.N_678\, B => \I2.N_654\, S => 
        \I2.PIPE7_DTL25R_682\, Y => \I2.N_686\);
    
    \I2.OFFSETl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_563_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETl3r_net_1\);
    
    \I2.EVNT_NUM_n10_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl10r_net_1\, B => 
        \I2.EVNT_NUM_c9_net_1\, Y => \I2.EVNT_NUM_n10_tz_i\);
    
    \I3.VDBoff_123\ : MUX2L
      port map(A => \I3.VDBoffl7r_net_1\, B => \I3.N_81\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_123_net_1\);
    
    \I1.N_113_adt_net_3714_\ : OR2
      port map(A => \I1.N_41_9\, B => 
        \I1.N_113_adt_net_126306__net_1\, Y => 
        \I1.N_113_adt_net_3714__net_1\);
    
    \I3.REG_44_IL88R_2303\ : AOI21FTT
      port map(A => REGl88r, B => \I3.N_98_0\, C => \I3.N_1671\, 
        Y => \I3.N_1634_adt_net_150223_\);
    
    \I2.un2_evnt_word_I_38\ : XOR2
      port map(A => \I2.WOFFSETl7r\, B => \I2.N_29\, Y => 
        \I2.I_38\);
    
    \I3.PIPEB_104_2319\ : NOR2FT
      port map(A => \I3.PIPEBl25r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_104_adt_net_159663_\);
    
    FID_padl13r : OB33PH
      port map(PAD => FID(13), A => FID_cl13r);
    
    \I2.N_4252_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4252\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4252_Rd1__net_1\);
    
    \I1.REG_1_sqmuxa_0_a2_1\ : OR2
      port map(A => \I1.PAGECNTL5R_311\, B => 
        \I1.N_237_adt_net_854804__net_1\, Y => \I1.N_255\);
    
    \I1.REG_74_0_IVL330R_1886\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l330r_adt_net_118088_\);
    
    \I4.STATE1_nsl0r\ : AO21FTT
      port map(A => END_TDC, B => \I4.STATE1l2r_net_1\, C => 
        \I4.STATE1l0r_net_1\, Y => \I4.STATE1_nsl0r_net_1\);
    
    \I2.PIPE2_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl2r_net_1\);
    
    \I2.LEAD_FLAG6_641_1602\ : NOR2FT
      port map(A => LEAD_FLAGl4r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_641_adt_net_64180_\);
    
    \I2.DT_SRAM_0l7r\ : MUX2L
      port map(A => \I2.PIPE10_DTl7r_net_1\, B => 
        \I2.PIPE5_DTl7r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, Y => 
        \I2.N_875\);
    
    \I2.DT_TEMP_7l6r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, B => 
        \I2.DT_SRAMl6r_net_1\, Y => \I2.DT_TEMP_7l6r_net_1\);
    
    \I1.REG_1_136\ : MUX2H
      port map(A => \REGl235r\, B => \I1.REG_74l235r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\, Y => 
        \I1.REG_1_136_net_1\);
    
    \I2.PIPE10_DT_17_i_0l15r\ : OAI21TTF
      port map(A => \I2.N_22_i_0_adt_net_855596__net_1\, B => 
        \I2.PIPE9_DTl15r_net_1\, C => \I2.N_26\, Y => 
        \I2.PIPE10_DT_17_i_0l15r_net_1\);
    
    \I1.REG_0_sqmuxa_i_0_a4_1_907\ : NAND2
      port map(A => \I1.N_598_23\, B => 
        \I1.sstate_ns_il5r_adt_net_107266_\, Y => 
        \I1.N_435_1_285\);
    
    REGl335r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_236_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl335r\);
    
    \I2.TDCGDBi_0_sqmuxa_i_o2\ : NOR2
      port map(A => \I2.CHAINB_EN244_c_0_adt_net_855240__net_1\, 
        B => \I2.N_3879_180\, Y => \I2.N_3883\);
    
    \I1.LUT_0_sqmuxa_i_0\ : OAI21FTF
      port map(A => \I1.sstatel4r_net_1\, B => \I1.N_359\, C => 
        \I1.N_1384\, Y => \I1.N_56\);
    
    \I3.REGMAPl13r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un54_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPl13r_net_1\);
    
    \I3.VDBi_57l7r_adt_net_143037_\ : AO21FTT
      port map(A => \I3.N_2017\, B => 
        \I3.VDBi_57l7r_adt_net_3750__net_1\, C => 
        \I3.VDBi_57l7r_adt_net_143023__net_1\, Y => 
        \I3.VDBi_57l7r_adt_net_143037__net_1\);
    
    \I2.PIPE1_DTl5r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_732_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl5r_net_1\);
    
    \I2.EVNT_WORDl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_721_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl8r_net_1\);
    
    REGl340r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_241_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl340r\);
    
    \I1.LOAD_RESi_50\ : OA21TTF
      port map(A => LOAD_RES, B => \I1.sstatel3r_net_1\, C => 
        \PULSEl0r_adt_net_854532__adt_net_855544__net_1\, Y => 
        \I1.LOAD_RESi_50_net_1\);
    
    REGl269r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_170_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl269r\);
    
    \I3.VDBi_57_iv_0_o3_i_o2l2r\ : NOR2
      port map(A => \I3.STATE1_IPL2R_886\, B => 
        \I3.STATE1_ipl3r_adt_net_854368__net_1\, Y => \I3.N_1904\);
    
    \I2.STATE1_NS_0L11R_1034\ : NOR2FT
      port map(A => \I2.STATE1L6R_630\, B => 
        \I2.END_CHAINB1_709_adt_net_2397__net_1\, Y => 
        \I2.STATE1_nsl11r_adt_net_23385_\);
    
    \I2.MIC_REG1l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_305_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1l4r_net_1\);
    
    \I1.REG_74_0_ivl392r\ : AO21
      port map(A => \REGl392r\, B => \I1.N_265\, C => 
        \I1.REG_74l392r_adt_net_110870_\, Y => \I1.REG_74l392r\);
    
    \I2.PIPE10_DT_17_0l30r\ : AO21
      port map(A => \I2.N_22_i_0_adt_net_855592__net_1\, B => 
        \I2.PIPE10_DT_17l29r\, C => \I2.PIPE9_DTl30r_net_1\, Y
         => \I2.PIPE10_DT_17l30r\);
    
    \I5.REG_1_17\ : MUX2H
      port map(A => REGl131r, B => REGl434r, S => 
        \I5.REG_2_sqmuxa_0_adt_net_975__adt_net_855872__net_1\, Y
         => \I5.REG_1_17_net_1\);
    
    \I1.PAGECNT_n2_0_0_x2\ : XOR2FT
      port map(A => \I1.PAGECNTl2r_adt_net_834908_Rd1__net_1\, B
         => \I1.N_300_Rd1__net_1\, Y => \I1.N_390_i_i_0_i\);
    
    \I2.DT_TEMP_7l8r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, B => 
        \I2.DT_SRAMl8r_net_1\, Y => \I2.DT_TEMP_7l8r_net_1\);
    
    \I2.PIPE4_DTl2r_1252_1753\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL2R_860\);
    
    \I1.REG_74L380R_1818\ : AND3FFT
      port map(A => \I1.REG_74_1_380_m8_i_0_Rd1__net_1\, B => 
        \I1.REG_74_1_380_N_15_i_i_i\, C => 
        \I1.REG_74_1_380_m8_i_0_0\, Y => 
        \I1.N_249_adt_net_112440_\);
    
    \I2.I_1337_ca_0_and2\ : NOR2FT
      port map(A => \I2.SUB8l5r_net_1\, B => \I2.OFFSETl2r_net_1\, 
        Y => \I2.N_3537_i_i\);
    
    \I2.STATE2_ns_0l1r\ : OR3FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855196__net_1\, 
        B => \I2.STATE2_nsl1r_adt_net_24963_\, C => 
        \I2.STATE2_nsl1r_adt_net_24965_\, Y => \I2.STATE2_nsl1r\);
    
    \I3.VDBOFFA_31_IV_0L3R_2571\ : AO21
      port map(A => \REGl200r\, B => \I3.REGMAPl22r_net_1\, C => 
        \I3.VDBoffa_31l3r_adt_net_164024_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164068_\);
    
    \I2.TDCDBSl15r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl15r, Q => 
        \I2.TDCDBSl15r_net_1\);
    
    DPR_padl21r : IB33
      port map(PAD => DPR(21), Y => DPR_cl21r);
    
    \I3.REG_1_i_il2r\ : AO21
      port map(A => \I3.REG3l2r_net_1\, B => \I3.REG2l2r_net_1\, 
        C => \REGl2r_adt_net_21315_\, Y => REGl2r);
    
    \I2.EVNT_NUMl1r_1135\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_962_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUML1R_397\);
    
    \I2.un1_tdc_res_26_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl410r, Y => 
        \I2.N_4607_i_0\);
    
    \I3.VDBOFFA_31_IV_0L4R_2557\ : AO21
      port map(A => \REGl257r\, B => \I3.REGMAPl29r_net_1\, C => 
        \I3.VDBoffa_31l4r_adt_net_163850_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163882_\);
    
    \I3.VDBI_57_0_IV_0L19R_2171\ : AND2FT
      port map(A => \I3.N_1917_adt_net_855336__net_1\, B => 
        \I3.REGl152r\, Y => \I3.VDBi_57l19r_adt_net_139383_\);
    
    \I3.PIPEA_8_0l6r\ : MUX2L
      port map(A => DPR_cl6r, B => \I3.PIPEA1l6r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855364__net_1\, Y => \I3.N_215\);
    
    \I3.STATE1_0l9r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl9r\);
    
    \I3.PIPEA1l17r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_315_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l17r_net_1\);
    
    \I2.PIPE3_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl30r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl30r_net_1\);
    
    \I3.PIPEA_8l21r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854464__net_1\, B => 
        \I3.N_230\, Y => \I3.PIPEA_8l21r_net_1\);
    
    \I3.VDBoffal5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_49_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal5r_net_1\);
    
    \I2.STATE1l5r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3214_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1l5r_net_1\);
    
    \I1.REG_74_0_ivl383r\ : AO21
      port map(A => \REGl383r\, B => \I1.N_257\, C => 
        \I1.REG_74l383r_adt_net_111749_\, Y => \I1.REG_74l383r\);
    
    \I2.BITCNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.BITCNT_940\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.BITCNT_c0\);
    
    \I3.STATE1_428_0\ : NAND2FT
      port map(A => \HWRES_3_ADT_NET_738__17\, B => 
        \I3.N_1310_i_0\, Y => \I3.N_1311_0\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I162_un1_Y\ : AND3FFT
      port map(A => \I2.N348\, B => \I2.N356\, C => \I2.N513\, Y
         => \I2.I162_un1_Y\);
    
    \I2.DTE_21_1_IV_0L20R_1261\ : OR3
      port map(A => \I2.DTO_16_1l20r_adt_net_30786_\, B => 
        \I2.DTE_21_1l20r_adt_net_37605_\, C => 
        \I2.DTE_21_1l20r_adt_net_37612_\, Y => 
        \I2.DTE_21_1l20r_adt_net_37614_\);
    
    \I2.N477_adt_net_302179_\ : AO21
      port map(A => \I2.N299_0\, B => \I2.N345\, C => 
        \I2.N477_adt_net_302171__net_1\, Y => 
        \I2.N477_adt_net_302179__net_1\);
    
    \I2.G_EVNT_NUMl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_932_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl2r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L4R_2559\ : AO21
      port map(A => \REGl273r\, B => \I3.REGMAPl31r_net_1\, C => 
        \I3.VDBoffa_31l4r_adt_net_163858_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163884_\);
    
    \I3.REG_1_I_IL1R_1005\ : OA21
      port map(A => \I3.REG3L1R_744\, B => \I3.REG2l1r_net_1\, C
         => \I3.REG1l1r_net_1\, Y => \REGl1r_adt_net_21137_\);
    
    \I3.REG_1_295\ : MUX2L
      port map(A => VDB_inl13r, B => REGl114r, S => 
        \I3.N_318_adt_net_855884__net_1\, Y => \I3.REG_1_295_0\);
    
    \I1.REG_23_sqmuxa_adt_net_855512_\ : BFR
      port map(A => \I1.REG_23_sqmuxa\, Y => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I182_Y\ : XOR2FT
      port map(A => \I2.N_42_1\, B => 
        \I2.ADD_21x21_fast_I182_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l12r\);
    
    \I2.DTO_16_1_iv_0_a2_2l21r_674\ : AND3
      port map(A => \I2.N_223_54\, B => \I2.N_4182\, C => 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_888__net_1\, Y => 
        \I2.N_196_52\);
    
    \I2.PIPE1_DT_12l2r\ : MUX2L
      port map(A => \I2.TDCDASl2r_net_1\, B => 
        \I2.TDCDASl0r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855092__net_1\, Y
         => \I2.PIPE1_DT_12l2r_net_1\);
    
    \I1.PAGECNTL9R_2975\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854856__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL9R_492\);
    
    \I0.CLEAR_936\ : NAND3FFT
      port map(A => \I0.CLEAR_adt_net_15816_\, B => PULSEl1r, C
         => LOAD_RES_1, Y => \I0.CLEAR_adt_net_15818_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I136_Y_0_o2_m4_2\ : AO21
      port map(A => \I2.RAMDT4L12R_827\, B => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_2_i_adt_net_271662_\, C
         => \I2.N_112_1\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_2_i_adt_net_56602_\);
    
    \I3.REG_0_sqmuxa_2_adt_net_855308_\ : BFR
      port map(A => \I3.REG_0_sqmuxa_2\, Y => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\);
    
    \I2.CRC32_12_i_x2l13r\ : XOR2FT
      port map(A => \I2.CRC32l13r_net_1\, B => \I2.N_3958_i_i\, Y
         => \I2.N_115_i_i_0\);
    
    \I2.DTO_16_1_IV_0L24R_1092\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855676__net_1\, B => 
        \I2.DTO_9l24r\, Y => \I2.DTO_16_1l24r_adt_net_29854_\);
    
    \I3.VDBI_57_0_IV_0_0L15R_2187\ : AO21
      port map(A => REGl47r, B => \I3.N_403_1\, C => 
        \I3.VDBi_57l15r_adt_net_139969_\, Y => 
        \I3.VDBi_57l15r_adt_net_139971_\);
    
    \I1.REG_1_288\ : MUX2H
      port map(A => \REGl387r\, B => \I1.REG_74l387r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855532__net_1\, Y => 
        \I1.REG_1_288_net_1\);
    
    \I2.PIPE6_DT_460\ : MUX2H
      port map(A => \I2.PIPE5_DTl6r_net_1\, B => 
        \I2.PIPE6_DTl6r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_460_net_1\);
    
    \I2.SUB8_510\ : MUX2H
      port map(A => \I2.SUB8l7r_net_1\, B => \I2.SUB8_2l7r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855148__net_1\, Y => 
        \I2.SUB8_510_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL13R_1443\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044__net_1\, 
        B => \I2.PIPE1_DT_12l13r_net_1\, Y => 
        \I2.PIPE1_DT_42l13r_adt_net_49195_\);
    
    \I1.REG_1_261\ : MUX2H
      port map(A => \REGl360r\, B => \I1.REG_74l360r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_261_net_1\);
    
    \I2.STATE1_ns_a3_i_o3l12r_801\ : NAND2
      port map(A => \I2.STATE1L7R_633\, B => 
        \I2.N_3883_adt_net_854632__net_1\, Y => \I2.N_3889_179\);
    
    \I2.ROFFSET_c7\ : NAND2
      port map(A => \I2.ROFFSETl7r_net_1\, B => 
        \I2.ROFFSET_c6_net_1\, Y => \I2.ROFFSET_c7_net_1\);
    
    \I3.VDBi_57_0_iv_0_a2_0_0_a2l19r\ : AND3FFT
      port map(A => \I3.N_1905_1_adt_net_855376__net_1\, B => 
        \I3.REGMAPl17r_adt_net_854292__net_1\, C => 
        \I3.REGMAPl9r_adt_net_854316__net_1\, Y => \I3.N_1839\);
    
    \I2.OFFSET_37_11l7r\ : MUX2L
      port map(A => \REGl380r\, B => \REGl316r\, S => 
        \I2.PIPE7_DTL27R_75\, Y => \I2.N_722\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I44_Y_1653\ : AO21
      port map(A => \I2.N_3537_i_i\, B => \I2.G_1_3\, C => 
        \I2.N_3539_i_i\, Y => \I2.N309_adt_net_70030_\);
    
    \I2.DTO_16_1_iv_0_a2_4_18_m7_0_a5\ : AND3
      port map(A => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, B => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        C => \I2.DTO_16_1_iv_0_a2_4_18_N_11\, Y => 
        \I2.DTO_16_1_iv_0_a2_4_18_N_12_i\);
    
    \I3.REG_1_211\ : MUX2L
      port map(A => VDB_inl30r, B => \I3.REGl163r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\, Y => 
        \I3.REG_1_211_0\);
    
    \I1.REG_74_0_ivl304r\ : AO21
      port map(A => \REGl304r\, B => \I1.N_177\, C => 
        \I1.REG_74l304r_adt_net_120524_\, Y => \I1.REG_74l304r\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2274\ : AND2
      port map(A => \I3.N_2045\, B => \I3.REGl91r\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146420_\);
    
    \I5.TEMPDATAl7r\ : DFFC
      port map(CLK => CLK_c, D => \I5.TEMPDATA_81_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.TEMPDATAl7r_net_1\);
    
    \I2.resyn_0_I2_FID_446\ : MUX2H
      port map(A => FID_cl30r, B => \I2.FID_7l30r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\, 
        Y => \I2.FID_446\);
    
    REGl361r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_262_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl361r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0\ : OR2
      port map(A => \I2.N_45_1\, B => \I2.N525_0_adt_net_58015_\, 
        Y => \I2.N525_0\);
    
    \I2.DT_TEMP_771\ : MUX2H
      port map(A => \I2.DT_TEMPl10r_net_1\, B => 
        \I2.DT_TEMP_7l10r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_771_net_1\);
    
    \I2.WOFFSET_13_il7r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_38\, Y => \I2.N_4250\);
    
    \I3.PIPEB_82\ : AO21
      port map(A => DPR_cl3r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_82_adt_net_160587_\, Y => 
        \I3.PIPEB_82_net_1\);
    
    \I2.END_CHAINB1_709_1536\ : NOR2FT
      port map(A => \I2.END_CHAINB1_net_1\, B => \I2.N_158\, Y
         => \I2.END_CHAINB1_709_adt_net_53455_\);
    
    \I1.REG_74_0_ivl170r\ : AO21
      port map(A => \REGl170r\, B => \I1.N_41\, C => 
        \I1.REG_74l170r_adt_net_133235_\, Y => \I1.REG_74l170r\);
    
    \I3.UN12_TCNT3_2641\ : NOR2
      port map(A => \I3.TCNT3_i_0_il6r_net_1\, B => 
        \I3.TCNT3l5r_net_1\, Y => \I3.un12_tcnt3_adt_net_165618_\);
    
    \I3.VDBi_57l6r_adt_net_3761_\ : AO21
      port map(A => REGl6r, B => 
        \I3.VDBi_57l7r_adt_net_142960__net_1\, C => 
        \I3.VDBi_57l6r_adt_net_143252__net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_3761__net_1\);
    
    \I2.DTO_9_IV_0_O2L2R_1205\ : NOR2
      port map(A => \I2.CRC32_1_SQMUXA_0_38\, B => 
        \I2.N_4193_377\, Y => \I2.DTO_9_ivl2r_adt_net_34812_\);
    
    \I2.PIPE1_DT_42_1_IVL21R_1388\ : OAI21FTF
      port map(A => REGl441r, B => 
        \I2.N_3234_adt_net_855648__net_1\, C => 
        \I2.PIPE1_DT_42l21r_adt_net_46867_\, Y => 
        \I2.PIPE1_DT_42l21r_adt_net_46873_\);
    
    \I2.DTESl11r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl11r, Q => 
        \I2.DTESl11r_net_1\);
    
    \I3.REGMAPl20r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un81_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl20r_net_1\);
    
    \I1.REG_74_0_iv_0l264r\ : AO21
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, C => 
        \I1.REG_74l264r_adt_net_124371_\, Y => \I1.REG_74l264r\);
    
    \I2.STATE3_ns_a7l13r\ : NOR2FT
      port map(A => \I2.STATE3l1r_net_1\, B => \I2.N_3015\, Y => 
        \I2.STATE3_nsl13r\);
    
    REGl375r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_276_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl375r\);
    
    \I5.REG_1l441r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_24_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl441r);
    
    \I1.REG_74_0_IV_0L371R_1830\ : AND2
      port map(A => \FBOUTl6r\, B => \I1.N_593\, Y => 
        \I1.REG_74l371r_adt_net_113396_\);
    
    \I2.CRC32_12_il20r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_111_i_i_0\, Y => 
        \I2.N_3937\);
    
    \I2.ROFFSETl1r_1244\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_917_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETL1R_506\);
    
    \I2.ROFFSETe_0_adt_net_27175_\ : NOR2
      port map(A => \I2.N_145\, B => \I2.N_3019\, Y => 
        \I2.ROFFSETe_0_adt_net_27175__net_1\);
    
    \I2.PIPE10_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_634_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl29r_net_1\);
    
    \I2.PIPE8_DT_16_0l13r\ : MUX2H
      port map(A => \I2.PIPE8_DTl13r_net_1\, B => 
        \I2.PIPE7_DTl13r_net_1\, S => 
        \I2.N_565_0_adt_net_855736__net_1\, Y => \I2.N_579\);
    
    \I1.BITCNT_315\ : MUX2L
      port map(A => \I1.BITCNTl2r_net_1\, B => \I1.N_415\, S => 
        \I1.N_68\, Y => \I1.BITCNT_315_net_1\);
    
    VDB_padl11r : IOB33PH
      port map(PAD => VDB(11), A => \I3.VDBml11r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl11r);
    
    \I1.PAGECNTl1r_adt_net_834904_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.PAGECNT_326_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNTl1r_adt_net_834904_Rd1__net_1\);
    
    \I2.G_EVNT_NUMl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_931_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl3r_net_1\);
    
    \I2.DT_TEMP_762\ : MUX2H
      port map(A => \I2.DT_TEMPl1r_net_1\, B => 
        \I2.DT_TEMP_7l1r_net_1\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.DT_TEMP_762_net_1\);
    
    REGl233r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_134_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl233r\);
    
    \I3.PIPEA1_12l24r\ : AND2
      port map(A => DPR_cl24r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854488__net_1\, Y => 
        \I3.PIPEA1_12l24r_net_1\);
    
    \I1.REG_18_sqmuxa_0_a2_0_0_a4\ : NAND2
      port map(A => \I1.N_238_RD1__314\, B => \I1.PAGECNTL9R_835\, 
        Y => \I1.N_267\);
    
    \I3.VDBOFFB_53_2474\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl1r_net_1\, Y => 
        \I3.VDBoffb_53_adt_net_162980_\);
    
    \I1.REG_74_0_IVL196R_2038\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.REG_4_sqmuxa\, 
        Y => \I1.REG_74l196r_adt_net_130925_\);
    
    \I2.LSRAM_WADDR_381\ : MUX2L
      port map(A => \I2.PIPE5_DTl21r_net_1\, B => 
        \I2.LSRAM_WADDRl0r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_WADDR_381_net_1\);
    
    \I2.LSRAM_RADDRil2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_RADDRi_501\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.LSRAM_RADDRil2r_net_1\);
    
    \I1.REG_1_161\ : MUX2H
      port map(A => \REGl260r\, B => \I1.REG_74l260r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_161_net_1\);
    
    \I3.VADm_0_a3l13r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl13r_net_1\, Y => \I3.VADml13r\);
    
    REGl360r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_261_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl360r\);
    
    \I2.BNC_IDl9r\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_52_0\, CLR => 
        \I2.N_4620_i_0\, SET => \I2.N_4608_i_0\, Q => 
        \I2.BNC_IDl9r_net_1\);
    
    \I3.REG_1_203\ : MUX2L
      port map(A => VDB_inl22r, B => \I3.REGl155r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\, Y => 
        \I3.REG_1_203_0\);
    
    \I2.OFFSET_37_26l0r\ : MUX2L
      port map(A => \REGl221r\, B => \I2.N_827\, S => 
        \I2.PIPE7_DTl26r_net_1\, Y => \I2.N_835\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I110_Y_1665\ : AOI21
      port map(A => \I2.I110_un1_Y_adt_net_71212_\, B => 
        \I2.N332\, C => \I2.ADD_18x18_fast_I110_Y_0\, Y => 
        \I2.N442_i_adt_net_71348_\);
    
    \I2.PIPE5_DT_6_0l1r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l1r\, B => 
        \I2.un27_pipe5_dt0l1r\, S => 
        \I2.dataout_0_adt_net_855800__net_1\, Y => \I2.N_1070\);
    
    \I2.FID_7_IVL4R_1724\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl52r, C => 
        \I2.STATE3l9r_net_1\, Y => \I2.FID_7l4r_adt_net_93158_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I92_Y\ : NOR2
      port map(A => \I2.N303_0_543\, B => \I2.N307_2\, Y => 
        \I2.N346_0\);
    
    \I2.UN1_ERR_WORDS_RDY_0_SQMUXA_0_0_A5_1032\ : AND3FTT
      port map(A => \I2.BITCNTl1r_net_1\, B => 
        \I2.BITCNTl5r_net_1\, C => \I2.STATE5l1r_net_1\, Y => 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23154_\);
    
    \I2.N_4669_adt_net_855052_\ : BFR
      port map(A => \I2.N_4669\, Y => 
        \I2.N_4669_adt_net_855052__net_1\);
    
    \I2.FID_7_0_IVL10R_971\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl10r_net_1\, 
        Y => \I2.FID_7l10r_adt_net_18363_\);
    
    \I1.REG_74_13_388_m8_i_a4_0\ : OR2
      port map(A => \I1.N_299_adt_net_833868_Rd1__net_1\, B => 
        \I1.REG_74_12_300_N_15_adt_net_3731__net_1\, Y => 
        \I1.REG_74_12_300_N_15\);
    
    \I1.PAGECNTL5R_2879\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_322_adt_net_854384__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL5R_311\);
    
    \I2.ADEl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl8r);
    
    \I1.PAGECNTlde_0_o2_2_1239\ : NAND2FT
      port map(A => \I1.N_310_RD1__335\, B => 
        \I1.N_311_i_i_Rd1__net_1\, Y => \I1.N_325_501\);
    
    \I1.REG_74_0_IV_0_0L259R_1966\ : AND2
      port map(A => \FBOUTl6r\, B => \I1.N_596\, Y => 
        \I1.REG_74l259r_adt_net_124884_\);
    
    \I3.REG_1_276\ : MUX2H
      port map(A => VDB_inl4r, B => \I3.REGl95r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_276_0\);
    
    \I3.REG_1_198\ : MUX2L
      port map(A => VDB_inl17r, B => \I3.REGl150r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\, Y => 
        \I3.REG_1_198_0\);
    
    \I2.PIPE7_DTL26R_2895\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl26r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL26R_349\);
    
    \I1.REG_74_0_IVL390R_1800\ : NOR2FT
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, Y => 
        \I1.REG_74l390r_adt_net_111042_\);
    
    \I2.STATE2_ns_o3_i_o2l1r\ : AND2FT
      port map(A => \I2.TEMPF_net_1\, B => 
        \I2.WR_SRAM_2_ADT_NET_748__39\, Y => \I2.N_4184\);
    
    \I2.LEAD_FLAG6_7_i_0l7r\ : AOI21
      port map(A => \I2.N_219\, B => \I2.N_484\, C => \I2.N_222\, 
        Y => \I2.N_4528_adt_net_63525_\);
    
    \I2.L2TYPEl13r_1553\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_602_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_I_0_IL13R_660\);
    
    \I3.REG3_129\ : MUX2L
      port map(A => VDB_inl4r, B => \I3.REG3l4r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855624__net_1\, Y => 
        \I3.REG3_129_net_1\);
    
    \I2.PIPE7_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl14r_net_1\);
    
    \I2.PIPE3_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl9r_net_1\);
    
    \I2.STATE2_NS_I_0L0R_1009\ : OAI21FTF
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, B => 
        \I2.N_4284\, C => \I2.N_2796_i_0_adt_net_21575_\, Y => 
        \I2.N_2796_i_0_adt_net_21536_\);
    
    \I2.DT_TEMP_7l26r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854236__net_1\, B => 
        \I2.DT_SRAMl26r_net_1\, Y => \I2.DT_TEMP_7l26r_net_1\);
    
    \I1.REG_74_0_IVL216R_2018\ : AND2
      port map(A => \FBOUTl3r\, B => \I1.REG_7_sqmuxa\, Y => 
        \I1.REG_74l216r_adt_net_129120_\);
    
    \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__2823\ : OR3
      port map(A => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_N_20_i\, B
         => \I2.DTE_cl_0_sqmuxa_2_adt_net_20059__net_1\, C => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20061__net_1\, Y => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__158\);
    
    \I2.SUB8l13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_516_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l13r_net_1\);
    
    \I2.PIPE7_DTl25r_1580\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL25R_687\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I164_Y_2655\ : OR3FFT
      port map(A => \I2.N309_0\, B => 
        \I2.N258_0_adt_net_854936__net_1\, C => 
        \I2.N495_i_adt_net_202144_\, Y => 
        \I2.N495_i_adt_net_207682_\);
    
    \I3.PIPEA_8l13r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854476__net_1\, B => 
        \I3.N_222\, Y => \I3.PIPEA_8l13r_net_1\);
    
    \I3.N_178_ADT_NET_1360__2806\ : OR2FT
      port map(A => \I3.N_2083\, B => 
        \I3.N_178_adt_net_134608__net_1\, Y => 
        \I3.N_178_ADT_NET_1360__126\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2513\ : AND2
      port map(A => \REGl219r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.N_2070_adt_net_163466_\);
    
    \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__2973\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__490\);
    
    \I2.un8_evread_1_adt_net_855780_\ : BFR
      port map(A => \I2.un8_evread_1\, Y => 
        \I2.un8_evread_1_adt_net_855780__net_1\);
    
    \I3.TCNT3l7r\ : DFFC
      port map(CLK => CLK_c, D => TCNT3_372, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT3l7r_net_1\);
    
    REGl256r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_157_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl256r\);
    
    \I2.PIPE1_DT_42_1_IVL18R_1400\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040__net_1\, 
        B => \I2.PIPE1_DT_12l18r_net_1\, Y => 
        \I2.PIPE1_DT_42l18r_adt_net_47441_\);
    
    \I2.PIPE6_DT_0_SQMUXA_I_O4_1595\ : AO21TTF
      port map(A => \I2.N_219\, B => \I2.N_4545\, C => 
        \I2.PIPE5_DTL30R_622\, Y => \I2.N_4551_adt_net_63757_\);
    
    \I2.STATE1_ns_a3l7r\ : NOR2FT
      port map(A => TDCDRYA_c, B => \I2.STATE1_ns_1l7r\, Y => 
        \I2.STATE1_nsl7r\);
    
    \I3.VASl8r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_70_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl8r_net_1\);
    
    \I2.NPRSFIF_328_1735\ : NOR3FTT
      port map(A => NMRSFIF_c_c, B => \I2.un1_STATE3_3\, C => 
        \I2.STATE3_i_il10r\, Y => \I2.NPRSFIF_328_adt_net_97261_\);
    
    \I2.DT_TEMP_779\ : MUX2H
      port map(A => \I2.DT_TEMPl18r_net_1\, B => 
        \I2.DT_TEMP_7l18r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__29\, Y => 
        \I2.DT_TEMP_779_net_1\);
    
    \I2.EVNT_WORDl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_724_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl11r_net_1\);
    
    \I3.VDBil15r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_355_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil15r_net_1\);
    
    \I1.REG_25_sqmuxa_0_a2_0_a2\ : AND2
      port map(A => \I1.N_590\, B => \I1.N_584\, Y => 
        \I1.REG_25_sqmuxa\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I214_Y\ : XOR2FT
      port map(A => \I2.N479\, B => \I2.SUB_21x21_fast_I214_Y_0\, 
        Y => \I2.SUB8_2l18r\);
    
    \I2.L2TYPE_4_0L15R_1615\ : NOR2
      port map(A => \I2.L2AS_adt_net_855724__net_1\, B => 
        \I2.N_4468\, Y => \I2.L2TYPE_4l15r_adt_net_66837_\);
    
    REGl273r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_174_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl273r\);
    
    \I2.un8_evread_1_adt_net_855784_\ : BFR
      port map(A => \I2.un8_evread_1\, Y => 
        \I2.un8_evread_1_adt_net_855784__net_1\);
    
    \I2.BNCID_VECTrff_7\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_7_258_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_7\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854196_\ : BFR
      port map(A => \I2.N_4667_1_ADT_NET_1046__35\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854196__net_1\);
    
    \I3.VDBI_31_I_A3_0_1L5R_2241\ : AO21
      port map(A => \I3.REGMAPL14R_735\, B => \I3.REGl96r\, C => 
        \I3.REGMAPl17r_adt_net_854292__net_1\, Y => 
        \I3.VDBi_31_i_a3_0_1l5r_adt_net_143654_\);
    
    \I2.PIPE1_DT_42_1_IVL11R_1459\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855752__net_1\, B => 
        \I2.PIPE1_DT_30l11r_net_1\, C => 
        \I2.PIPE1_DT_42l11r_adt_net_49689_\, Y => 
        \I2.PIPE1_DT_42l11r_adt_net_49705_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2699\ : OA21
      port map(A => \I2.PIPE4_DTL10R_476\, B => 
        \I2.PIPE4_DTL9R_472\, C => \I2.RAMDT4L12R_825\, Y => 
        \I2.N_152_i_0_adt_net_502546_\);
    
    \I1.REG_74l172r\ : OR3
      port map(A => \I1.N_41_8\, B => 
        \I1.N_113_adt_net_3714__net_1\, C => \I1.REG_2_sqmuxa\, Y
         => \I1.N_41\);
    
    \I3.N_1309_i\ : DFFCI
      port map(CLK => CLK_c, D => \I3.N_1193_ip\, CLR => 
        \HWRES_3_adt_net_738__net_1\, QBAR => \I3.N_1309_i_net_1\);
    
    \I2.ROFFSETl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_911_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl7r_net_1\);
    
    \I3.un171_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_558\, B => \I3.N_583\, Y => 
        \I3.un171_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_2672\ : NOR2
      port map(A => \I2.N_72_0\, B => \I2.N_95_0\, Y => 
        \I2.N525_0_adt_net_318530_\);
    
    \I2.resyn_0_I2_FID_443\ : MUX2H
      port map(A => FID_cl27r, B => \I2.FID_7l27r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855828__net_1\, 
        Y => \I2.FID_443\);
    
    \I2.DTESl23r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl23r, Q => 
        \I2.DTESl23r_net_1\);
    
    \I1.REG_74_0_ivl265r\ : AO21
      port map(A => \REGl265r\, B => 
        \I1.N_137_adt_net_854760__net_1\, C => 
        \I1.REG_74l265r_adt_net_124285_\, Y => \I1.REG_74l265r\);
    
    VDB_padl0r : IOB33PH
      port map(PAD => VDB(0), A => \I3.VDBml0r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl0r);
    
    \I3.N_1905_1_adt_net_855384_\ : BFR
      port map(A => \I3.N_1905_1\, Y => 
        \I3.N_1905_1_adt_net_855384__net_1\);
    
    \I3.PIPEA1l10r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_308_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l10r_net_1\);
    
    \I2.PIPE5_DT_6l18r\ : MUX2L
      port map(A => \I2.PIPE5_DT_6_dl18r_net_1\, B => 
        \I2.un27_pipe5_dt0l18r\, S => \I2.PIPE5_DT_6_sl19r_net_1\, 
        Y => \I2.PIPE5_DT_6l18r_net_1\);
    
    REGl229r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_130_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl229r\);
    
    \I2.OFFSET_37_21l7r\ : MUX2L
      port map(A => \I2.N_794\, B => \I2.N_770\, S => 
        \I2.PIPE7_DTL25R_683\, Y => \I2.N_802\);
    
    \I2.OFFSET_37_15l6r\ : MUX2L
      port map(A => \REGl235r\, B => \REGl171r\, S => 
        \I2.PIPE7_DTL27R_68\, Y => \I2.N_753\);
    
    \I2.PIPE3_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl23r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl23r_net_1\);
    
    \I2.PIPE10_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_614_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl9r_net_1\);
    
    \I1.REG_74_0_IV_0L365R_1836\ : AND2
      port map(A => \FBOUTl0r\, B => \I1.N_593\, Y => 
        \I1.REG_74l365r_adt_net_113912_\);
    
    \I2.PIPE8_DT_539\ : MUX2L
      port map(A => \I2.PIPE8_DTl11r_net_1\, B => 
        \I2.PIPE8_DT_21l11r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_539_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL23R_1376\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_339\, B => 
        \I2.EVNT_NUMl7r_net_1\, Y => 
        \I2.PIPE1_DT_42l23r_adt_net_46641_\);
    
    \I2.REG_1_C5_I_1742\ : AND2
      port map(A => REGl37r, B => 
        \I2.N_3834_i_0_adt_net_1384__net_1\, Y => 
        \I2.N_3834_i_0_adt_net_101432_\);
    
    \I2.CRC32l16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_811_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l16r_net_1\);
    
    \I2.MIC_REG3_321\ : MUX2L
      port map(A => \I2.MIC_REG3l5r_net_1\, B => 
        \I2.MIC_REG3l4r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\, Y => 
        \I2.MIC_REG3_321_net_1\);
    
    \I1.PAGECNT_n6_i_i_a4_0_826\ : OR2FT
      port map(A => \I1.UN1_SBYTE13_1_I_1_208\, B => 
        \I1.N_656_495\, Y => \I1.N_473_204\);
    
    \I2.TDCDBSl13r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl13r, Q => 
        \I2.TDCDBSl13r_net_1\);
    
    \I2.DTE_21_1_IV_0L6R_1323\ : AO21
      port map(A => \I2.DT_TEMPl6r_net_1\, B => \I2.N_4038\, C
         => \I2.DTE_21_1l6r_adt_net_38967_\, Y => 
        \I2.DTE_21_1l6r_adt_net_38981_\);
    
    \I4.bcnt_3l0r\ : AND2FT
      port map(A => \I4.bcntl0r_net_1\, B => \I4.N_48_3\, Y => 
        \I4.bcnt_3l0r_net_1\);
    
    \I3.VDBi_57l6r_adt_net_143252_\ : AO21FTT
      port map(A => \I2.N_4424\, B => \I3.N_2040\, C => 
        \I3.VDBi_57l6r_adt_net_143243__net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143252__net_1\);
    
    \I3.VDBi_29_0_a2_0l9r\ : NOR3FTT
      port map(A => \I3.REGMAPl2r_net_1\, B => 
        \I3.REGMAPl7r_net_1\, C => \I3.N_1907_262\, Y => 
        \I3.N_2040\);
    
    \I3.VAS_77\ : MUX2L
      port map(A => VAD_inl15r, B => \I3.VAS_i_0_il15r\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_77_net_1\);
    
    \I2.MIC_ERR_REGS_347\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl19r_net_1\, B => 
        \I2.MIC_ERR_REGSl18r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_347_net_1\);
    
    \I3.STATE1_TR24_I_0_A3_5_2113\ : AND3FFT
      port map(A => \I3.REGMAPl13r_net_1\, B => \I3.N_303\, C => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_1570__net_1\, Y => 
        \I3.STATE1_tr24_i_0_a3_5_i_adt_net_135637_\);
    
    \I2.DTO_16_1_IV_0_0L12R_1157\ : AND2FT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        B => \I2.DT_TEMPl12r_net_1\, Y => 
        \I2.DTO_16_1l12r_adt_net_32622_\);
    
    \I2.LSRAM_RADDRil0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_RADDRi_499\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.LSRAM_RADDRil0r_net_1\);
    
    \I3.VASl7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_69_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VAS_i_0_il7r\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_2673\ : AND2FT
      port map(A => 
        \I2.N_3_0_adt_net_1070__adt_net_855604__net_1\, B => 
        \I2.N525_0_adt_net_318487_\, Y => 
        \I2.N525_0_adt_net_58018_\);
    
    \I3.REG3l4r_1170\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_129_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3L4R_432\);
    
    \I3.TICKi_2l0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.un6_tcnt1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => TICKL0R_3);
    
    \I1.BYTECNT_n4_i\ : AND2FT
      port map(A => \I1.N_223\, B => \I1.N_1381_adt_net_109130_\, 
        Y => \I1.N_1381\);
    
    \I2.DT_TEMP_7l0r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, B => 
        \I2.DT_SRAMl0r_net_1\, Y => \I2.DT_TEMP_7l0r_net_1\);
    
    TDCDB_padl22r : IB33
      port map(PAD => TDCDB(22), Y => TDCDB_cl22r);
    
    \I2.STATE2_ns_i_0l0r\ : AND2FT
      port map(A => \I2.STATE2_ns_i_0_1_il0r\, B => 
        \I2.N_2796_i_0_adt_net_21536_\, Y => \I2.N_2796_i_0\);
    
    \I2.EVNT_NUM_n2_tz\ : XOR2FT
      port map(A => \I2.EVNT_NUMl2r_net_1\, B => 
        \I2.EVNT_NUM_c1_net_1\, Y => \I2.EVNT_NUM_n2_tz_i\);
    
    \I3.VDBI_57_0_IV_0_0L13R_2199\ : AO21
      port map(A => REGl61r, B => \I3.N_402_1\, C => 
        \I3.VDBi_57l13r_adt_net_140592_\, Y => 
        \I3.VDBi_57l13r_adt_net_140594_\);
    
    \I2.un21_pipe5_dt_2\ : XOR2
      port map(A => \I2.RAMDT4l4r_net_1\, B => 
        \I2.RAMDT4l3r_net_1\, Y => \I2.un21_pipe5_dt_2_net_1\);
    
    \I2.CRC32_12_i_x2l15r\ : XOR2FT
      port map(A => \I2.CRC32l15r_net_1\, B => \I2.N_3960_i_i\, Y
         => \I2.N_113_i_i_0\);
    
    \I2.PIPE5_DT_6_0l12r\ : MUX2L
      port map(A => \I2.un27_pipe5_dt1l12r\, B => 
        \I2.un27_pipe5_dt0l12r\, S => 
        \I2.dataout_0_adt_net_855804__net_1\, Y => \I2.N_1081\);
    
    \I3.STATE2_0_sqmuxa_0_a2_i\ : NAND2
      port map(A => \I3.DSS_425\, B => \I3.STATE2L0R_720\, Y => 
        \I3.N_1896\);
    
    \I1.REG_1_83\ : MUX2H
      port map(A => \REGl182r\, B => \I1.REG_74l182r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855396__net_1\, Y => 
        \I1.REG_1_83_net_1\);
    
    \I2.DTESl16r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl16r, Q => 
        \I2.DTESl16r_net_1\);
    
    \I3.PIPEA1_304\ : MUX2L
      port map(A => \I3.PIPEA1l6r_net_1\, B => 
        \I3.PIPEA1_12l6r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__254\, Y => 
        \I3.PIPEA1_304_net_1\);
    
    \I1.UN1_SBYTE13_2_I_I_A2_I_1776\ : AO21
      port map(A => \I1.N_341_Rd1__net_1\, B => \I1.N_332\, C => 
        \I1.N_223_adt_net_108706_\, Y => 
        \I1.N_223_adt_net_108707_\);
    
    \I3.un96_reg_ads_0_a2_0_a2\ : NAND3FFT
      port map(A => \I3.VASl4r_net_1\, B => \I3.N_549_364\, C => 
        \I3.VASl1r_net_1\, Y => \I3.N_585\);
    
    \I2.DTO_9_iv_0_o2_0l5r\ : MUX2H
      port map(A => \I2.DT_TEMP_7l5r_net_1\, B => 
        \I2.DT_TEMPl5r_net_1\, S => 
        \I2.TEMPF_adt_net_855740__adt_net_855896__net_1\, Y => 
        \I2.N_4266\);
    
    REGl321r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_222_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl321r\);
    
    \I2.PIPE1_DT_42_1_IV_2L27R_1364\ : NOR2
      port map(A => REGl431r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855816__net_1\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il27r_adt_net_46033_\);
    
    \I1.REG_74_0_ivl305r\ : AO21
      port map(A => \REGl305r\, B => \I1.N_177\, C => 
        \I1.REG_74l305r_adt_net_120438_\, Y => \I1.REG_74l305r\);
    
    \I2.PIPE5_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_685_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl9r_net_1\);
    
    \I3.REGMAPL25R_3022\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un106_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL25R_776\);
    
    \I2.L2SERVl1r_1504\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_921_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL13R_611\);
    
    \I2.RAMAD1_660\ : MUX2L
      port map(A => \I2.RAMAD1_12l6r_net_1\, B => 
        \I2.RAMAD1l6r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__172\, Y => 
        \I2.RAMAD1_660_net_1\);
    
    \I2.PIPE1_DT_757\ : MUX2L
      port map(A => \I2.PIPE1_DTl30r_net_1\, B => 
        \I2.PIPE1_DT_42l30r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854560__net_1\, 
        Y => \I2.PIPE1_DT_757_net_1\);
    
    \I2.PIPE1_DT_42_0_0l27r_963\ : NOR3
      port map(A => \I2.PIPE1_DT_42_0l27r_net_1\, B => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\, C => \I2.N_12169_i\, Y => 
        \I2.PIPE1_DT_42_3_0L28R_341\);
    
    \I2.PIPE1_DT_12l6r\ : MUX2L
      port map(A => \I2.TDCDASl6r_net_1\, B => 
        \I2.TDCDASl4r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855112__net_1\, Y
         => \I2.PIPE1_DT_12l6r_net_1\);
    
    \I2.N_4283_i_0_a2_m1_e_0\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854444__net_1\, 
        B => \I2.TEMPF_adt_net_855744__net_1\, Y => 
        \I2.N_4283_i_0\);
    
    \I2.SUB9_0_SQMUXA_0_A2_0_0_1001\ : NOR2
      port map(A => \I2.NWPIPE8_I_0_I_0_0_5\, B => 
        \I2.PIPE8_DTl30r_net_1\, Y => 
        \I2.SUB9_0_sqmuxa_0_adt_net_20771_\);
    
    \I2.SRAM_EVNT_c1_i\ : OAI21
      port map(A => \I2.N_3855\, B => \I2.N_128_1\, C => 
        \I2.N_135\, Y => \I2.N_3826\);
    
    \I3.VDBm_0l9r\ : MUX2L
      port map(A => \I3.PIPEAl9r_net_1\, B => \I3.PIPEBl9r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_151\);
    
    DPR_padl31r : IB33
      port map(PAD => DPR(31), Y => DPR_cl31r);
    
    REGl179r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_80_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl179r\);
    
    \I3.STATE2_nsl3r\ : AO21FTF
      port map(A => \I3.N_1465\, B => \I3.STATE2l1r_net_1\, C => 
        \I3.N_1463_i_1_adt_net_855356__net_1\, Y => 
        \I3.STATE2_nsl3r_net_1\);
    
    \I2.RAMADl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l0r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl0r);
    
    \I0.CLEARF1\ : DFFC
      port map(CLK => CLK_c, D => \I0.CLEAR_i_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I0.CLEARF1_net_1\);
    
    \I2.PIPE1_DT_42_1_ivl2r\ : OR2
      port map(A => \I2.PIPE1_DT_42l2r_adt_net_51838_\, B => 
        \I2.PIPE1_DT_42l2r_adt_net_51839_\, Y => 
        \I2.PIPE1_DT_42l2r\);
    
    \I1.REG_74_1_a0_0l228r_adt_net_854832_\ : BFR
      port map(A => \I1.REG_74_1_a0_0l228r\, Y => 
        \I1.REG_74_1_a0_0l228r_adt_net_854832__net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2433\ : AO21
      port map(A => \REGl336r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l3r_adt_net_162528_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162554_\);
    
    \I3.VDBI_57_0_IV_0_0L15R_2188\ : AO21
      port map(A => REGl63r, B => \I3.N_402_1\, C => 
        \I3.VDBi_57l15r_adt_net_139970_\, Y => 
        \I3.VDBi_57l15r_adt_net_139972_\);
    
    SYSRESB_pad : IB33
      port map(PAD => SYSRESB, Y => SYSRESB_c);
    
    \I3.VDBoffal3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_47_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal3r_net_1\);
    
    \I1.BYTECNT_I_0_IL1R_2918\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_313_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.BYTECNT_I_0_IL1R_435\);
    
    \I2.CRC32l20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_815_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l20r_net_1\);
    
    \I1.REG_74l188r_890\ : OR2
      port map(A => \I1.REG_4_sqmuxa\, B => 
        \I1.N_65_ADT_NET_1433__217\, Y => \I1.N_57_268\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I60_Y_1657\ : AND2
      port map(A => \I2.N294\, B => \I2.N297\, Y => 
        \I2.N328_adt_net_70573_\);
    
    \I2.OFFSET_37_6l3r\ : MUX2L
      port map(A => \I2.N_670\, B => \I2.N_662\, S => 
        \I2.PIPE7_DTL26R_353\, Y => \I2.N_678\);
    
    \I2.DTE_1l18r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l18r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l18r_Rd1__net_1\);
    
    \I3.VAS_71\ : MUX2L
      port map(A => VAD_inl9r, B => \I3.VASl9r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_71_net_1\);
    
    \I2.N_2828_adt_net_39955_\ : AO21FTF
      port map(A => \I2.N_176_i\, B => \I2.STATE2l5r_net_1\, C
         => \I2.N_4293\, Y => \I2.N_2828_adt_net_39955__net_1\);
    
    \I1.REG_1_301\ : MUX2H
      port map(A => \REGl400r\, B => \I1.REG_74l400r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855524__net_1\, Y => 
        \I1.REG_1_301_net_1\);
    
    \I2.BNCID_VECTrff_3\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_3_262_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_3\);
    
    \I3.VDBi_57_0_ivl25r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l25r_net_1\, C
         => \I3.VDBi_57l25r_adt_net_138713_\, Y => 
        \I3.VDBi_57l25r\);
    
    TDCDA_padl2r : IB33
      port map(PAD => TDCDA(2), Y => TDCDA_cl2r);
    
    \I3.TCNT1l0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT1_i_0l0r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT1l0r_net_1\);
    
    \I2.SUB8l7r_1598\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_510_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8L7R_705\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855424_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__22\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855424__net_1\);
    
    \I2.LSRAM_INl5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_389_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl5r_net_1\);
    
    \I2.SUB9_586\ : MUX2H
      port map(A => \I2.SUB9l18r_net_1\, B => \I2.SUB9_1l18r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_586_net_1\);
    
    \I3.PIPEA1l12r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_310_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l12r_net_1\);
    
    \I2.PIPE1_DT_42_1_IV_2L26R_1367\ : NOR2
      port map(A => \I2.TDCDASl26r_net_1\, B => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855036__net_1\, 
        Y => \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46167_\);
    
    \I2.OFFSETl6r_1566\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_566_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL6R_673\);
    
    \I3.REG_1_207\ : MUX2L
      port map(A => VDB_inl26r, B => \I3.REGl159r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\, Y => 
        \I3.REG_1_207_0\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I167_Y_1689\ : AND2
      port map(A => \I2.N319_0\, B => \I2.N315\, Y => 
        \I2.N504_adt_net_88887_\);
    
    \I2.STATEE_NSL3R_1024\ : AND2
      port map(A => \I2.CHAIN_ERRS_net_1\, B => \I2.STATEe_ipl1r\, 
        Y => \I2.STATEe_nsl3r_adt_net_22965_\);
    
    \I2.ROFFSET_n11\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855700__net_1\, B => 
        \I2.ROFFSET_n11_tz_i\, Y => \I2.ROFFSET_n11_net_1\);
    
    \I2.END_TDC1\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.END_TDC1_711_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.END_TDC1_net_1\);
    
    \I2.SUB9_588\ : MUX2H
      port map(A => \I2.SUB9l20r_net_1\, B => \I2.SUB9_1l20r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_588_net_1\);
    
    \I2.SRAM_EVNTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SRAM_EVNT_n4_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.SRAM_EVNTl4r_net_1\);
    
    \I2.DTO_16_1_IVL11R_1165\ : AND2FT
      port map(A => \I2.N_223\, B => \I2.DTE_2_1l11r_net_1\, Y
         => \I2.DTO_16_1l11r_adt_net_32872_\);
    
    \I1.REG_1_275\ : MUX2H
      port map(A => \REGl374r\, B => \I1.REG_74l374r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_275_net_1\);
    
    \I1.REG_74_0_IVL281R_1938\ : NOR2FT
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l281r_adt_net_122635_\);
    
    REGl320r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_221_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl320r\);
    
    \I2.PIPE8_DT_558_1671\ : AND2
      port map(A => \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, B => 
        \I2.PIPE8_DTl30r_net_1\, Y => 
        \I2.PIPE8_DT_558_adt_net_82590_\);
    
    \I2.FCNT_106\ : NOR2
      port map(A => \I2.FCNTl1r_net_1\, B => \I2.un1_STATE1_22\, 
        Y => \I2.N_1237\);
    
    \I2.RAMDT4L1R_3015\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl1r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L1R_769\);
    
    \I2.OFFSET_37_11l5r\ : MUX2L
      port map(A => \REGl378r\, B => \REGl314r\, S => 
        \I2.PIPE7_DTL27R_78\, Y => \I2.N_720\);
    
    \I2.DT_TEMP_772\ : MUX2H
      port map(A => \I2.DT_TEMPl11r_net_1\, B => 
        \I2.DT_TEMP_7l11r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__30\, Y => 
        \I2.DT_TEMP_772_net_1\);
    
    \I1.PAGECNTL6R_3080\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_321_adt_net_854880__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL6R_836\);
    
    \I2.DTO_16_1_iv_0_0l16r\ : OR2
      port map(A => \I2.DTO_16_1l16r_adt_net_31717_\, B => 
        \I2.DTO_16_1l16r_adt_net_31718_\, Y => \I2.DTO_16_1l16r\);
    
    \I2.PIPE7_DTl31r_1240\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl31r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL31R_502\);
    
    \I3.VDBi_4_il0r\ : AND2
      port map(A => REGl0r, B => \I3.REGMAPL1R_725\, Y => 
        \I3.N_2063_i\);
    
    \I2.PIPE10_DT_17_I_A3_2L13R_1611\ : OR3
      port map(A => \I2.N_3822_adt_net_64759_\, B => 
        \I2.SUB9_i_0_il9r\, C => \I2.SUB9l8r_net_1\, Y => 
        \I2.N_3822_adt_net_64764_\);
    
    \I2.DTO_16_1_iv_0l8r\ : OR2
      port map(A => \I2.DTO_16_1l8r_adt_net_33489_\, B => 
        \I2.DTO_16_1l8r_adt_net_33490_\, Y => \I2.DTO_16_1l8r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I73_Y\ : AND2
      port map(A => \I2.N243_0\, B => \I2.N240_0\, Y => 
        \I2.N323_0\);
    
    \I2.G_EVNT_NUM_n6_i_o2_1291\ : AND2FT
      port map(A => \I2.N_4669\, B => \I2.G_EVNT_NUMl5r_net_1\, Y
         => \I2.N_4672_553\);
    
    \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835180_Rd1_\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__net_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_775__adt_net_835180_Rd1__net_1\);
    
    REGl237r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_138_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl237r\);
    
    \I3.VDBOFFB_57_2402\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl5r_net_1\, Y => 
        \I3.VDBoffb_57_adt_net_162220_\);
    
    \I2.PIPE3_DTl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl25r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl25r_net_1\);
    
    \I1.REG_74_0_iv_0_0_o2l253r\ : OR2
      port map(A => \I1.N_661_adt_net_114476_\, B => 
        \I1.N_658_adt_net_124758_\, Y => \I1.N_658\);
    
    \I3.PIPEA_245\ : MUX2L
      port map(A => \I3.PIPEAl14r_net_1\, B => 
        \I3.PIPEA_8l14r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854668__net_1\, Y
         => \I3.PIPEA_245_net_1\);
    
    \I2.DTO_9_IV_0L23R_1098\ : AO21FTT
      port map(A => \I2.CRC32_1_sqmuxa_0\, B => 
        \I2.DT_SRAMl23r_net_1\, C => 
        \I2.DTO_9l23r_adt_net_30040_\, Y => 
        \I2.DTO_9l23r_adt_net_30048_\);
    
    \I1.REG_74_0_ivl277r\ : AO21
      port map(A => \REGl277r\, B => \I1.N_153\, C => 
        \I1.REG_74l277r_adt_net_122979_\, Y => \I1.REG_74l277r\);
    
    \I2.WROi_10_0_0\ : NAND2
      port map(A => \I2.WROi_10_1\, B => \I2.N_2836\, Y => 
        \I2.WROi_10\);
    
    \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_888_\ : AO21FTF
      port map(A => \I2.STATE2L2R_589\, B => 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_28083__net_1\, C
         => \I2.WOFFSETl0r_adt_net_854640__net_1\, Y => 
        \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_888__net_1\);
    
    \I2.SUB8_509\ : MUX2H
      port map(A => \I2.SUB8l6r_net_1\, B => \I2.SUB8_2l6r\, S
         => \I2.SUB8_1_sqmuxa_0_adt_net_855148__net_1\, Y => 
        \I2.SUB8_509_net_1\);
    
    \I1.REG_74_2_2L340R_1874\ : OR3FTT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__761\, B
         => \PULSE_0L0R_ADT_NET_834380_RD1__540\, C => 
        \I1.REG_74_2_2_il340r_adt_net_117061_\, Y => 
        \I1.REG_74_2_2_il340r_adt_net_117067_\);
    
    \I2.un1_DTO_cl_1_sqmuxa_2_0_o2_1_0\ : NOR2
      port map(A => NOESRAME_C_239, B => 
        \I2.WOFFSETl0r_adt_net_854644__net_1\, Y => \I2.N_4241_1\);
    
    \I2.PIPE8_DTl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_532_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl4r_net_1\);
    
    \I2.DTO_16_1_iv_0_0l19r\ : OR2
      port map(A => \I2.DTO_16_1l19r_adt_net_30979_\, B => 
        \I2.DTO_16_1l19r_adt_net_30980_\, Y => \I2.DTO_16_1l19r\);
    
    \I1.REG_74_0_iv_0_o2_0_a2l253r\ : AND3FFT
      port map(A => \I1.PAGECNT_0l9r_adt_net_835128_Rd1__net_1\, 
        B => \I1.PAGECNTl8r_net_1\, C => 
        \I1.PAGECNTl6r_adt_net_854924__net_1\, Y => \I1.N_4867_i\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_2679\ : OA21
      port map(A => \I2.N_107_adt_net_256840_\, B => 
        \I2.N525_adt_net_335996_\, C => \I2.N_2360_tz_tz\, Y => 
        \I2.N525_adt_net_57834_\);
    
    \I2.TRGSERVl2r_1475\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l2r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVL2R_582\);
    
    \I2.L2SERVl2r_1506\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_920_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL14R_613\);
    
    \I2.OFFSET_37_8l4r\ : MUX2L
      port map(A => \REGl361r\, B => \REGl297r\, S => 
        \I2.PIPE7_DTL27R_70\, Y => \I2.N_695\);
    
    \I2.TRGSERVl2r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l2r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVl2r_net_1\);
    
    \I2.OFFSET_37_16l6r\ : MUX2L
      port map(A => \REGl267r\, B => \REGl203r\, S => 
        \I2.PIPE7_DTL27R_77\, Y => \I2.N_761\);
    
    DTO_padl9r : IOB33PH
      port map(PAD => DTO(9), A => \I2.DTO_1l9r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl9r);
    
    \I2.FIDl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_425_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl9r);
    
    \I3.PIPEB_100_2323\ : NOR2FT
      port map(A => \I3.PIPEBl21r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_100_adt_net_159831_\);
    
    \I1.SBYTE_60\ : MUX2L
      port map(A => \FBOUTl2r\, B => \I1.N_190\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_60_net_1\);
    
    \I1.REG_74_0_IV_0L220R_2014\ : AND2
      port map(A => \REGl220r\, B => \I1.N_89_164\, Y => 
        \I1.REG_74l220r_adt_net_128776_\);
    
    \I1.BYTECNT_n1_i_0\ : NOR2
      port map(A => \I1.N_223_adt_net_854848__net_1\, B => 
        \I1.N_386_i_i_0\, Y => \I1.N_1161\);
    
    \I3.VDBOFFA_31_IV_0L1R_2601\ : AND2
      port map(A => \REGl238r\, B => \I3.REGMAPl27r_net_1\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164408_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I120_Y_0_76_TZ_TZ_1561\ : 
        AND2
      port map(A => \I2.RAMDT4L9R_768\, B => \I2.PIPE4_DTL2R_513\, 
        Y => \I2.N_2358_tz_tz_adt_net_55567_\);
    
    RAMDT_padl9r : IOB33PH
      port map(PAD => RAMDT(9), A => \I1.RAMDT_SPI_1l2r_net_1\, 
        EN => \I1.RAMDT_SPI_e_net_1\, Y => RAMDT_inl9r);
    
    \I2.PIPE1_DTl26r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_753_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl26r_net_1\);
    
    \I3.VDBil1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_341_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil1r_net_1\);
    
    \I3.REGMAPl3r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un17_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPl3r_net_1\);
    
    \I3.REG_1l74r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_175_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl74r);
    
    \I2.EVNT_NUM_957\ : MUX2L
      port map(A => \I2.EVNT_NUMl6r_net_1\, B => 
        \I2.EVNT_NUM_n6_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_957_net_1\);
    
    \I3.WRITES_23\ : MUX2L
      port map(A => WRITEB_c, B => \I3.WRITES_8\, S => 
        \I3.VSEL_0\, Y => \I3.WRITES_23_net_1\);
    
    \I2.BNCID_VECT_tile_DIN_REG1l0r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl0r_net_1\, Q => 
        \I2.DIN_REG1_0l0r\);
    
    \I2.DT_SRAM_0l19r\ : MUX2L
      port map(A => \I2.PIPE10_DTl19r_net_1\, B => 
        \I2.PIPE5_DTl19r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854220__net_1\, Y => 
        \I2.N_887\);
    
    \I2.CRC32_12_i_0_a2_1l6r\ : AND2
      port map(A => \I2.STATE2L0R_588\, B => 
        \I2.WR_SRAM_2_ADT_NET_748__39\, Y => \I2.N_2867_1\);
    
    \I2.TRGARR_3_I_11\ : XOR2
      port map(A => TDCTRG_c, B => \I2.TRGARRl0r_net_1\, Y => 
        \I2.DWACT_ADD_CI_0_partial_sum_2l0r\);
    
    \I2.OFFSET_37_19l3r\ : MUX2L
      port map(A => \REGl280r\, B => \REGl216r\, S => 
        \I2.PIPE7_DTL27R_90\, Y => \I2.N_782\);
    
    \I2.BITCNTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.BITCNT_937\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.BITCNTl3r_net_1\);
    
    \I2.PIPE1_DT_751\ : MUX2L
      port map(A => \I2.PIPE1_DTl24r_net_1\, B => 
        \I2.PIPE1_DT_42_1_iv_i_0l24r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854564__net_1\, 
        Y => \I2.PIPE1_DT_751_net_1\);
    
    \I2.WOFFSETl0r\ : DFFS
      port map(CLK => CLK_c, D => \I2.WOFFSET_827_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl0r_net_1\);
    
    \I2.LSRAM_WADDR_383\ : MUX2L
      port map(A => \I2.PIPE5_DTl23r_net_1\, B => 
        \I2.LSRAM_WADDRl2r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_WADDR_383_net_1\);
    
    \I4.un4_bcnt_I_12\ : AND2
      port map(A => \I4.bcnt_i_0_il2r_net_1\, B => \I4.N_7\, Y
         => \I4.N_4_0\);
    
    \I3.PIPEAl14r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_245_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl14r_net_1\);
    
    \I2.TEMPF_adt_net_855744_\ : BFR
      port map(A => \I2.TEMPF_net_1\, Y => 
        \I2.TEMPF_adt_net_855744__net_1\);
    
    \I2.OFFSET_37_25l6r\ : MUX2L
      port map(A => \REGl259r\, B => \REGl195r\, S => 
        \I2.PIPE7_DTL27R_88\, Y => \I2.N_833\);
    
    \I2.RAMAD_4l3r\ : MUX2L
      port map(A => \I2.N_530\, B => \I1.BYTECNTl3r_net_1\, S => 
        LOAD_RES, Y => \I2.RAMAD_4l3r_net_1\);
    
    \I3.N_178_adt_net_134608_\ : NAND2
      port map(A => \I3.N_2086\, B => \I3.N_177\, Y => 
        \I3.N_178_adt_net_134608__net_1\);
    
    \I3.PULSE_46_0_iv_i_il7r\ : AO21
      port map(A => PULSEl7r, B => 
        \I3.N_311_adt_net_854752__net_1\, C => \I3.N_318\, Y => 
        \I3.N_1897\);
    
    REGl176r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_77_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl176r\);
    
    FID_padl6r : OB33PH
      port map(PAD => FID(6), A => FID_cl6r);
    
    \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760_\ : BFR
      port map(A => \I2.PIPE1_DT_2_sqmuxa_1_1_net_1\, Y => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855760__net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I141_Y_0_O4_2682\ : 
        NAND2FT
      port map(A => \I2.N522_0_adt_net_329219_\, B => 
        \I2.N_96_0_adt_net_469923_\, Y => \I2.N522_0\);
    
    \I2.LEAD_FLAG6_641\ : AO21
      port map(A => \I2.N_4531_adt_net_1150__net_1\, B => 
        \I2.N_4531_adt_net_64140_\, C => 
        \I2.LEAD_FLAG6_641_adt_net_64180_\, Y => 
        \I2.LEAD_FLAG6_641_net_1\);
    
    SDAB_pad : IOB33PH
      port map(PAD => SDAB, A => \I5.SDAout_net_1\, EN => 
        un1_sdab_0_a2, Y => SDAB_in);
    
    \I1.PAGECNT_n6_i_i_o2_0\ : NAND2
      port map(A => \I1.PAGECNT_323_net_1\, B => \I1.N_308_Ra1_\, 
        Y => \I1.N_310_Ra1_\);
    
    \I3.un131_reg_ads_0_a2_1_a2\ : OR2
      port map(A => \I3.N_549\, B => \I3.N_586_adt_net_165970_\, 
        Y => \I3.N_586\);
    
    \I3.un47_reg_ads_0_a2_0_a2_991\ : OR2FT
      port map(A => \I3.WRITES_8\, B => \I3.N_546_373\, Y => 
        \I3.N_547_369\);
    
    \I3.REGMAPl2r_1630\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un13_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL2R_737\);
    
    \I3.REG3_226\ : OAI21FTF
      port map(A => \I3.REG3l405r_net_1\, B => \I3.N_1563\, C => 
        \I3.REG2_15l405r\, Y => \I3.REG3_226_net_1\);
    
    \I3.RAMAD_VME_31\ : MUX2H
      port map(A => RAMAD_VMEl7r, B => \I3.VASl8r_net_1\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_31_net_1\);
    
    \I3.un1_STATE2_7_1_adt_net_1473_\ : NAND2FT
      port map(A => \I3.STATE2l2r_net_1\, B => 
        \I3.NRDMEBi_0_sqmuxa_net_1\, Y => 
        \I3.un1_STATE2_7_1_adt_net_1473__net_1\);
    
    \I3.PIPEA1_303\ : MUX2L
      port map(A => \I3.PIPEA1l5r_net_1\, B => 
        \I3.PIPEA1_12l5r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__254\, Y => 
        \I3.PIPEA1_303_net_1\);
    
    \I3.RAMAD_VMEl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.RAMAD_VME_26_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => RAMAD_VMEl2r);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_499\ : MUX2H
      port map(A => \I2.PIPE4_DTl21r_net_1\, B => 
        \I2.LSRAM_RADDRil0r_net_1\, S => \I2.N_4642\, Y => 
        \I2.LSRAM_RADDRi_499\);
    
    \I3.REG_44_il85r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_1631_adt_net_150433_\, Y => \I3.N_1631\);
    
    \I2.resyn_0_I2_LSRAM_RADDRi_1_sqmuxa_0_a4_i_o2_46_tz\ : MUX2L
      port map(A => LEAD_FLAGl5r, B => LEAD_FLAGl4r, S => 
        \I2.PIPE4_DTl21r_net_1\, Y => \I2.N_2328_tz\);
    
    \I2.DTE_0_sqmuxa_i_o2_m6_i_1tt_m3_859\ : MUX2H
      port map(A => \I2.MIC_REG2L3R_ADT_NET_834020_RD1__491\, B
         => \I2.MIC_REG3L3R_484\, S => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_N_8_RD1__485\, Y => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_1TT_M3_237\);
    
    \I2.PIPE1_DT_30l8r\ : MUX2L
      port map(A => \I2.TDCDBSl8r_net_1\, B => 
        \I2.TDCDBSl6r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, Y
         => \I2.PIPE1_DT_30l8r_net_1\);
    
    \I2.CHAIN_ERRS\ : NOR2
      port map(A => \I2.CHAINA_ERRS_net_1\, B => 
        \I2.CHAINB_ERRS_net_1\, Y => \I2.CHAIN_ERRS_net_1\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2512\ : AND2
      port map(A => \REGl235r\, B => \I3.REGMAPl26r_net_1\, Y => 
        \I3.N_2070_adt_net_163462_\);
    
    \I2.PIPE1_DT_42_1_ivl11r\ : OR3
      port map(A => \I2.PIPE1_DT_42l11r_adt_net_49695_\, B => 
        \I2.PIPE1_DT_42l11r_adt_net_49704_\, C => 
        \I2.PIPE1_DT_42l11r_adt_net_49705_\, Y => 
        \I2.PIPE1_DT_42l11r\);
    
    \I2.N_4533_adt_net_1164_\ : AO21
      port map(A => \I2.PIPE5_DTl22r_net_1\, B => \I2.N_217\, C
         => LEAD_FLAGl2r, Y => \I2.N_4533_adt_net_1164__net_1\);
    
    REGl277r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_178_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl277r\);
    
    \I3.UN2_VSEL_1_I_0_2104\ : NOR3FFT
      port map(A => AMB_cl1r, B => AMB_cl0r, C => \I3.N_2055\, Y
         => \I3.N_1508_adt_net_135122_\);
    
    \I3.REG_1l65r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_166_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl65r);
    
    \I3.REGMAPL57R_2767\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un231_reg_ads_0_a2_4_a3_net_1\, Q => 
        \I3.REGMAPL57R_50\);
    
    \I1.REG_74_0_IVL265R_1958\ : AND2
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_13_sqmuxa_adt_net_855440__net_1\, Y => 
        \I1.REG_74l265r_adt_net_124285_\);
    
    \I3.VDBi_31l23r\ : MUX2L
      port map(A => \I3.REGl156r\, B => \I3.VDBi_20l23r\, S => 
        \I3.REGMAPl17r_adt_net_854284__net_1\, Y => 
        \I3.VDBi_31l23r_net_1\);
    
    \I1.REG_74_I_O2L364R_1841\ : AND3FTT
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536__net_1\, 
        B => \I1.REG_74_i_o2_0_0_364_m9_i_1_net_1\, C => 
        \I1.REG_74_i_o2_0_0_m9_i_0_0_net_1\, Y => 
        \I1.N_661_adt_net_114478_\);
    
    \I3.VDBI_57_0_IV_0_0L15R_2185\ : AO21
      port map(A => \I3.VDBil15r_net_1\, B => 
        \I3.N_1910_0_adt_net_854348__net_1\, C => 
        \I3.VDBi_57l15r_adt_net_139959_\, Y => 
        \I3.VDBi_57l15r_adt_net_139969_\);
    
    \I3.VDBOFFA_31_IV_0L0R_2627\ : AO21
      port map(A => \REGl221r\, B => \I3.REGMAPl25r_net_1\, C => 
        \I3.VDBoffa_31l0r_adt_net_164602_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164640_\);
    
    \I3.PIPEA_8l23r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854460__net_1\, B => 
        \I3.N_232\, Y => \I3.PIPEA_8l23r_net_1\);
    
    \I1.SBYTE_58\ : MUX2L
      port map(A => \FBOUTl0r\, B => \I1.N_186\, S => 
        \I1.SBYTE_0_sqmuxa\, Y => \I1.SBYTE_58_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL9R_1470\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855228__net_1\, B => 
        \I2.MIC_ERR_REGSl9r_net_1\, C => 
        \I2.PIPE1_DT_42l9r_adt_net_50197_\, Y => 
        \I2.PIPE1_DT_42l9r_adt_net_50198_\);
    
    \I2.PIPE1_DT_42_1_IVL4R_1499\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl36r_net_1\, C => 
        \I2.PIPE1_DT_42l4r_adt_net_51414_\, Y => 
        \I2.PIPE1_DT_42l4r_adt_net_51432_\);
    
    TOKOUTB_BP_pad : IB33
      port map(PAD => TOKOUTB_BP, Y => TOKOUTB_BP_c);
    
    \I5.sstate2se_3_i\ : MUX2L
      port map(A => \I5.sstate2l0r_net_1\, B => 
        \I5.sstate2l1r_net_1\, S => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\, Y => 
        \I5.sstate2se_3_i_net_1\);
    
    \I5.REG_1l424r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_37_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl424r);
    
    \I2.DTO_1_885\ : MUX2L
      port map(A => \I2.DTO_1l11r_Rd1__net_1\, B => 
        \I2.DTO_16_1l11r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834772_Rd1__net_1\, Y
         => \I2.DTO_1l11r\);
    
    \I3.TCNT2l1r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT2_395_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNT2l1r_net_1\);
    
    \I1.REG_1_70\ : MUX2H
      port map(A => \REGl169r\, B => \I1.REG_74l169r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855404__net_1\, Y => 
        \I1.REG_1_70_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I61_Y\ : NAND2
      port map(A => \I2.N261_0\, B => \I2.N258_0\, Y => 
        \I2.N311_0\);
    
    \I4.un1_lead_flag_1_2_0\ : MUX2L
      port map(A => LEAD_FLAGl6r, B => LEAD_FLAGl2r, S => 
        \I4.bcnt_i_0_il2r_net_1\, Y => \I4.N_2\);
    
    \I2.PIPE3_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl31r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl31r_net_1\);
    
    \I2.PIPE10_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_616_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl11r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I174_Y\ : XOR2
      port map(A => \I2.N394\, B => \I2.ADD_21x21_fast_I174_Y_0\, 
        Y => \I2.un27_pipe5_dt0l4r\);
    
    \I3.VDBml22r\ : MUX2L
      port map(A => \I3.VDBil22r_net_1\, B => \I3.N_164\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml22r_net_1\);
    
    \I2.PIPE5_DT_6l6r\ : MUX2L
      port map(A => \I2.PIPE4_DTl6r_net_1\, B => \I2.N_1075\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855620__net_1\, Y
         => \I2.PIPE5_DT_6l6r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I151_Y_i_a4_0\ : NAND3FFT
      port map(A => \I2.N_41_0_adt_net_55923_\, B => 
        \I2.N_41_0_adt_net_55921_\, C => \I2.N_163_0\, Y => 
        \I2.N_41_0\);
    
    \I2.WR_SRAM_2_adt_net_748__adt_net_854252_\ : BFR
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854260__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\);
    
    \I2.RAMADl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l13r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl13r);
    
    \I3.PIPEA_8_0l0r\ : MUX2L
      port map(A => DPR_cl0r, B => \I3.PIPEA1l0r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855364__net_1\, Y => \I3.N_209\);
    
    \I2.DTO_1_894\ : MUX2L
      port map(A => \I2.DTO_1l20r_Rd1__net_1\, B => 
        \I2.DTO_16_1l20r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834760_Rd1__net_1\, Y
         => \I2.DTO_1l20r\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I161_Y_1690\ : OA21FTF
      port map(A => \I2.N346_0\, B => \I2.N353\, C => \I2.N345\, 
        Y => \I2.N486_i_adt_net_89208_\);
    
    \I5.REG_1l426r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_39_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl426r);
    
    \I2.DTO_16_1_IV_0L8R_1179\ : AND2
      port map(A => \I2.N_182_ADT_NET_1007__386\, B => 
        \I2.DT_SRAMl8r_net_1\, Y => 
        \I2.DTO_16_1l8r_adt_net_33480_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I33_P0N_1762\ : OR2FT
      port map(A => \I2.LSRAM_OUTl12r\, B => 
        \I2.PIPE7_DTL12R_693\, Y => \I2.N267_0_869\);
    
    DTE_padl8r : IOB33PH
      port map(PAD => DTE(8), A => \I2.DTE_1l8r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl8r);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2715\ : AO21
      port map(A => \I2.N_45_1\, B => 
        \I2.N_152_i_0_adt_net_502543_\, C => 
        \I2.N_152_i_0_adt_net_610542_\, Y => 
        \I2.N_152_i_0_adt_net_610543_\);
    
    \I1.REG_74_9l356r\ : NAND3FTT
      port map(A => \I1.N_374\, B => \I1.N_1366\, C => 
        \I1.N_347_adt_net_854792__net_1\, Y => \I1.N_41_8\);
    
    \I2.PIPE9_DT_298\ : MUX2H
      port map(A => \I2.PIPE8_DTl29r_net_1\, B => 
        \I2.PIPE9_DTl29r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_298_net_1\);
    
    \I2.un3_tdcgda1_1_adt_net_821_\ : OR3FTT
      port map(A => \I2.TDCDASl30r_net_1\, B => 
        \I2.TDCDASl31r_net_1\, C => \I2.TDCDASl29r_net_1\, Y => 
        \I2.un3_tdcgda1_1_adt_net_821__net_1\);
    
    \I2.OFFSET_563\ : MUX2L
      port map(A => \I2.OFFSETl3r_net_1\, B => \I2.OFFSET_37l3r\, 
        S => \I2.UN1_NWPIPE7_2_298\, Y => \I2.OFFSET_563_net_1\);
    
    \I3.MYBERRi_62\ : MUX2H
      port map(A => MYBERR_c, B => \I3.DSS_9\, S => 
        \I3.un1_MYBERRi_1_sqmuxa\, Y => \I3.MYBERRi_62_net_1\);
    
    \I1.ISI_7_i_0_o4\ : OAI21FTF
      port map(A => \I1.sstatel6r_net_1\, B => 
        \I1.sstatel9r_net_1\, C => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854908__net_1\, Y
         => \I1.N_337\);
    
    \I3.UN6_TCNT1_2100\ : NOR3FTT
      port map(A => \I3.un6_tcnt1_adt_net_134941_\, B => 
        \I3.TCNT1l5r_net_1\, C => \I3.TCNT1_i_0_il3r_net_1\, Y
         => \I3.un6_tcnt1_adt_net_134944_\);
    
    \I2.RAMDT4L12R_3041\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_795\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I138_Y_0_0_1578\ : NOR3FFT
      port map(A => \I2.N_2360_tz_tz_adt_net_54584_\, B => 
        \I2.N_53\, C => \I2.N_80\, Y => 
        \I2.ADD_21x21_fast_I138_Y_0_0_adt_net_58475_\);
    
    \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__2830\ : OR3FFT
      port map(A => \I2.N_2870\, B => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\, C => 
        \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35789__net_1\, Y => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__174\);
    
    \I2.SUB9_1_ADD_18x18_fast_I26_Y\ : AND2FT
      port map(A => \I2.N_3558_i_net_1\, B => 
        \I2.N291_adt_net_4302__net_1\, Y => \I2.N291\);
    
    \I3.REG_1_169\ : MUX2L
      port map(A => VDB_inl20r, B => REGl68r, S => 
        \I3.N_1935_adt_net_855320__net_1\, Y => \I3.REG_1_169_0\);
    
    \I2.resyn_0_I2_BITCNT_n5_i\ : NOR2
      port map(A => \I2.ERR_WORDS_RDY_0_sqmuxa\, B => 
        \I2.N_28_i_0\, Y => \I2.N_4326\);
    
    \I2.PIPE4_DTl29r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl29r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl29r_net_1\);
    
    \I2.LEAD_FLAG6_7_i_0l1r\ : AOI21
      port map(A => \I2.N_4673\, B => \I2.N_483\, C => \I2.N_222\, 
        Y => \I2.N_4534_adt_net_64476_\);
    
    TDCDB_padl11r : IB33
      port map(PAD => TDCDB(11), Y => TDCDB_cl11r);
    
    \I2.SRAM_EVNT_c2_i_o2\ : AND2
      port map(A => \I2.N_3855\, B => \I2.SRAM_EVNTl2r_net_1\, Y
         => \I2.N_3858\);
    
    \I1.REG_74_0_ivl303r\ : AO21
      port map(A => \REGl303r\, B => \I1.N_177\, C => 
        \I1.REG_74l303r_adt_net_120610_\, Y => \I1.REG_74l303r\);
    
    \I3.VDBOFFA_31_IV_0L4R_2561\ : OR2
      port map(A => \I3.VDBoffa_31l4r_adt_net_163881_\, B => 
        \I3.VDBoffa_31l4r_adt_net_163882_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163887_\);
    
    \I2.un7_bnc_id_1_I_37\ : AND2
      port map(A => \I2.BNC_IDl6r_net_1\, B => \I2.N_29_0\, Y => 
        \I2.N_24_1\);
    
    \I2.L_LUT_498_1695\ : NOR3
      port map(A => \I2.NWPIPE4_576\, B => 
        \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\, C => 
        \I2.N_4595\, Y => \I2.L_LUT_498_adt_net_90208_\);
    
    \I2.PIPE1_DT_12l14r\ : MUX2L
      port map(A => \I2.TDCDASl14r_net_1\, B => 
        \I2.TDCDASl12r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, Y
         => \I2.PIPE1_DT_12l14r_net_1\);
    
    \I2.BITCNT_n2_i\ : NOR3
      port map(A => \I2.ERR_WORDS_RDY_0_sqmuxa\, B => \I2.N_4335\, 
        C => \I2.N_4328\, Y => \I2.N_4323\);
    
    VDB_padl4r : IOB33PH
      port map(PAD => VDB(4), A => \I3.VDBml4r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl4r);
    
    \I2.OFFSET_37_2l1r\ : MUX2L
      port map(A => \REGl382r\, B => \REGl318r\, S => 
        \I2.PIPE7_DTL27R_73\, Y => \I2.N_644\);
    
    \I2.STATE3_nsl6r\ : OAI21FTF
      port map(A => \I2.STATE3l5r_net_1\, B => 
        \I3.N_203_adt_net_854976__net_1\, C => 
        \I2.STATE3_nsl6r_adt_net_24857_\, Y => 
        \I2.STATE3_nsl6r_net_1\);
    
    \I3.VDBI_57_0_IV_0_0L24R_2157\ : AO21
      port map(A => REGl72r, B => \I3.N_1839\, C => 
        \I3.VDBi_57l24r_adt_net_138807_\, Y => 
        \I3.VDBi_57l24r_adt_net_138814_\);
    
    TDCDB_padl2r : IB33
      port map(PAD => TDCDB(2), Y => TDCDB_cl2r);
    
    \I2.L2TYPE_589\ : MUX2L
      port map(A => \I2.L2TYPEl0r_net_1\, B => \I2.N_4452\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_589_net_1\);
    
    \I2.PIPE9_DT_274\ : MUX2L
      port map(A => \I2.PIPE9_DTl5r_net_1\, B => 
        \I2.PIPE8_DTl5r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_274_net_1\);
    
    \I1.REG_74_0_IVL219R_2015\ : AND2
      port map(A => \FBOUTl6r\, B => \I1.REG_7_sqmuxa\, Y => 
        \I1.REG_74l219r_adt_net_128862_\);
    
    \I2.un15_clear_stat\ : OR2FT
      port map(A => CLEAR_STAT_12, B => \I2.CHAINB_ERRS_net_1\, Y
         => \I2.un15_clear_stat_i\);
    
    \I2.OFFSET_37_21l5r\ : MUX2L
      port map(A => \I2.N_792\, B => \I2.N_768\, S => 
        \I2.PIPE7_DTL25R_684\, Y => \I2.N_800\);
    
    \I1.REG_74_0_ivl227r\ : AO21
      port map(A => \REGl227r\, B => \I1.N_97\, C => 
        \I1.REG_74l227r_adt_net_128050_\, Y => \I1.REG_74l227r\);
    
    \I2.MIC_ERR_REGS_348\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl20r_net_1\, B => 
        \I2.MIC_ERR_REGSl19r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_348_net_1\);
    
    \I3.VDBil20r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_360_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil20r_net_1\);
    
    \I2.un7_bnc_id_1_I_56\ : XOR2
      port map(A => \I2.BNC_IDl10r_net_1\, B => \I2.N_11_1\, Y
         => \I2.I_56_0\);
    
    VDB_padl23r : IOB33PH
      port map(PAD => VDB(23), A => \I3.VDBml23r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl23r);
    
    \I2.EVNT_WORDl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_715_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl2r_net_1\);
    
    \I2.BNCID_VECTrff_7_258_0\ : AO21
      port map(A => \I2.BNCID_VECTwa15_1_net_1\, B => 
        \I2.BNCID_VECTrff_7_258_0_a2_0\, C => \I2.BNCID_VECTro_7\, 
        Y => \I2.BNCID_VECTrff_7_258_0_net_1\);
    
    \I5.SSTATE2SE_0_0_902\ : AOI21FTF
      port map(A => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\, B => 
        \I5.AIR_START_net_1\, C => \I5.sstate2l3r_net_1\, Y => 
        \I5.sstate2_ns_el1r_adt_net_8563_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I18_P0N_i_o2\ : NOR2
      port map(A => \I2.RAMDT4L12R_798\, B => 
        \I2.PIPE4_DTl18r_net_1\, Y => \I2.N_63_0\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608_\ : BFR
      port map(A => \I2.DTO_cl_1_sqmuxa_adt_net_1022__net_1\, Y
         => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608__net_1\);
    
    \I2.DTO_1_887\ : MUX2L
      port map(A => \I2.DTO_1l13r_Rd1__net_1\, B => 
        \I2.DTO_16_1l13r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834768_Rd1__net_1\, Y
         => \I2.DTO_1l13r\);
    
    \I2.LSRAM_INl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_392_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl8r_net_1\);
    
    \I2.FID_7_0_IVL22R_992\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl70r, C => 
        \I2.FID_7l22r_adt_net_19303_\, Y => 
        \I2.FID_7l22r_adt_net_19311_\);
    
    \I1.BITCNTlde_i_a2_0\ : OR2FT
      port map(A => \I1.N_457\, B => \I1.N_68_adt_net_108395_\, Y
         => \I1.N_68\);
    
    \I3.PIPEAl20r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_251_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl20r_net_1\);
    
    \I2.LSRAM_IN_394\ : MUX2L
      port map(A => \I2.PIPE5_DTl10r_net_1\, B => 
        \I2.LSRAM_INl10r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_394_net_1\);
    
    \I2.FID_418\ : MUX2H
      port map(A => FID_cl2r, B => \I2.FID_7l2r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855836__net_1\, 
        Y => \I2.FID_418_net_1\);
    
    \I1.sstate_ns_0_iv_0_il3r\ : AND2FT
      port map(A => 
        \PULSEl0r_adt_net_854532__adt_net_855544__net_1\, B => 
        \I1.N_420_i\, Y => \I1.sstate_ns_0_iv_0_il3r_net_1\);
    
    \I3.REG_1_212\ : MUX2L
      port map(A => VDB_inl31r, B => \I3.REGl164r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855292__net_1\, Y => 
        \I3.REG_1_212_0\);
    
    \I2.OFFSET_37_26l6r\ : MUX2L
      port map(A => \REGl227r\, B => \I2.N_833\, S => 
        \I2.PIPE7_DTL26R_360\, Y => \I2.N_841\);
    
    \I2.FCNT_945\ : MUX2L
      port map(A => \I2.FCNTl2r_net_1\, B => \I2.FCNT_n2_i\, S
         => \I2.N_3267\, Y => \I2.FCNT_945_net_1\);
    
    \I2.DTO_16_1_iv_0_a2_5l6r\ : AO21TTF
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855000__net_1\, 
        B => \I2.STATE2l4r_net_1\, C => \I2.N_223_156\, Y => 
        \I2.N_457\);
    
    \I2.DTE_21_1_IV_0L5R_1329\ : AO21
      port map(A => \I2.STATE2L3R_440\, B => \I2.DTO_9l5r\, C => 
        \I2.DTE_21_1l5r_adt_net_39100_\, Y => 
        \I2.DTE_21_1l5r_adt_net_39101_\);
    
    \I1.FBOUTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_65_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.FBOUTl7r_net_1\);
    
    \I1.REG_74_0_iv_i_a2_il206r\ : AO21
      port map(A => \REGl206r\, B => \I1.N_183_i_0\, C => 
        \I1.N_282_adt_net_130017_\, Y => \I1.N_282\);
    
    \I3.VDBOFFB_30_IV_0L7R_2350\ : AND2
      port map(A => \REGl380r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161752_\);
    
    \I2.sram_empty_1\ : XOR2
      port map(A => \I2.RPAGEL13R_611\, B => \I2.WPAGEL13R_751\, 
        Y => \I2.sram_empty_1_i_0_i\);
    
    \I2.DTO_1_879\ : MUX2L
      port map(A => \I2.DTO_1l5r_net_1\, B => \I2.DTO_16_1l5r\, S
         => \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => 
        \I2.DTO_1_879_net_1\);
    
    REGl165r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_66_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl165r\);
    
    \I2.DTE_1_859\ : MUX2L
      port map(A => \I2.DTE_1l21r_Rd1__net_1\, B => 
        \I2.DTE_21_1l21r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\, Y => 
        \I2.DTE_1l21r\);
    
    \I2.PIPE2_DTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl1r_net_1\);
    
    \I2.PIPE8_DT_547\ : MUX2L
      port map(A => \I2.PIPE8_DTl19r_net_1\, B => 
        \I2.PIPE8_DT_21l19r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_547_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2611\ : AO21
      port map(A => \REGl254r\, B => \I3.REGMAPl29r_net_1\, C => 
        \I3.VDBoffa_31l1r_adt_net_164420_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164452_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I22_Y\ : OA21TTF
      port map(A => \I2.N_3560_i_net_1\, B => 
        \I2.N_3558_i_adt_net_855584__net_1\, C => \I2.N_3562_i\, 
        Y => \I2.N287\);
    
    \I3.VDBOFFB_30_IV_0L6R_2383\ : OR3
      port map(A => \I3.VDBoffb_30l6r_adt_net_161987_\, B => 
        \I3.VDBoffb_30l6r_adt_net_161983_\, C => 
        \I3.VDBoffb_30l6r_adt_net_161984_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161990_\);
    
    \I2.PIPE1_DT_42_0_0l27r\ : NOR3
      port map(A => \I2.PIPE1_DT_42_0l27r_net_1\, B => 
        \I2.un1_PIPE1_DT_1_sqmuxa_2\, C => \I2.N_12169_i\, Y => 
        \I2.PIPE1_DT_42_3_0l28r\);
    
    \I2.END_TDC4\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_TDC3_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_TDC4_net_1\);
    
    \I2.TDCDASl3r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl3r, Q => 
        \I2.TDCDASl3r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2594\ : AO21
      port map(A => \REGl167r\, B => \I3.REGMAPl18r_net_1\, C => 
        \I3.VDBoffa_31l2r_adt_net_164234_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164263_\);
    
    \I5.sstate1l13r\ : DFFS
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el0r\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SSTATE1L13R_4\);
    
    \I3.VDBi_43l11r\ : MUX2L
      port map(A => REGl417r, B => \I3.VDBi_40l11r_net_1\, S => 
        \I3.REGMAPl55r_net_1\, Y => \I3.VDBi_43l11r_net_1\);
    
    \I2.MIC_ERR_REGSl35r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_364_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl35r_net_1\);
    
    \I3.REG_1l150r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_198_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl150r\);
    
    \I3.VDBoffl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoff_119_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffl3r_net_1\);
    
    \I2.un78_pipe5_dt_4\ : XOR2
      port map(A => \I2.un78_pipe5_dt_3_net_1\, B => 
        \I2.un78_pipe5_dt_2_net_1\, Y => 
        \I2.un78_pipe5_dt_4_net_1\);
    
    \I2.DTE_21_1l27r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l27r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l27r_Rd1__net_1\);
    
    \I3.VDBi_57_0_iv_0_a2_3l13r_742\ : OR2
      port map(A => \I3.REGMAPl17r_net_1\, B => \I3.N_2014_122\, 
        Y => \I3.N_2015_120\);
    
    \I2.OFFSET_37_29l3r\ : MUX2L
      port map(A => \I2.N_854\, B => \I2.N_742\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l3r\);
    
    \I2.EVNT_NUM_952\ : MUX2L
      port map(A => \I2.EVNT_NUMl11r_net_1\, B => 
        \I2.EVNT_NUM_n11_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_952_net_1\);
    
    \I2.OFFSET_37_4l1r\ : MUX2L
      port map(A => \REGl366r\, B => \REGl302r\, S => 
        \I2.PIPE7_DTL27R_73\, Y => \I2.N_660\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I154_Y_0\ : AOI21
      port map(A => \I2.N_65\, B => \I2.N_82\, C => \I2.N307\, Y
         => \I2.N502_i\);
    
    \I3.RAMDTSl4r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl4r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl4r_net_1\);
    
    \I2.DTO_cl_0_sqmuxa_0_adt_net_855192_\ : BFR
      port map(A => \I2.DTO_cl_0_sqmuxa_0\, Y => 
        \I2.DTO_cl_0_sqmuxa_0_adt_net_855192__net_1\);
    
    \I3.PIPEA_8l1r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854464__net_1\, B => 
        \I3.N_210\, Y => \I3.PIPEA_8l1r_net_1\);
    
    \I2.PIPE9_DT_297\ : MUX2L
      port map(A => \I2.PIPE9_DTl28r_net_1\, B => 
        \I2.PIPE8_DTl28r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_297_net_1\);
    
    \I2.PIPE1_DT_12l12r\ : MUX2L
      port map(A => \I2.TDCDASl12r_net_1\, B => 
        \I2.TDCDASl10r_net_1\, S => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855108__net_1\, Y
         => \I2.PIPE1_DT_12l12r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2436\ : OR3
      port map(A => \I3.VDBoffb_30l3r_adt_net_162555_\, B => 
        \I3.VDBoffb_30l3r_adt_net_162549_\, C => 
        \I3.VDBoffb_30l3r_adt_net_162550_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162559_\);
    
    \I2.PIPE1_DT_42_1_IVL15R_1434\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855224__net_1\, B => 
        \I2.MIC_ERR_REGSl15r_net_1\, C => 
        \I2.PIPE1_DT_42l15r_adt_net_48715_\, Y => 
        \I2.PIPE1_DT_42l15r_adt_net_48716_\);
    
    \I3.VDBOFFA_31_IV_0L4R_2554\ : AO21
      port map(A => \REGl193r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.VDBoffa_31l4r_adt_net_163838_\, Y => 
        \I3.VDBoffa_31l4r_adt_net_163879_\);
    
    VDB_padl10r : IOB33PH
      port map(PAD => VDB(10), A => \I3.VDBml10r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl10r);
    
    \I3.REGMAP_i_0_il58r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un235_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il58r_net_1\);
    
    \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__2909\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_320_adt_net_854876__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__363\);
    
    \I2.FID_7_IVL4R_1725\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl4r_net_1\, 
        C => \I2.FID_7l4r_adt_net_93151_\, Y => 
        \I2.FID_7l4r_adt_net_93159_\);
    
    \I2.DTE_21_1_IVL15R_1276\ : OR3
      port map(A => \I2.DTO_16_1l15r_adt_net_31956_\, B => 
        \I2.DTE_21_1l15r_adt_net_37943_\, C => 
        \I2.DTE_21_1l15r_adt_net_37950_\, Y => 
        \I2.DTE_21_1l15r_adt_net_37952_\);
    
    \I2.STATE1l12r_1539\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl6r_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STATE1L12R_646\);
    
    \I2.TOKOUTBS\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKOUTBS_3_i_net_1\, 
        Q => \I2.TOKOUTBS_net_1\);
    
    \I2.DTE_21_1_IV_2L0R_1346\ : OAI21TTF
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_290\, B => 
        \I2.DT_SRAMl0r_net_1\, C => 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39732_\, Y => 
        \I2.DTE_21_1_iv_2_il0r_adt_net_39733_\);
    
    \I3.UN1_MYBERRI_1_SQMUXA_0_0_2346\ : AND3FTT
      port map(A => \I3.DSS_net_1\, B => \I3.STATE1_ipl5r\, C => 
        \I3.un1_MYBERRi_1_sqmuxa_adt_net_161483_\, Y => 
        \I3.un1_MYBERRi_1_sqmuxa_adt_net_161480_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I58_Y_1679\ : AND2FT
      port map(A => \I2.LSRAM_OUTl11r\, B => 
        \I2.PIPE7_DTl11r_net_1\, Y => \I2.N308_0_adt_net_86492_\);
    
    \I2.PIPE1_DT_752\ : MUX2L
      port map(A => \I2.PIPE1_DTl25r_net_1\, B => 
        \I2.PIPE1_DT_42_1_iv_i_0l25r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854564__net_1\, 
        Y => \I2.PIPE1_DT_752_net_1\);
    
    AMB_padl0r : IB33
      port map(PAD => AMB(0), Y => AMB_cl0r);
    
    \I3.PULSEl3r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_333_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEl3r);
    
    \I2.PIPE8_DT_21l2r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl2r\, B => \I2.N_568\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l2r_net_1\);
    
    \I3.TCNT2_n2\ : XOR2
      port map(A => \I3.TCNT2_i_0_il2r_net_1\, B => \I3.TCNT2_c1\, 
        Y => \I3.TCNT2_n2_net_1\);
    
    \I3.un1_STATE1_13_1_adt_net_1351_\ : OR3
      port map(A => \I3.un1_STATE1_13_1_adt_net_137890__net_1\, B
         => \I3.un1_STATE1_13_1_adt_net_137896__net_1\, C => 
        \I3.un1_STATE1_13_1_adt_net_137902__net_1\, Y => 
        \I3.un1_STATE1_13_1_adt_net_1351__net_1\);
    
    \I2.LSRAM_IN_396\ : MUX2L
      port map(A => \I2.PIPE5_DTl12r_net_1\, B => 
        \I2.LSRAM_INl12r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_396_net_1\);
    
    \I2.DT_TEMP_7l4r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, B => 
        \I2.DT_SRAMl4r_net_1\, Y => \I2.DT_TEMP_7l4r_net_1\);
    
    \I5.TEMPDATA_79\ : MUX2L
      port map(A => \I5.TEMPDATAl5r_net_1\, B => REGl130r, S => 
        \I5.N_443\, Y => \I5.TEMPDATA_79_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I165_Y\ : AO21TTF
      port map(A => \I2.N510\, B => \I2.N498_1_adt_net_88035_\, C
         => \I2.N353\, Y => \I2.N498_1\);
    
    \I2.PIPE1_DT_42_1_IVL10R_1464\ : AO21FTT
      port map(A => \I2.N_3279_0_adt_net_855228__net_1\, B => 
        \I2.MIC_ERR_REGSl10r_net_1\, C => 
        \I2.PIPE1_DT_42l10r_adt_net_49950_\, Y => 
        \I2.PIPE1_DT_42l10r_adt_net_49951_\);
    
    \I0.EV_RESF2_i_0\ : NAND2FT
      port map(A => \HWRES_3_ADT_NET_738__17\, B => CLEAR_STAT_12, 
        Y => \I0.un4_hwresi_i\);
    
    \I2.un2_evnt_word_I_19\ : AND2
      port map(A => \I2.WOFFSETl3r_adt_net_854988__net_1\, B => 
        \I2.DWACT_FINC_E_0l0r\, Y => \I2.N_42\);
    
    \I2.PIPE1_DT_42_1_IVL3R_1502\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl19r_net_1\, Y => 
        \I2.PIPE1_DT_42l3r_adt_net_51617_\);
    
    \I1.BYTECNT_i_0_il1r\ : DFFC
      port map(CLK => CLK_c, D => \I1.BYTECNT_313_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.BYTECNT_i_0_il1r_net_1\);
    
    \I2.DTO_16_1_iv_0_1l2r\ : AO21FTT
      port map(A => \I2.DTO_1l2r_net_1\, B => \I2.N_196_53\, C
         => \I2.DTO_16_1_iv_0_1l2r_adt_net_34868_\, Y => 
        \I2.DTO_16_1_iv_0_1l2r_net_1\);
    
    \I1.REG_1_201\ : MUX2H
      port map(A => \REGl300r\, B => \I1.REG_74l300r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\, Y
         => \I1.REG_1_201_net_1\);
    
    \I2.EVNT_NUMl3r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.EVNT_NUM_960_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.EVNT_NUMl3r_net_1\);
    
    \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834760_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_0_sqmuxa_i_0_N_3_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834760_Rd1__net_1\);
    
    \I2.resyn_0_I2_FID_440\ : MUX2H
      port map(A => FID_cl24r, B => \I2.FID_7l24r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855832__net_1\, 
        Y => \I2.FID_440\);
    
    \I3.un37_reg_ads_0_a2_1_a2_1\ : NAND2
      port map(A => \I3.VASl4r_net_1\, B => \I3.VASl1r_net_1\, Y
         => \I3.N_555\);
    
    \I3.REG1l6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG1_139_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l6r_net_1\);
    
    \I2.DTOSl24r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl24r, Q => 
        \I2.DTOSl24r_net_1\);
    
    \I3.VDBoffal7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBoffa_51_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBoffal7r_net_1\);
    
    \I2.RAMDT4L9R_3014\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl9r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L9R_768\);
    
    \I3.REGMAPL43R_2928\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un196_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAPL43R_445\);
    
    \I3.PIPEA1l15r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_313_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l15r_net_1\);
    
    \I2.DTO_1l26r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l26r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l26r_Rd1__net_1\);
    
    \I1.REG_74_12_284_m10_i_0\ : OR2
      port map(A => \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_1_Ra1_\, B
         => \I3.PULSE_330_net_1\, Y => 
        \I1.REG_74_1_380_m8_i_0_Ra1_\);
    
    \I2.FIRST_TDC_1_sqmuxa_1_0_923\ : OR2FT
      port map(A => \I2.STATE1l12r_net_1\, B => 
        \I2.END_CHAINA1_1_sqmuxa_3\, Y => 
        \I2.NWPIPE1_4_SQMUXA_1_0_301\);
    
    \I2.FID_7_0_IVL16R_959\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl16r_net_1\, 
        Y => \I2.FID_7l16r_adt_net_17799_\);
    
    \I1.BYTECNT_N6_I_0_1781\ : XOR2FT
      port map(A => \I1.BYTECNTl6r_net_1\, B => \I1.N_335\, Y => 
        \I1.N_77_adt_net_109270_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I32_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl11r\, B => 
        \I2.PIPE7_DTL11R_694\, Y => \I2.N264_0\);
    
    \I3.VDBOFFB_30_IV_0L0R_2486\ : AO21
      port map(A => \REGl309r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        C => \I3.VDBoffb_30l0r_adt_net_163094_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163123_\);
    
    \I2.STATE2_NS_4_0L2R_1048\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.N_4282\, Y => \I2.STATE2_nsl2r_adt_net_24907_\);
    
    \I2.DTO_1l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1_876_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l2r_net_1\);
    
    \I2.PIPE1_DTl28r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_755_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl28r_net_1\);
    
    \I2.DTE_1_865\ : MUX2L
      port map(A => \I2.DTE_1l27r_Rd1__net_1\, B => 
        \I2.DTE_21_1l27r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\, Y => 
        \I2.DTE_1l27r\);
    
    ADO_padl2r : OB33PH
      port map(PAD => ADO(2), A => ADO_cl2r);
    
    \I1.REG_74_1_396_m7_i_3_adt_net_854840_\ : BFR
      port map(A => \I1.REG_74_1_396_m7_i_3\, Y => 
        \I1.REG_74_1_396_m7_i_3_adt_net_854840__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I175_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_801\, B => 
        \I2.PIPE4_DTl5r_adt_net_854412__adt_net_855600__net_1\, Y
         => \I2.ADD_21x21_fast_I175_Y_0_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I138_Y_0_a2_2\ : AO21
      port map(A => \I2.PIPE4_DTL11R_842\, B => 
        \I2.PIPE4_DTL12R_856\, C => \I2.RAMDT4L5R_812\, Y => 
        \I2.N_114_adt_net_275711_\);
    
    \I2.BNCID_VECT_tile_0_I_1\ : RAM256x9SA
      port map(DO8 => OPEN, DO7 => OPEN, DO6 => OPEN, DO5 => OPEN, 
        DO4 => OPEN, DO3 => \I2.DOUT_TMPl3r\, DO2 => 
        \I2.DOUT_TMPl2r\, DO1 => \I2.DOUT_TMPl1r\, DO0 => 
        \I2.DOUT_TMPl0r\, WPE => OPEN, RPE => OPEN, DOS => OPEN, 
        WADDR7 => \GND\, WADDR6 => \GND\, WADDR5 => \GND\, WADDR4
         => \GND\, WADDR3 => \I2.TRGARRl3r_net_1\, WADDR2 => 
        \I2.TRGARRl2r_net_1\, WADDR1 => \I2.TRGARRl1r_net_1\, 
        WADDR0 => \I2.TRGARRl0r_net_1\, RADDR7 => \GND\, RADDR6
         => \GND\, RADDR5 => \GND\, RADDR4 => \GND\, RADDR3 => 
        \I2.TRGSERVl3r_net_1\, RADDR2 => \I2.TRGSERVL2R_584\, 
        RADDR1 => \I2.TRGSERVl1r_net_1\, RADDR0 => 
        \I2.TRGSERVl0r_net_1\, DI8 => \GND\, DI7 => \GND\, DI6
         => \GND\, DI5 => \GND\, DI4 => \GND\, DI3 => 
        \I2.BNC_IDl11r_net_1\, DI2 => \I2.BNC_IDl10r_net_1\, DI1
         => \I2.BNC_IDl9r_net_1\, DI0 => \I2.BNC_IDl8r_net_1\, 
        WRB => \I2.TDCTRG_c_i_0\, RDB => \GND\, WBLKB => \GND\, 
        RBLKB => \GND\, PARODD => \VCC\, WCLKS => CLK_c, DIS => 
        \VCC\);
    
    \I1.REG_74_0_iv_0_0l253r\ : AO21
      port map(A => \REGl253r\, B => \I1.N_658\, C => 
        \I1.REG_74l253r_adt_net_125400_\, Y => \I1.REG_74l253r\);
    
    \I2.PIPE3_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl28r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl28r_net_1\);
    
    \I2.N_2826_1_adt_net_40738_\ : OA21FTT
      port map(A => \I2.N_176_I_157\, B => 
        \I2.WR_SRAM_2_ADT_NET_748__39\, C => \I2.STATE2l5r_net_1\, 
        Y => \I2.N_2826_1_adt_net_40738__net_1\);
    
    \I2.PIPE1_DT_42_1_IVL15R_1430\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044__net_1\, 
        B => \I2.PIPE1_DT_12l15r_net_1\, Y => 
        \I2.PIPE1_DT_42l15r_adt_net_48701_\);
    
    \I3.PIPEA_249\ : MUX2L
      port map(A => \I3.PIPEAl18r_net_1\, B => 
        \I3.PIPEA_8l18r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854664__net_1\, Y
         => \I3.PIPEA_249_net_1\);
    
    \I2.N_176_i_adt_net_855708_\ : BFR
      port map(A => \I2.N_176_i\, Y => 
        \I2.N_176_i_adt_net_855708__net_1\);
    
    \I2.OFFSETl6r_1565\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_566_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL6R_672\);
    
    \I2.OFFSET_37_19l4r\ : MUX2L
      port map(A => \REGl281r\, B => \REGl217r\, S => 
        \I2.PIPE7_DTL27R_89\, Y => \I2.N_783\);
    
    \I3.VDBi_40_1l4r\ : AND2FT
      port map(A => \I3.REGMAPl16r_net_1\, B => 
        \I3.VDBi_31l4r_net_1\, Y => \I3.N_342\);
    
    N_1_I3_TCNT2_390 : MUX2H
      port map(A => \I3.TCNT2_i_0_il6r_net_1\, B => 
        \N_1.I3.TCNT2_n6\, S => TICKL0R_558, Y => TCNT2_390);
    
    \I2.OFFSET_37_15l0r\ : MUX2L
      port map(A => \REGl229r\, B => \REGl165r\, S => 
        \I2.PIPE7_DTL27R_68\, Y => \I2.N_747\);
    
    \I2.RAMAD1_12l16r\ : MUX2L
      port map(A => \I2.TDCDASl27r_net_1\, B => 
        \I2.TDCDBSl27r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855184__net_1\, Y => 
        \I2.RAMAD1_12l16r_net_1\);
    
    \I1.REG_1_75\ : MUX2H
      port map(A => \REGl174r\, B => \I1.REG_74l174r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855400__net_1\, Y => 
        \I1.REG_1_75_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I152_Y_0\ : AND3FFT
      port map(A => \I2.N313\, B => \I2.N_103\, C => 
        \I2.N498_adt_net_56484_\, Y => \I2.N498\);
    
    \I2.DTE_21_1_IVL15R_1274\ : AND2FT
      port map(A => \I2.DTE_CL_0_SQMUXA_2_0_288\, B => 
        \I2.DT_SRAMl15r_net_1\, Y => 
        \I2.DTE_21_1l15r_adt_net_37943_\);
    
    \I2.L2TYPE_4_IL13R_1618\ : OR2
      port map(A => \I2.N_4455\, B => \I2.N_4457\, Y => 
        \I2.N_4439_adt_net_67071_\);
    
    \I1.REG_74_0_ivl330r\ : AO21
      port map(A => \REGl330r\, B => \I1.N_201\, C => 
        \I1.REG_74l330r_adt_net_118088_\, Y => \I1.REG_74l330r\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2516\ : AND2
      port map(A => \REGl283r\, B => \I3.REGMAP_i_0_il32r_net_1\, 
        Y => \I3.N_2070_adt_net_163478_\);
    
    VDB_padl29r : IOB33PH
      port map(PAD => VDB(29), A => \I3.VDBml29r_net_1\, EN => 
        NOE32R_c_i_0, Y => VDB_inl29r);
    
    \I3.REG_1_i_il18r\ : AO21
      port map(A => \I3.REG3l405r_net_1\, B => 
        \I3.REG2l405r_net_1\, C => \REGl18r_adt_net_15773_\, Y
         => REGl18r);
    
    \I3.REG_1l147r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_195_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl147r\);
    
    \I2.N_4283_i_0_adt_net_854968_\ : BFR
      port map(A => \I2.N_4283_I_0_235\, Y => 
        \I2.N_4283_i_0_adt_net_854968__net_1\);
    
    \I2.DTO_16_1_IV_0_0L25R_1089\ : AO21
      port map(A => \I2.N_197_150\, B => \I2.DT_SRAMl25r_net_1\, 
        C => \I2.DTO_16_1l25r_adt_net_29614_\, Y => 
        \I2.DTO_16_1l25r_adt_net_29624_\);
    
    \I2.DTE_21_1_IV_0_0L22R_1253\ : AO21FTT
      port map(A => \I2.DTE_cl_0_sqmuxa_2_0\, B => 
        \I2.DT_SRAMl22r_net_1\, C => 
        \I2.DTE_21_1l22r_adt_net_37393_\, Y => 
        \I2.DTE_21_1l22r_adt_net_37394_\);
    
    \I1.REG_1_101\ : MUX2H
      port map(A => \REGl200r\, B => \I1.N_1339\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\, Y => 
        \I1.REG_1_101_net_1\);
    
    \I2.TRGCNTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TRGCNT_n3\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGCNT_i_0_il3r\);
    
    \I1.REG_74_0_IVL334R_1882\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l334r_adt_net_117744_\);
    
    \I3.REGMAPl23r_adt_net_855012_\ : BFR
      port map(A => \I3.REGMAPl23r_adt_net_855016__net_1\, Y => 
        \I3.REGMAPl23r_adt_net_855012__net_1\);
    
    \I3.TCNT3_376\ : MUX2H
      port map(A => \I3.TCNT3l3r_net_1\, B => \I3.TCNT3_n3_net_1\, 
        S => \TICKl1r\, Y => \I3.TCNT3_376_net_1\);
    
    \I3.un6_asb_NE\ : NOR3FTT
      port map(A => \I3.un6_asb_NE_adt_net_135785_\, B => 
        \I3.N_260_i_0\, C => \I3.N_186_i_0\, Y => 
        \I3.un6_asb_NE_net_1\);
    
    \I2.PIPE8_DT_545\ : MUX2L
      port map(A => \I2.PIPE8_DTl17r_net_1\, B => 
        \I2.PIPE8_DT_21l17r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_545_net_1\);
    
    \I1.REG_74_0_iv_0l360r\ : AO21
      port map(A => \REGl360r\, B => \I1.N_661\, C => 
        \I1.REG_74l360r_adt_net_114869_\, Y => \I1.REG_74l360r\);
    
    \I3.REG_1_151\ : MUX2L
      port map(A => VDB_inl2r, B => REGl50r, S => 
        \I3.N_1935_adt_net_855332__net_1\, Y => \I3.REG_1_151_0\);
    
    \I2.BNCID_VECT_tile_DOUTl2r\ : MUX2L
      port map(A => \I2.DIN_REG1_0l2r\, B => \I2.DOUT_TMP_0l2r\, 
        S => \I2.N_13\, Y => \I2.BNCID_VECTrxl2r\);
    
    \I3.REGMAP_I_0_IL36R_2982\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un161_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL36R_529\);
    
    \I1.REG_0_sqmuxa_i_0_a4_1_906\ : NAND2
      port map(A => \I1.N_598_23\, B => 
        \I1.sstate_ns_il5r_adt_net_107266_\, Y => 
        \I1.N_435_1_284\);
    
    \I2.END_EVNT2\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT1_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT2_net_1\);
    
    \I2.PIPE10_DT_611\ : MUX2L
      port map(A => \I2.PIPE10_DTl6r_net_1\, B => 
        \I2.PIPE9_DTl6r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_611_net_1\);
    
    \I2.PLL_sram_del.Core\ : PLLCORE
      port map(SDOUT => OPEN, SCLK => \GND\, SDIN => \GND\, 
        SSHIFT => \GND\, SUPDATE => \GND\, GLB => \I2.CLK_sram\, 
        CLK => CLK_c, GLA => OPEN, CLKA => \GND\, LOCK => 
        \I2.PLL_LOCK_sram\, MODE => \GND\, FBDIV5 => \GND\, EXTFB
         => \GND\, FBSEL0 => \GND\, FBSEL1 => \VCC\, FINDIV0 => 
        \GND\, FINDIV1 => \GND\, FINDIV2 => \GND\, FINDIV3 => 
        \GND\, FINDIV4 => \GND\, FBDIV0 => \GND\, FBDIV1 => \GND\, 
        FBDIV2 => \GND\, FBDIV3 => \GND\, FBDIV4 => \GND\, 
        STATBSEL => \GND\, DLYB0 => \GND\, DLYB1 => \GND\, OBDIV0
         => \GND\, OBDIV1 => \GND\, STATASEL => \GND\, DLYA0 => 
        \GND\, DLYA1 => \GND\, OADIV0 => \GND\, OADIV1 => \GND\, 
        OAMUX0 => \GND\, OAMUX1 => \GND\, OBMUX0 => \GND\, OBMUX1
         => \GND\, OBMUX2 => \VCC\, FBDLY0 => \VCC\, FBDLY1 => 
        \VCC\, FBDLY2 => \VCC\, FBDLY3 => \VCC\, XDLYSEL => \VCC\);
    
    \I2.PIPE1_DTl4r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_731_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl4r_net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__3077\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__831\);
    
    \I3.VDBi_57_0_iv_0l19r\ : OR2
      port map(A => \I3.VDBi_57l19r_adt_net_139392_\, B => 
        \I3.VDBi_57l19r_adt_net_139393_\, Y => \I3.VDBi_57l19r\);
    
    \I2.PIPE6_DT_0_sqmuxa_i_o4\ : OR2
      port map(A => \I2.N_4551_adt_net_63758_\, B => 
        \I2.N_4551_adt_net_63759_\, Y => \I2.N_4551\);
    
    \I2.PIPE4_DTl3r_adt_net_854544_\ : BFR
      port map(A => \I2.PIPE4_DTl3r_adt_net_854548__net_1\, Y => 
        \I2.PIPE4_DTl3r_adt_net_854544__net_1\);
    
    ADE_padl12r : OB33PH
      port map(PAD => ADE(12), A => ADE_cl12r);
    
    \I1.REG_74_0_ivl236r\ : AO21
      port map(A => \REGl236r\, B => \I1.N_105\, C => 
        \I1.REG_74l236r_adt_net_127108_\, Y => 
        \I1.REG_74l236r_net_1\);
    
    \I2.WR_SRAM_2_adt_net_748_\ : OAI21FTF
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__149\, B => 
        \I2.N_4030\, C => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_20049__net_1\, Y => 
        \I2.WR_SRAM_2_adt_net_748__net_1\);
    
    \I2.DTO_16_1_IV_0L21R_1112\ : AND2
      port map(A => \I2.DTO_1l21r\, B => \I2.N_196_51\, Y => 
        \I2.DTO_16_1l21r_adt_net_30538_\);
    
    \I2.DT_TEMP_7l7r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, B => 
        \I2.DT_SRAMl7r_net_1\, Y => \I2.DT_TEMP_7l7r_net_1\);
    
    \I1.REG_1_225\ : MUX2H
      port map(A => \REGl324r\, B => \I1.REG_74l324r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y
         => \I1.REG_1_225_net_1\);
    
    \I1.REG_74_0_IVL170R_2064\ : AND2
      port map(A => \FBOUTl5r\, B => 
        \I1.REG_1_sqmuxa_adt_net_855388__net_1\, Y => 
        \I1.REG_74l170r_adt_net_133235_\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I109_Y_1662\ : AOI21
      port map(A => \I2.I109_un1_Y_adt_net_70914_\, B => 
        \I2.N330\, C => \I2.ADD_18x18_fast_I109_Y_0\, Y => 
        \I2.N439_i_adt_net_71055_\);
    
    TDCDB_padl30r : IB33
      port map(PAD => TDCDB(30), Y => TDCDB_cl30r);
    
    \I3.VDBI_57_IV_0_0L6R_2237\ : AO21
      port map(A => \I3.N_2034_adt_net_854684__net_1\, B => 
        \I3.RAMDTSl6r_net_1\, C => 
        \I3.VDBi_57l6r_adt_net_143401_\, Y => 
        \I3.VDBi_57l6r_adt_net_143402_\);
    
    \I3.PIPEA_8l2r\ : AND2
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854464__net_1\, B => 
        \I3.N_211\, Y => \I3.PIPEA_8l2r_net_1\);
    
    \I2.STATE2_NS_I_0L0R_1010\ : AND2FT
      port map(A => \I2.N_176_i_adt_net_855708__net_1\, B => 
        \I2.N_4284\, Y => \I2.N_2796_i_0_adt_net_21575_\);
    
    \I1.REG_74_0_ivl288r\ : AO21
      port map(A => \REGl288r\, B => \I1.N_161\, C => 
        \I1.REG_74l288r_adt_net_122033_\, Y => \I1.REG_74l288r\);
    
    \I2.CRC32_12_i_x2l8r\ : XOR2FT
      port map(A => \I2.CRC32l8r_net_1\, B => \I2.N_3956_i_i\, Y
         => \I2.N_117_i_i_0\);
    
    \I2.DTO_9_IVL3R_1202\ : NOR2
      port map(A => \I2.N_4283_I_0_235\, B => 
        \I2.DT_TEMPl3r_net_1\, Y => 
        \I2.DTO_9_ivl3r_adt_net_34552_\);
    
    \I2.PIPE1_DTl23r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_750_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl23r_net_1\);
    
    REGl404r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_305_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl404r\);
    
    \I2.ROFFSET_c2\ : AND3
      port map(A => \I2.ROFFSETL0R_505\, B => \I2.ROFFSETL1R_506\, 
        C => \I2.ROFFSETL2R_400\, Y => \I2.ROFFSET_c2_net_1\);
    
    \I3.VDBOFFB_30_IV_0L7R_2353\ : AND2
      port map(A => \REGl348r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        Y => \I3.VDBoffb_30l7r_adt_net_161764_\);
    
    \I2.PIPE4_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl16r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl16r_net_1\);
    
    \I5.sstate1se_13_0\ : AO21
      port map(A => TICKL0R_3, B => 
        \I5.sstate1_ns_el0r_adt_net_7898_\, C => 
        \I5.sstate1_ns_el0r_adt_net_8036_\, Y => 
        \I5.sstate1_ns_el0r\);
    
    \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772_\ : BFR
      port map(A => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855772__net_1\);
    
    \I3.REGMAPl28r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un121_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl28r_net_1\);
    
    \I2.CRC32_12_il18r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_52_i_0_i_0\, Y => 
        \I2.N_3935\);
    
    \I2.CRC32_7l3r\ : XOR2
      port map(A => \I2.CRC32l3r_net_1\, B => 
        \I2.DT_TEMPl3r_net_1\, Y => \I2.CRC32_7l3r_net_1\);
    
    \I2.I_1339_G_1\ : XOR2FT
      port map(A => \I2.OFFSETL4R_676\, B => \I2.SUB8L7R_705\, Y
         => \I2.G_1_2\);
    
    \I2.DTO_16_1_IV_0L7R_1185\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855680__net_1\, B => 
        \I2.DTO_9l7r\, Y => \I2.DTO_16_1l7r_adt_net_33720_\);
    
    \I2.PIPE7_DTl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl28r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl28r_net_1\);
    
    \I2.MIC_ERR_REGS_343\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl15r_net_1\, B => 
        \I2.MIC_ERR_REGSl14r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\, Y => 
        \I2.MIC_ERR_REGS_343_net_1\);
    
    \I2.DTE_1l24r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l24r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l24r_Rd1__net_1\);
    
    NLD_pad : OB33PH
      port map(PAD => NLD, A => NLD_c);
    
    \I2.EVNT_WORDl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_722_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl9r_net_1\);
    
    \I2.RAMADl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.RAMAD_4l15r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => RAMAD_cl15r);
    
    \I2.PIPE7_DTL27R_2790\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_83\);
    
    \I1.REG_1_194\ : MUX2H
      port map(A => \REGl293r\, B => \I1.REG_74l293r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\, Y => 
        \I1.REG_1_194_net_1\);
    
    \I3.PIPEA1_300\ : MUX2L
      port map(A => \I3.PIPEA1l2r_net_1\, B => 
        \I3.PIPEA1_12l2r_net_1\, S => 
        \I3.un1_STATE2_15_1_adt_net_1342__net_1\, Y => 
        \I3.PIPEA1_300_net_1\);
    
    \I2.PIPE6_DTl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_464_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl10r_net_1\);
    
    REGl202r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_103_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl202r\);
    
    \I3.CYCS\ : DFFC
      port map(CLK => CLK_c, D => \I3.CYCSF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.CYCS_net_1\);
    
    \I2.ROFFSET_n4\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855704__net_1\, B => 
        \I2.ROFFSET_n4_tz_i\, Y => \I2.ROFFSET_n4_net_1\);
    
    \I2.PIPE8_DT_16_0l0r\ : MUX2H
      port map(A => \I2.PIPE8_DTl0r_net_1\, B => 
        \I2.PIPE7_DTl0r_net_1\, S => 
        \I2.N_565_0_adt_net_855728__net_1\, Y => \I2.N_566\);
    
    \I2.SUB8_1_sqmuxa_0_adt_net_855148_\ : BFR
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855152__net_1\, Y
         => \I2.SUB8_1_sqmuxa_0_adt_net_855148__net_1\);
    
    \I3.PULSE_330_2098\ : AND2
      port map(A => \PULSEl0r_adt_net_854532__net_1\, B => 
        \I3.N_1409\, Y => \I3.PULSE_330_adt_net_134909_\);
    
    \I2.CRC32_12_0_0_m2l29r\ : MUX2L
      port map(A => \I2.DT_TEMPl29r_net_1\, B => 
        \I2.DT_SRAMl29r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854188__net_1\, Y => 
        \I2.N_4157_i_i\);
    
    \I1.REG_74_0_IVL323R_1893\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l323r_adt_net_118787_\);
    
    \I2.PIPE4_DTL9R_3083\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL9R_847\);
    
    \I3.VDBi_31_i_a3_0_1l5r\ : NOR3FFT
      port map(A => REGl53r, B => 
        \I3.REGMAPl9r_adt_net_854328__net_1\, C => 
        \I3.REGMAPL14R_735\, Y => 
        \I3.VDBi_31_i_a3_0_1l5r_adt_net_143649_\);
    
    \I2.I_1340_ca_0_and2\ : AND2FT
      port map(A => \I2.OFFSETl5r_net_1\, B => \I2.SUB8l8r_net_1\, 
        Y => \I2.N_3543_i_i\);
    
    \I1.BYTECNT_n7_i_0_o2_0\ : NAND2
      port map(A => \I1.BYTECNTl7r_net_1\, B => \I1.N_358\, Y => 
        \I1.N_363\);
    
    \I3.VADm_0_a3l16r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl16r_net_1\, Y => \I3.VADml16r\);
    
    \I2.STATE1l7r_1525\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.STATE1_nsl11r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE1L7R_632\);
    
    \I1.N_50_0_adt_net_1409__adt_net_855528_\ : BFR
      port map(A => \I1.N_50_0_ADT_NET_1409__281\, Y => 
        \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\);
    
    \I3.VDBI_57_0_IVL12R_2207\ : AO21
      port map(A => \I3.STATE1_ipl2r_net_1\, B => 
        \I3.VDBi_55l12r_net_1\, C => 
        \I3.VDBi_57l12r_adt_net_140997_\, Y => 
        \I3.VDBi_57l12r_adt_net_140998_\);
    
    \I2.CHAINB_EN244_c_0_adt_net_855248_\ : BFR
      port map(A => \I2.CHAINB_EN244_c_0\, Y => 
        \I2.CHAINB_EN244_c_0_adt_net_855248__net_1\);
    
    \I1.REG_14_sqmuxa_adt_net_855436_\ : BFR
      port map(A => \I1.REG_14_sqmuxa\, Y => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\);
    
    \I2.OFFSET_37_3l7r\ : MUX2L
      port map(A => \I2.N_650\, B => \I2.N_642\, S => 
        \I2.PIPE7_DTL26R_349\, Y => \I2.N_658\);
    
    DTE_padl11r : IOB33PH
      port map(PAD => DTE(11), A => \I2.DTE_1l11r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl11r);
    
    \I2.BNC_IDl4r_1605\ : DFFB
      port map(CLK => CLK_c, D => \I2.I_20_0\, CLR => 
        \I2.N_4627_i_0\, SET => \I2.N_4607_i_0\, Q => 
        \I2.BNC_IDL4R_712\);
    
    \I3.UN15_ANYCYC_2297\ : NOR3FFT
      port map(A => \I3.PIPEBl28r_net_1\, B => 
        \I3.un15_anycyc_adt_net_147620_\, C => 
        \I3.PIPEB_i_0_il31r\, Y => 
        \I3.un15_anycyc_adt_net_147613_\);
    
    \I2.UN21_SRAM_EMPTY_NE_1037\ : NOR2
      port map(A => \I2.un21_sram_empty_3_net_1\, B => 
        \I2.un21_sram_empty_2_net_1\, Y => 
        \I2.un21_sram_empty_NE_adt_net_24173_\);
    
    \I2.SUB8l11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_514_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l11r_net_1\);
    
    \I2.DTO_1_888\ : MUX2L
      port map(A => \I2.DTO_1l14r_Rd1__net_1\, B => 
        \I2.DTO_16_1l14r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834768_Rd1__net_1\, Y
         => \I2.DTO_1l14r\);
    
    \I2.DTO_16_1_IV_0_0L12R_1158\ : AND2
      port map(A => \I2.N_182_ADT_NET_1007__385\, B => 
        \I2.DT_SRAMl12r_net_1\, Y => 
        \I2.DTO_16_1l12r_adt_net_32624_\);
    
    REGl168r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_69_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl168r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I139_Y_i\ : AO21FTF
      port map(A => \I2.N_96_0_adt_net_58152_\, B => 
        \I2.N_40_0_adt_net_577252_\, C => \I2.N_91_0\, Y => 
        \I2.N_42_1\);
    
    \I2.PIPE10_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_624_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl19r_net_1\);
    
    \I2.SUB8_523_2706\ : NOR3FTT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855136__net_1\, B
         => \I2.SUB_21x21_fast_I216_Y_0\, C => 
        \I2.N475_adt_net_87372_\, Y => 
        \I2.SUB8_523_adt_net_566476_\);
    
    \I2.OFFSET_37_4l3r\ : MUX2L
      port map(A => \REGl368r\, B => \REGl304r\, S => 
        \I2.PIPE7_DTL27R_71\, Y => \I2.N_662\);
    
    \I2.FID_7_0_IVL9R_1714\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl9r_net_1\, 
        Y => \I2.FID_7l9r_adt_net_92645_\);
    
    \I2.INT_ERRS\ : OR3
      port map(A => \I2.INT_ERRS_adt_net_22801_\, B => 
        \I2.INT_ERRBS_i_i\, C => \I2.INT_ERRAS_net_1\, Y => 
        \I2.INT_ERRS_net_1\);
    
    \I5.SSTATE1SE_7_0_0_904\ : AND3
      port map(A => TICKL0R_558, B => \I5.sstate1l3r_net_1\, C
         => \I5.N_67\, Y => \I5.sstate1_ns_el8r_adt_net_8886_\);
    
    REGl309r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_210_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl309r\);
    
    \I2.PIPE4_DTl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl11r_net_1\);
    
    \I2.CRC32_12_0_0_x2l24r\ : XOR2FT
      port map(A => \I2.CRC32l24r_net_1\, B => \I2.N_4270_i_i\, Y
         => \I2.N_128_i_0_i_0\);
    
    \I1.REG_74L404R_1784\ : AOI21TTF
      port map(A => \I1.PAGECNTl7r_net_1\, B => 
        \I1.REG_74_1_404_m7_i_a5_0_net_1\, C => 
        \I1.REG_74_1_396_N_12\, Y => \I1.N_273_adt_net_109616_\);
    
    \I3.VDBOFFA_31_IV_0L3R_2575\ : AO21
      port map(A => \REGl256r\, B => \I3.REGMAPl29r_net_1\, C => 
        \I3.VDBoffa_31l3r_adt_net_164040_\, Y => 
        \I3.VDBoffa_31l3r_adt_net_164072_\);
    
    \I2.TDCDASl30r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl30r, Q => 
        \I2.TDCDASl30r_net_1\);
    
    \I3.RAMAD_VME_29\ : MUX2H
      port map(A => RAMAD_VMEl5r, B => \I3.VASl6r_net_1\, S => 
        \I3.TCNT_0_sqmuxa\, Y => \I3.RAMAD_VME_29_net_1\);
    
    \I2.PIPE6_DT_470\ : MUX2H
      port map(A => \I2.PIPE5_DTl16r_net_1\, B => 
        \I2.PIPE6_DTl16r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_470_net_1\);
    
    REGl246r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_147_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl246r\);
    
    \I2.N_4541_i_0_o2\ : NOR2
      port map(A => \I2.PIPE5_DTL23R_623\, B => 
        \I2.PIPE5_DTL21R_625\, Y => \I2.N_217\);
    
    \I1.REG_74_0_IVL294R_1924\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l294r_adt_net_121384_\);
    
    \I2.LEAD_FLAG6_7_i_0l3r\ : AOI21
      port map(A => \I2.N_4673\, B => \I2.N_484\, C => \I2.N_222\, 
        Y => \I2.N_4532_adt_net_64252_\);
    
    \I3.REG_1_274\ : MUX2H
      port map(A => VDB_inl2r, B => \I3.REGl93r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_274_0\);
    
    \I3.REG_1l110r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_291_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl110r);
    
    \I2.DTESl8r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl8r, Q => 
        \I2.DTESl8r_net_1\);
    
    \I2.REG_0l3r_adt_net_848_\ : AO21
      port map(A => \I3.REG1l3r_net_1\, B => \I3.REG2l3r_net_1\, 
        C => \I2.REG_0l3r_adt_net_19773_Rd1__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__net_1\);
    
    \I3.PIPEA_242\ : MUX2L
      port map(A => \I3.PIPEAl11r_net_1\, B => 
        \I3.PIPEA_8l11r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854672__net_1\, Y
         => \I3.PIPEA_242_net_1\);
    
    \I2.PIPE8_DT_543\ : MUX2L
      port map(A => \I2.PIPE8_DTl15r_net_1\, B => 
        \I2.PIPE8_DT_21l15r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_543_net_1\);
    
    \I3.REG3l7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG3_132_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l7r_net_1\);
    
    \I4.resyn_0_I4_un1_bcnt_2\ : NAND3FFT
      port map(A => \I4.N_48_3_adt_net_14719_\, B => 
        \I4.bcntl0r_net_1\, C => \I4.bcntl3r_net_1\, Y => 
        \I4.N_48_3\);
    
    \I5.SCL_63\ : MUX2H
      port map(A => \I5.SCL_net_1\, B => \I5.N_484\, S => TICKl0r, 
        Y => \I5.SCL_63_net_1\);
    
    \I2.LSRAM_INl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_384_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl0r_net_1\);
    
    DTO_padl17r : IOB33PH
      port map(PAD => DTO(17), A => \I2.DTO_1l17r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl17r);
    
    \I3.NOEDTKi_111\ : OAI21FTF
      port map(A => NOEDTK_C_14, B => \I3.un1_NOEDTKi_0_sqmuxa_1\, 
        C => \I3.un1_NOEDTKi_0_sqmuxa\, Y => 
        \I3.NOEDTKi_111_net_1\);
    
    \I1.REG_74L388R_1804\ : OR3
      port map(A => \I1.REG_30_sqmuxa_adt_net_854376__net_1\, B
         => \I1.N_257_adt_net_111267_\, C => \I1.REG_27_sqmuxa\, 
        Y => \I1.N_257_adt_net_111279_\);
    
    \I3.DSS_1163\ : DFFS
      port map(CLK => CLK_c, D => \I3.DSSF1_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.DSS_425\);
    
    \I2.SRAM_EVNT_n1_0\ : XOR2FT
      port map(A => \I2.SRAM_EVNTl1r_net_1\, B => \I2.N_128_1\, Y
         => \I2.SRAM_EVNT_n1_0_net_1\);
    
    \I2.SUB8_1_sqmuxa_0_a2_0_0\ : NOR2
      port map(A => \I2.NWPIPE7_689\, B => 
        \I2.N_587_adt_net_1201__net_1\, Y => \I2.SUB8_1_sqmuxa_0\);
    
    \I3.REG_1_ml79r\ : AND2
      port map(A => REGl79r, B => 
        \I3.REGMAPl9r_adt_net_854324__net_1\, Y => 
        \I3.VDBi_20l31r\);
    
    \I2.PIPE1_DT_42_1_IVL7R_1479\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        B => \I2.PIPE1_DT_12l7r_net_1\, Y => 
        \I2.PIPE1_DT_42l7r_adt_net_50677_\);
    
    \I2.ENDF\ : DFFC
      port map(CLK => CLK_c, D => \I2.ENDF_712_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ENDF_net_1\);
    
    \I2.FID_7_0_IVL13R_965\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl13r_net_1\, 
        Y => \I2.FID_7l13r_adt_net_18081_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I197_Y\ : XOR2FT
      port map(A => \I2.N411_adt_net_194931__net_1\, B => 
        \I2.SUB_21x21_fast_I197_Y_0\, Y => \I2.SUB8_2l1r\);
    
    \I2.OFFSET_37_29l4r\ : MUX2L
      port map(A => \I2.N_855\, B => \I2.N_743\, S => 
        \I2.CHA_DATA8_net_1\, Y => \I2.OFFSET_37l4r\);
    
    \I3.un111_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_586\, B => \I3.N_553\, Y => 
        \I3.un111_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.OFFSET_37_25l0r\ : MUX2L
      port map(A => \REGl253r\, B => \REGl189r\, S => 
        \I2.PIPE7_DTL27R_88\, Y => \I2.N_827\);
    
    \I3.VDBi_31l30r\ : MUX2L
      port map(A => \I3.REGl163r\, B => \I3.VDBi_20l30r\, S => 
        \I3.REGMAPl17r_adt_net_854280__net_1\, Y => 
        \I3.VDBi_31l30r_net_1\);
    
    \I5.SCLA_i_a2\ : OR2
      port map(A => \I5.SCL_net_1\, B => \I5.CHAIN_SELECT_net_1\, 
        Y => \I5.N_107\);
    
    \I2.LSRAM_IN_391\ : MUX2L
      port map(A => \I2.PIPE5_DTl7r_net_1\, B => 
        \I2.LSRAM_INl7r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_391_net_1\);
    
    REGl358r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_259_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl358r\);
    
    \I2.ROFFSET_n0\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855700__net_1\, B => 
        \I2.ROFFSETl0r_net_1\, Y => \I2.ROFFSET_n0_net_1\);
    
    \I1.REG_1_251\ : MUX2H
      port map(A => \REGl350r\, B => \I1.REG_74l350r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_251_net_1\);
    
    \I2.DT_SRAM_0l12r\ : MUX2L
      port map(A => \I2.PIPE10_DTl12r_net_1\, B => 
        \I2.PIPE5_DTl12r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854212__net_1\, Y => 
        \I2.N_880\);
    
    \I1.PAGECNTl6r_adt_net_854928_\ : BFR
      port map(A => \I1.PAGECNTl6r_adt_net_854932__net_1\, Y => 
        \I1.PAGECNTl6r_adt_net_854928__net_1\);
    
    \I3.VDBi_40l9r\ : MUX2L
      port map(A => \I3.N_347\, B => \I3.N_1854\, S => 
        \I3.N_354_0_adt_net_855368__net_1\, Y => 
        \I3.VDBi_40l9r_net_1\);
    
    \I1.REG_21_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_260_222\, B => \I1.N_243\, Y => 
        \I1.REG_21_sqmuxa\);
    
    \I1.REG_74_0_ivl352r\ : AO21
      port map(A => \REGl352r\, B => \I1.N_225\, C => 
        \I1.REG_74l352r_adt_net_115945_\, Y => \I1.REG_74l352r\);
    
    \I1.REG_74_0_IVL310R_1906\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_19_sqmuxa_adt_net_855488__net_1\, Y => 
        \I1.REG_74l310r_adt_net_119905_\);
    
    \I2.TDCDASl10r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl10r, Q => 
        \I2.TDCDASl10r_net_1\);
    
    \I3.STATE1_tr22_17_0_i2_0_a2_i_o3_0_o3\ : NAND2
      port map(A => \I3.N_277\, B => \I3.STATE1_IPL9R_731\, Y => 
        \I3.N_303\);
    
    \I2.REG_1_c8_i\ : AOI21FTT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => \I2.N_3852\, C => \I2.N_129\, Y => \I2.N_3837_i_0\);
    
    \I5.SSTATE1SE_0_0_0_909\ : AND3FFT
      port map(A => \I5.N_64_adt_net_855868__net_1\, B => 
        \I5.COMMANDl0r_net_1\, C => 
        \I5.sstate1_ns_el1r_adt_net_9246_\, Y => 
        \I5.sstate1_ns_el1r_adt_net_9243_\);
    
    \I2.DT_SRAM_i_m_0l28r\ : NOR2FT
      port map(A => \I2.N_182_ADT_NET_1007__385\, B => 
        \I2.DT_SRAMl28r_net_1\, Y => \I2.DT_SRAM_i_m_0l28r_net_1\);
    
    \I3.VDBoffb_30_iv_0l7r\ : AND2
      port map(A => \REGl372r\, B => \I3.REGMAPl43r_net_1\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161744_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I203_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl7r\, B => 
        \I2.PIPE7_DTl7r_net_1\, Y => \I2.SUB_21x21_fast_I203_Y_0\);
    
    \I2.STATE3_nsl12r\ : AO21
      port map(A => \I2.STATE3l1r_net_1\, B => \I2.N_3015\, C => 
        \I2.STATE3_nsl12r_adt_net_24672_\, Y => 
        \I2.STATE3_nsl12r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I208_Y\ : XOR2
      port map(A => \I2.N495_i\, B => 
        \I2.SUB_21x21_fast_I208_Y_0\, Y => \I2.SUB8_2l12r\);
    
    \I2.PIPE1_DT_30l9r\ : MUX2L
      port map(A => \I2.TDCDBSl9r_net_1\, B => 
        \I2.TDCDBSl7r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, Y
         => \I2.PIPE1_DT_30l9r_net_1\);
    
    \I2.TOKENB_CNTl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TOKENB_CNT_3l1r\, CLR => 
        \I2.un12_clear_stat_i\, Q => \I2.TOKENB_CNTl1r_net_1\);
    
    \I3.REG_1_280\ : MUX2H
      port map(A => VDB_inl8r, B => \I3.REGl99r\, S => 
        \I3.N_2297_i\, Y => \I3.REG_1_280_0\);
    
    \I2.CRC32_12_0l1r\ : MUX2L
      port map(A => \I2.CRC32_7_il1r\, B => \I2.CRC32_2_il1r\, S
         => \I2.N_4667_1_adt_net_1046__adt_net_854424__net_1\, Y
         => \I2.N_999\);
    
    \I2.ENDF_1140_1731\ : DFFC
      port map(CLK => CLK_c, D => \I2.ENDF_712_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ENDF_838\);
    
    \I1.REG_30_sqmuxa_adt_net_854376_\ : BFR
      port map(A => \I1.REG_30_sqmuxa\, Y => 
        \I1.REG_30_sqmuxa_adt_net_854376__net_1\);
    
    \I2.DTE_21_1_IV_0L5R_1328\ : OR3
      port map(A => \I2.DTO_16_1l5r_adt_net_34192_\, B => 
        \I2.DTE_21_1l5r_adt_net_39091_\, C => 
        \I2.DTE_21_1l5r_adt_net_39098_\, Y => 
        \I2.DTE_21_1l5r_adt_net_39100_\);
    
    REGl231r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_132_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl231r\);
    
    \I3.VDBOFFA_47_2582\ : AND2
      port map(A => \I3.un1_REGMAP_30_adt_net_855008__net_1\, B
         => \I3.VDBoffal3r_net_1\, Y => 
        \I3.VDBoffa_47_adt_net_164118_\);
    
    \I3.VDBi_40_0_i_m2l3r\ : MUX2L
      port map(A => REGl421r, B => REGl437r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_135\);
    
    \I3.END_PK_1773\ : DFFC
      port map(CLK => CLK_c, D => \I3.END_PK_229_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.END_PK_879\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I163_un1_Y\ : AND3
      port map(A => \I2.N516\, B => \I2.N350\, C => 
        \I2.N504_adt_net_88887_\, Y => \I2.I163_un1_Y\);
    
    \I5.SDANOE_8_0_916\ : NOR3FFT
      port map(A => \I5.N_64_adt_net_855868__net_1\, B => 
        \I5.SDAnoe_8_adt_net_9738_\, C => \I5.N_74\, Y => 
        \I5.SDAnoe_8_adt_net_9739_\);
    
    \I3.PIPEA1_12l1r\ : AND2
      port map(A => DPR_cl1r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, Y => 
        \I3.PIPEA1_12l1r_net_1\);
    
    \I2.TRGARRl0r\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.DWACT_ADD_CI_0_partial_sum_2l0r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.TRGARRl0r_net_1\);
    
    \I2.DTE_cl_0_sqmuxa_2_0_a2_0_a2_0_908\ : OR2FT
      port map(A => \I2.N_4241_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, Y => 
        \I2.DTE_CL_0_SQMUXA_2_0_286\);
    
    \I2.PIPE1_DT_42_1_IVL2R_1511\ : OAI21TTF
      port map(A => GA_cl2r, B => \I2.N_3238\, C => 
        \I2.PIPE1_DT_42l2r_adt_net_51836_\, Y => 
        \I2.PIPE1_DT_42l2r_adt_net_51837_\);
    
    \I3.REG_1_201\ : MUX2L
      port map(A => VDB_inl20r, B => \I3.REGl153r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\, Y => 
        \I3.REG_1_201_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I15_G0N_i_o4\ : NAND2
      port map(A => \I2.RAMDT4L5R_818\, B => 
        \I2.PIPE4_DTl15r_net_1\, Y => \I2.N_8\);
    
    \I2.STATE1_NS_I_0L13R_1017\ : OA21
      port map(A => \I2.N_3272\, B => \I2.N_3351\, C => 
        \I2.STATE1l5r_net_1\, Y => \I2.N_3214_i_0_adt_net_22011_\);
    
    \I2.WOFFSETl10r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl10r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl10r_Rd1__net_1\);
    
    \I1.REG_74_0_IV_0_0L260R_1965\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.N_596\, Y => 
        \I1.REG_74l260r_adt_net_124798_\);
    
    \I3.UN1_REGMAP_30_0_A2_2083\ : NOR2
      port map(A => \I3.REGMAPL20R_780\, B => \I3.REGMAPL21R_779\, 
        Y => \I3.un1_REGMAP_30_adt_net_134453_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I138_Y_0_o2_2\ : AOI21
      port map(A => \I2.PIPE4_DTL10R_475\, B => 
        \I2.PIPE4_DTL11R_841\, C => \I2.RAMDT4L5R_811\, Y => 
        \I2.N_80\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I137_Y_I_2709\ : NOR3FFT
      port map(A => \I2.N_40_0_adt_net_58199_\, B => 
        \I2.N_40_0_adt_net_577252_\, C => 
        \I2.N_96_0_adt_net_58152_\, Y => 
        \I2.N_40_0_adt_net_577295_\);
    
    \I2.un8_evread_0_a2_1\ : OR2FT
      port map(A => \I2.FIFO_END_EVNT_579\, B => EVREAD_562, Y
         => \I2.un8_evread_1\);
    
    \I2.CRC32_799\ : MUX2L
      port map(A => \I2.CRC32l4r_net_1\, B => \I2.N_3921\, S => 
        \I2.N_2826_1_adt_net_794__net_1\, Y => 
        \I2.CRC32_799_net_1\);
    
    \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892_\ : BFR
      port map(A => \I3.N_1906_i_0_0_adt_net_855636__net_1\, Y
         => 
        \I3.N_1906_i_0_0_adt_net_855636__adt_net_855892__net_1\);
    
    \I3.PIPEA1_12l26r\ : AND2
      port map(A => DPR_cl26r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854488__net_1\, Y => 
        \I3.PIPEA1_12l26r_net_1\);
    
    \I1.REG_74_2_4l228r\ : OR3
      port map(A => \I1.REG_74_1_380_m8_i_0_Rd1__net_1\, B => 
        \I1.REG_74_2_4_il228r_adt_net_115255_\, C => 
        \I1.REG_74_2_4_il228r_adt_net_115250_\, Y => 
        \I1.REG_74_2_4_il228r\);
    
    \I3.REG_1_192\ : MUX2L
      port map(A => VDB_inl11r, B => \I3.REGl144r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, Y => 
        \I3.REG_1_192_0\);
    
    \I1.PAGECNT_318\ : MUX2H
      port map(A => \I1.PAGECNTl9r_net_1\, B => \I1.N_1380\, S
         => \I1.PAGECNTe_adt_net_854896__net_1\, Y => 
        \I1.PAGECNT_318_net_1\);
    
    \I5.BITCNT_n2_i_o4\ : AND2
      port map(A => \I5.BITCNT_C0_573\, B => \I5.BITCNTl1r_net_1\, 
        Y => \I5.N_65\);
    
    \I2.EVNT_NUM_c2\ : AND2
      port map(A => \I2.EVNT_NUML2R_596\, B => 
        \I2.EVNT_NUM_c1_net_1\, Y => \I2.EVNT_NUM_c2_net_1\);
    
    \I3.REG_44_il84r\ : AND2
      port map(A => \I3.REG_1_sqmuxa_3_adt_net_855340__net_1\, B
         => \I3.N_1630_adt_net_150503_\, Y => \I3.N_1630\);
    
    \I3.VDBI_40_0L5R_2243\ : AND2FT
      port map(A => \I3.N_354_0_adt_net_855372__net_1\, B => 
        \I3.N_137\, Y => \I3.VDBi_40l5r_adt_net_143744_\);
    
    \I3.REG_1_196\ : MUX2L
      port map(A => VDB_inl15r, B => \I3.REGl148r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\, Y => 
        \I3.REG_1_196_0\);
    
    \I2.PIPE8_DT_16l14r\ : AND2
      port map(A => 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\, B => 
        \I2.N_580\, Y => \I2.PIPE8_DT_16l14r_net_1\);
    
    \I3.STATE1_ns_0_iv_0l4r\ : AO21FTT
      port map(A => \I3.DSS_net_1\, B => \I3.STATE1_ipl6r\, C => 
        \I3.N_1516\, Y => \I3.STATE1_nsl4r\);
    
    \I2.N_4646_1_ADT_NET_1645_RD1__2750\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_ADT_NET_1645_RD1__26\);
    
    \I1.REG_1_151\ : MUX2H
      port map(A => \REGl250r\, B => \I1.REG_74l250r\, S => 
        \I1.N_50_0_ADT_NET_1409__293\, Y => \I1.REG_1_151_net_1\);
    
    \I2.PIPE1_DT_748\ : MUX2L
      port map(A => \I2.PIPE1_DTl21r_net_1\, B => 
        \I2.PIPE1_DT_42l21r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854568__net_1\, 
        Y => \I2.PIPE1_DT_748_net_1\);
    
    \I3.un191_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_586\, Y => 
        \I3.un191_reg_ads_0_a2_0_a3_net_1\);
    
    FBOUTl5r : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_63_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \FBOUTl5r\);
    
    REGl266r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_167_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl266r\);
    
    \I1.REG_74_0_ivl291r\ : AO21
      port map(A => \REGl291r\, B => \I1.N_161\, C => 
        \I1.REG_74l291r_adt_net_121775_\, Y => \I1.REG_74l291r\);
    
    \I3.STATE1_nsl2r_adt_net_1586_\ : AO21TTF
      port map(A => \I3.un1_REGMAP_30\, B => 
        \I3.STATE1_nsl2r_adt_net_134736__net_1\, C => 
        \I3.WRITES_8\, Y => \I3.STATE1_nsl2r_adt_net_1586__net_1\);
    
    \I1.REG_74_0_IVL229R_1997\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_9_sqmuxa_adt_net_854728__net_1\, Y => 
        \I1.REG_74l229r_adt_net_127710_\);
    
    \I1.REG_74_0_iv_0_0l252r\ : AO21
      port map(A => \REGl252r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l252r_adt_net_125605_\, Y => \I1.REG_74l252r\);
    
    \I2.un1_DTO_cl_1_sqmuxa_2_0_o2_1_0_x2_779\ : XOR2FT
      port map(A => NOESRAME_C_241, B => 
        \I2.WOFFSETl0r_adt_net_854644__net_1\, Y => 
        \I2.N_176_I_157\);
    
    \I1.REG_1_210\ : MUX2H
      port map(A => \REGl309r\, B => \I1.REG_74l309r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_210_net_1\);
    
    \I2.PIPE10_DT_612\ : MUX2L
      port map(A => \I2.PIPE10_DTl7r_net_1\, B => 
        \I2.PIPE9_DTl7r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_612_net_1\);
    
    \I1.REG_74_0_IVL358R_1849\ : AND2
      port map(A => \FBOUTl1r\, B => \I1.REG_25_sqmuxa\, Y => 
        \I1.REG_74l358r_adt_net_115041_\);
    
    VDB_padl6r : IOB33PH
      port map(PAD => VDB(6), A => \I3.VDBml6r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl6r);
    
    \I2.RAMDT4l2r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl2r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l2r_net_1\);
    
    \I2.N475_adt_net_442371_\ : AND3
      port map(A => \I2.N285\, B => \I2.N479_adt_net_642172_\, C
         => \I2.N479_adt_net_642225_\, Y => 
        \I2.N475_adt_net_442371__net_1\);
    
    \I2.PIPE9_DTl16r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_285_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl16r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL29R_1358\ : AO21
      port map(A => \I2.PIPE1_DT_2_SQMUXA_1_1_177\, B => 
        \I2.TDCDBSl29r_net_1\, C => 
        \I2.PIPE1_DT_42l29r_adt_net_45835_\, Y => 
        \I2.PIPE1_DT_42l29r_adt_net_45837_\);
    
    \I2.PIPE4_DTl17r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl17r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl17r_net_1\);
    
    \I1.REG_74_0_IVL190R_2044\ : AND2
      port map(A => \FBOUTl1r\, B => \I1.REG_4_sqmuxa\, Y => 
        \I1.REG_74l190r_adt_net_131441_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I8_P0N_i_a2\ : OR2
      port map(A => \I2.RAMDT4L5R_137\, B => 
        \I2.PIPE4_DTl8r_adt_net_854556__net_1\, Y => \I2.N_95\);
    
    \I3.STATE1_ns_0_iv_0_0_a3l6r\ : AND2FT
      port map(A => \I3.DSS_net_1\, B => \I3.N_1920\, Y => 
        \I3.STATE1_nsl6r\);
    
    ADE_padl15r : OB33PH
      port map(PAD => ADE(15), A => ADE_cl15r);
    
    \I2.DTO_16_1_IV_0_0L29R_1072\ : AND2FT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        B => \I2.DT_TEMPl29r_net_1\, Y => 
        \I2.DTO_16_1l29r_adt_net_28732_\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854468_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854472__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854468__net_1\);
    
    \I4.un1_lead_flag_1_1_0\ : MUX2L
      port map(A => LEAD_FLAGl4r, B => LEAD_FLAGl0r, S => 
        \I4.bcnt_i_0_il2r_net_1\, Y => \I4.N_1\);
    
    \I1.LOAD_RESi\ : DFFC
      port map(CLK => CLK_c, D => \I1.LOAD_RESi_50_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => LOAD_RES);
    
    \I2.N_4246_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4246\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4246_Rd1__net_1\);
    
    \I2.MIC_ERR_REGS_342\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl14r_net_1\, B => 
        \I2.MIC_ERR_REGSl13r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855856__net_1\, Y => 
        \I2.MIC_ERR_REGS_342_net_1\);
    
    \I1.REG_74_0_IVL296R_1922\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_17_sqmuxa_adt_net_855480__net_1\, Y => 
        \I1.REG_74l296r_adt_net_121212_\);
    
    \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820_\ : BFR
      port map(A => \I2.un1_STATE3_10_1_adt_net_999__net_1\, Y
         => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\);
    
    \I1.REG_74_2_I_A2_0L404R_1813\ : OR3
      port map(A => PULSEL0R_756, B => 
        \I1.REG_74_12_300_N_13_Rd1__net_1\, C => 
        \I1.REG_74_4_I_A2_404_N_4_I_ADT_NET_1465__193\, Y => 
        \I1.N_1366_adt_net_112007_\);
    
    \I3.STATE1_NS_0_IV_0L1R_2079\ : AO21FTT
      port map(A => \I3.N_268\, B => \I3.STATE1_ipl9r\, C => 
        \I3.STATE1_nsl1r_adt_net_134330_\, Y => 
        \I3.STATE1_nsl1r_adt_net_134337_\);
    
    \I3.VDBOFFA_31_IV_0L2R_2585\ : AND2
      port map(A => \REGl247r\, B => \I3.REGMAPl28r_net_1\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164226_\);
    
    \I2.REG_1_n12\ : XOR2
      port map(A => \I2.N_3840\, B => \I2.REG_1_n12_0_net_1\, Y
         => \I2.REG_1_n12_net_1\);
    
    \I2.BNCID_VECTrff_9\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_9_256_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_9\);
    
    \I2.RAMDT4L5R_2811\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_139\);
    
    \I2.FID_7_IVL3R_1726\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl3r_net_1\, 
        Y => \I2.FID_7l3r_adt_net_93251_\);
    
    \I1.REG_74_0_IVL393R_1797\ : NOR2FT
      port map(A => \FBOUTl4r\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, Y => 
        \I1.REG_74l393r_adt_net_110784_\);
    
    \I3.VDBOFFA_31_IV_0L2R_2589\ : AO21
      port map(A => \REGl199r\, B => \I3.REGMAPl22r_net_1\, C => 
        \I3.VDBoffa_31l2r_adt_net_164214_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164258_\);
    
    \I2.PIPE8_DT_21l17r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl17r\, B => 
        \I2.PIPE8_DT_16l17r_net_1\, S => \I2.NWPIPE7_net_1\, Y
         => \I2.PIPE8_DT_21l17r_net_1\);
    
    \I2.PIPE7_DTL27R_2772\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_65\);
    
    \I1.REG_74_0_IVL336R_1880\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\, Y => 
        \I1.REG_74l336r_adt_net_117572_\);
    
    REGl271r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_172_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl271r\);
    
    \I2.FIRST_TDC_1_sqmuxa\ : NOR2FT
      port map(A => \I2.PIPE1_DT_2_SQMUXA_1_1_177\, B => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855076__net_1\, Y
         => \I2.FIRST_TDC_1_sqmuxa_net_1\);
    
    \I2.MIC_REG2l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG2_311_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2l2r_net_1\);
    
    \I3.un51_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_573\, B => 
        \I3.un41_reg_ads_0_a2_3_a3_0\, Y => 
        \I3.un51_reg_ads_0_a2_0_a3_net_1\);
    
    \I1.LUT_0_sqmuxa_i_0_o2_i_0_834\ : NOR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__186\, B
         => \I1.N_325_499\, Y => \I1.N_328_I_0_212\);
    
    \I3.STATE2_ns_o2l3r\ : NOR2
      port map(A => \I3.ADACKCYC_net_1\, B => \I3.N_281\, Y => 
        \I3.N_1465\);
    
    \I1.REG_1_213\ : MUX2H
      port map(A => \REGl312r\, B => \I1.REG_74l312r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_213_net_1\);
    
    \I2.DTO_cl_0_sqmuxa_0_adt_net_855196_\ : BFR
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855200__net_1\, 
        Y => \I2.DTO_cl_0_sqmuxa_0_adt_net_855196__net_1\);
    
    \I4.STATE1_nsl1r\ : NOR2
      port map(A => \I4.STATE1_nsl2r\, B => 
        \I4.STATE1_nsl0r_net_1\, Y => \I4.STATE1_nsl1r_net_1\);
    
    \I2.DT_TEMP_7l24r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854236__net_1\, B => 
        \I2.N_4194\, Y => \I2.DT_TEMP_7l24r_net_1\);
    
    \I2.PIPE1_DTl30r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_757_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl30r_net_1\);
    
    \I2.DTO_1l16r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_1l16r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_1l16r_Rd1__net_1\);
    
    DTO_pad_i_1l31r : AND2
      port map(A => \I2.DTO_cl_32l31r\, B => \I2.DTO_cll31r\, Y
         => \I2.N_4239_i_0_1\);
    
    \I3.RAMDTSl9r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl9r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl9r_net_1\);
    
    \I3.STATE1l9r_1771\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl1r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL9R_877\);
    
    \I1.sstate_tr18_0_a2_0_a4_945\ : AND2FT
      port map(A => \I1.COMMAND_716\, B => \I1.LUT_net_1\, Y => 
        \I1.SSTATE_NS_IL5R_ADT_NET_107266__323\);
    
    \I1.REG_74l284r\ : OR2FT
      port map(A => \I1.REG_16_sqmuxa\, B => 
        \I1.N_161_adt_net_1449__net_1\, Y => \I1.N_153\);
    
    \I3.STATE1_IPL2R_3099\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl8r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL2R_885\);
    
    \I1.N_50_0_ADT_NET_1409__2872\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__541\, B => 
        \I1.N_50_0_ADT_NET_109751__257\, Y => 
        \I1.N_50_0_ADT_NET_1409__294\);
    
    \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854612_\ : BFR
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854620__net_1\, 
        Y => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854612__net_1\);
    
    \I2.DT_TEMP_7l23r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854236__net_1\, B => 
        \I2.DT_SRAMl23r_net_1\, Y => \I2.DT_TEMP_7l23r_net_1\);
    
    \I1.ISI_0_sqmuxa_1_0_i_a2\ : OR3FTT
      port map(A => \I1.sstatel9r_net_1\, B => \I1.N_321\, C => 
        \I1.sstatel0r_net_1\, Y => \I1.N_653\);
    
    \I2.OFFSET_37_3l2r\ : MUX2L
      port map(A => \I2.N_645\, B => \I2.N_637\, S => 
        \I2.PIPE7_DTL26R_350\, Y => \I2.N_653\);
    
    REGl282r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_183_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl282r\);
    
    \I1.PAGECNTl2r_adt_net_834908_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.PAGECNT_325_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNTl2r_adt_net_834908_Rd1__net_1\);
    
    \I2.SRAM_EVNT_C3_I_1746\ : NOR3
      port map(A => \I2.SRAM_EVNTl2r_net_1\, B => 
        \I2.SRAM_EVNTl3r_net_1\, C => \I2.N_135\, Y => 
        \I2.N_3828_adt_net_101749_\);
    
    \I1.REG_74_0_IV_0L176R_2058\ : AND2
      port map(A => \REGl176r\, B => \I1.N_49_267\, Y => 
        \I1.REG_74l176r_adt_net_132682_\);
    
    \I1.REG_74_0_ivl339r\ : AO21
      port map(A => \REGl339r\, B => \I1.N_209\, C => 
        \I1.REG_74l339r_adt_net_117314_\, Y => \I1.REG_74l339r\);
    
    \I2.EVNT_NUM_n2\ : NOR2
      port map(A => EV_RES_C_569, B => \I2.EVNT_NUM_n2_tz_i\, Y
         => \I2.EVNT_NUM_n2_net_1\);
    
    \I3.N_1409_adt_net_854744_\ : BFR
      port map(A => \I3.N_1409\, Y => 
        \I3.N_1409_adt_net_854744__net_1\);
    
    \I2.PIPE7_DTL27R_2797\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_90\);
    
    \I2.PIPE5_DT_6l13r\ : MUX2L
      port map(A => \I2.PIPE4_DTl13r_net_1\, B => \I2.N_1082\, S
         => \I2.N_4547_1_adt_net_1209__adt_net_855608__net_1\, Y
         => \I2.PIPE5_DT_6l13r_net_1\);
    
    \I2.LEAD_FLAG6_644\ : AO21
      port map(A => \I2.N_4528_adt_net_1129__net_1\, B => 
        \I2.N_4528_adt_net_63525_\, C => 
        \I2.LEAD_FLAG6_644_adt_net_63844_\, Y => 
        \I2.LEAD_FLAG6_644_net_1\);
    
    \I4.FLUSH\ : DFFC
      port map(CLK => CLK_c, D => \I4.FLUSH_3_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FLUSH);
    
    \I2.CRC32_12_IL3R_1350\ : OA21FTF
      port map(A => 
        \I2.N_4667_1_adt_net_1046__adt_net_854424__net_1\, B => 
        \I2.CRC32_7l3r_net_1\, C => 
        \I2.N_2867_1_adt_net_854960__net_1\, Y => 
        \I2.N_3920_adt_net_43068_\);
    
    \I3.TCNT3_375\ : MUX2H
      port map(A => \I3.TCNT3_i_0_il4r_net_1\, B => 
        \I3.TCNT3_n4_net_1\, S => \TICKl1r\, Y => 
        \I3.TCNT3_375_net_1\);
    
    \I3.VDBi_29_0l9r\ : MUX2L
      port map(A => \I3.REGl100r\, B => 
        \I3.VDBi_29l9r_adt_net_1596__net_1\, S => 
        \I3.REGMAPl14r_net_1\, Y => \I3.VDBi_29l9r\);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854668_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854668__net_1\);
    
    \I2.PIPE4_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl30r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl30r_net_1\);
    
    \I1.REG_1_279\ : MUX2H
      port map(A => \REGl378r\, B => \I1.REG_74l378r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_279_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I10_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L12R_828\, B => 
        \I2.PIPE4_DTL10R_791\, Y => \I2.N_59_0\);
    
    \I2.PIPE2_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl0r_net_1\);
    
    \I3.VDBoff_120\ : MUX2L
      port map(A => \I3.VDBoffl4r_net_1\, B => \I3.N_2068\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_120_net_1\);
    
    \I5.AIR_WDATAl9r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_59_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl9r_net_1\);
    
    \I2.N_2826_1_ADT_NET_794__2890\ : OAI21FTF
      port map(A => \I2.N_4261_304\, B => \I2.N_4282\, C => 
        \I2.N_2826_1_adt_net_40744__net_1\, Y => 
        \I2.N_2826_1_ADT_NET_794__331\);
    
    GA_padl3r : IB33
      port map(PAD => GA(3), Y => GA_cl3r);
    
    \I2.WOFFSET_13_il1r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_5_0\, Y => 
        \I2.N_4244\);
    
    \I2.LSRAM_IN_393\ : MUX2L
      port map(A => \I2.PIPE5_DTl9r_net_1\, B => 
        \I2.LSRAM_INl9r_net_1\, S => \I2.LEAD_FLAG6_0_sqmuxa_1_1\, 
        Y => \I2.LSRAM_IN_393_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I9_G0N_0_o3\ : AND2
      port map(A => \I2.RAMDT4L12R_826\, B => 
        \I2.PIPE4_DTL9R_790\, Y => \I2.N_16_0\);
    
    \I1.BITCNT_n2_i_i_o2\ : AND2
      port map(A => \I1.BITCNTL0R_18\, B => \I1.BITCNTl1r_net_1\, 
        Y => \I1.N_324\);
    
    \I2.MIC_ERR_REGSl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_340_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl11r_net_1\);
    
    \I3.VDBi_40_0_i_m2l0r\ : MUX2L
      port map(A => REGl418r, B => REGl434r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_132\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_A2_1_2666\ : AND2
      port map(A => \I2.RAMDT4L4R_883\, B => \I2.PIPE4_DTL4R_478\, 
        Y => \I2.N_107_adt_net_276024_\);
    
    \I3.VDBm_0l11r\ : MUX2L
      port map(A => \I3.PIPEAl11r_net_1\, B => 
        \I3.PIPEBl11r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_153\);
    
    REGl389r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_290_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl389r\);
    
    \I2.SUB8_520\ : AND2
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855160__net_1\, B
         => \I2.SUB_21x21_fast_I213_Y_0\, Y => 
        \I2.SUB8_520_adt_net_531295_\);
    
    \I2.DTO_16_1_iv_0l7r\ : OR2
      port map(A => \I2.DTO_16_1l7r_adt_net_33735_\, B => 
        \I2.DTO_16_1l7r_adt_net_33736_\, Y => \I2.DTO_16_1l7r\);
    
    \I2.PIPE8_DT_21l27r\ : MUX2H
      port map(A => \I2.PIPE7_DTl27r_net_1\, B => 
        \I2.LSRAM_OUTl27r\, S => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l27r_net_1\);
    
    \I1.REG_1_134\ : MUX2H
      port map(A => \REGl233r\, B => \I1.REG_74l233r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\, Y => 
        \I1.REG_1_134_net_1\);
    
    \I3.REGMAPl21r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un86_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl21r_net_1\);
    
    \I2.WROi_10_0_0_o2\ : OA21FTF
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.N_2838_i_0\, C => \I2.N_2867_1_adt_net_854960__net_1\, 
        Y => \I2.N_2836\);
    
    \I1.PAGECNTl0r_adt_net_833884_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I1.PAGECNT_327_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.PAGECNTl0r_adt_net_833884_Rd1__net_1\);
    
    \I5.REG_1l445r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_28_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl445r);
    
    \I3.VDBOFFB_30_IV_0L4R_2414\ : AO21
      port map(A => \REGl313r\, B => \I3.REGMAP_i_0_il36r_net_1\, 
        C => \I3.VDBoffb_30l4r_adt_net_162334_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162363_\);
    
    \I3.PIPEA1_315\ : MUX2L
      port map(A => \I3.PIPEA1l17r_net_1\, B => 
        \I3.PIPEA1_12l17r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__252\, Y => 
        \I3.PIPEA1_315_net_1\);
    
    \I1.N_238_Rd1__adt_net_854884_\ : BFR
      port map(A => \I1.N_238_Rd1__adt_net_854888__net_1\, Y => 
        \I1.N_238_Rd1__adt_net_854884__net_1\);
    
    \I3.PIPEB_91\ : AO21
      port map(A => DPR_cl12r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_91_adt_net_160209_\, Y => 
        \I3.PIPEB_91_net_1\);
    
    \I2.L2SERVl3r_1260\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_919_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL15R_522\);
    
    \I2.DTE_21_1_ivl2r\ : AOI21FTT
      port map(A => \I2.DTE_1l2r_net_1\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\, C => 
        \I2.DTE_21_1_iv_2_il2r\, Y => \I2.DTE_21_1_iv_i_0l2r\);
    
    \I2.SUB9_1_ADD_18x18_fast_I29_Y\ : AO21TTF
      port map(A => \I2.SUB8l14r_net_1\, B => \I2.SUB8l13r_net_1\, 
        C => \I2.N291_adt_net_4302__net_1\, Y => \I2.N294\);
    
    \I1.PAGECNT_n6_i_i_a2_853\ : AND2FT
      port map(A => \I1.PAGECNTL6R_248\, B => \I1.PAGECNTL5R_308\, 
        Y => \I1.N_590_231\);
    
    \I5.SBYTE_67\ : MUX2H
      port map(A => \I5.SBYTEl2r_net_1\, B => \I5.N_18\, S => 
        \I5.N_406\, Y => \I5.SBYTE_67_net_1\);
    
    \I0.HWCLEARi\ : DFFC
      port map(CLK => CLK_c, D => PLL_LOCK, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => HWCLEAR);
    
    \I3.un13_reg_ads_0_a2_0_a3\ : NOR2FT
      port map(A => \I3.un221_reg_ads_0_a2_0_a3_adt_net_165933_\, 
        B => \I3.N_637\, Y => \I3.un13_reg_ads_0_a2_0_a3_net_1\);
    
    \I1.REG_74_I_O2L364R_1842\ : OR3FTT
      port map(A => \I1.REG_29_sqmuxa\, B => 
        \I1.N_661_adt_net_114478_\, C => 
        \I1.N_661_adt_net_114476_\, Y => 
        \I1.N_661_adt_net_114485_\);
    
    \I1.REG_74_0_ivl361r\ : AO21
      port map(A => \REGl361r\, B => \I1.N_661\, C => 
        \I1.REG_74l361r_adt_net_114783_\, Y => \I1.REG_74l361r\);
    
    TDCDA_padl11r : IB33
      port map(PAD => TDCDA(11), Y => TDCDA_cl11r);
    
    \I2.PIPE1_DT_42_1_IV_2L26R_1370\ : OAI21FTF
      port map(A => \I2.PIPE1_DT_2_SQMUXA_1_1_177\, B => 
        \I2.TDCDBSl26r_net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46167_\, Y => 
        \I2.PIPE1_DT_42_1_iv_2_il26r_adt_net_46179_\);
    
    \I2.OFFSET_37_5l5r\ : MUX2L
      port map(A => \REGl402r\, B => \REGl338r\, S => 
        \I2.PIPE7_DTL27R_78\, Y => \I2.N_672\);
    
    \I1.sstatel4r_1608\ : DFFC
      port map(CLK => CLK_c, D => \I1.sstate_nsl6r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.SSTATEL4R_715\);
    
    \I2.UN1_END_CHAINA1_0_SQMUXA_I_O3_1535\ : NOR2
      port map(A => \I2.N_3351\, B => \I2.N_3275\, Y => 
        \I2.N_3281_adt_net_53327_\);
    
    \I2.DTE_21_1_IV_0L24R_1248\ : AO21
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.DTO_9l24r\, C
         => \I2.DTE_21_1l24r_adt_net_37174_\, Y => 
        \I2.DTE_21_1l24r_adt_net_37175_\);
    
    \I2.ROFFSETl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_910_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl8r_net_1\);
    
    \I5.COMMANDl0r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_12_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl0r_net_1\);
    
    \I2.LSRAM_INl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_399_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl15r_net_1\);
    
    \I2.PIPE8_DT_21_i_a2l31r\ : OR2
      port map(A => \I2.NWPIPE7_689\, B => 
        \I2.PIPE7_DTl31r_net_1\, Y => \I2.N_4418\);
    
    \I2.WOFFSET_13_il9r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_52\, Y => \I2.N_4252\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I122_Y_0_o2\ : OAI21FTT
      port map(A => \I2.N_64_0_adt_net_855028__net_1\, B => 
        \I2.N_17_0\, C => \I2.N_67\, Y => \I2.N_84_0\);
    
    \I2.DTO_16_1l18r_adt_net_756_\ : MUX2L
      port map(A => \I2.N_202_i\, B => \I2.PIPE2_DTl18r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.DTO_16_1l18r_adt_net_756__net_1\);
    
    \I2.OFFSET_37_10l6r\ : MUX2L
      port map(A => \I2.N_705\, B => \I2.N_697\, S => 
        \I2.PIPE7_DTL26R_352\, Y => \I2.N_713\);
    
    \I2.FID_7_0_IVL29R_977\ : AND2
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl29r_net_1\, 
        Y => \I2.FID_7l29r_adt_net_18645_\);
    
    \I1.REG_1_276\ : MUX2H
      port map(A => \REGl375r\, B => \I1.REG_74l375r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_276_net_1\);
    
    \I2.WOFFSET_13_il8r\ : AND2
      port map(A => \I2.N_4262\, B => \I2.I_45\, Y => \I2.N_4251\);
    
    \I1.REG_74_0_IVL285R_1934\ : NOR2FT
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_16_sqmuxa_adt_net_855456__net_1\, Y => 
        \I1.REG_74l285r_adt_net_122291_\);
    
    \I1.N_50_0_ADT_NET_109751__2861\ : NOR3FFT
      port map(A => \I1.N_232_1\, B => 
        \I1.N_50_0_adt_net_109760__net_1\, C => \I1.N_435_1_283\, 
        Y => \I1.N_50_0_ADT_NET_109751__256\);
    
    \I3.PIPEB_83\ : AO21
      port map(A => DPR_cl4r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_83_adt_net_160545_\, Y => 
        \I3.PIPEB_83_net_1\);
    
    \I1.LUT_0_sqmuxa_i_0_o2_i_0_833\ : NOR2FT
      port map(A => \I1.PAGECNT_0L9R_ADT_NET_835128_RD1__186\, B
         => \I1.N_325\, Y => \I1.N_328_I_0_211\);
    
    \I3.VDBi_369\ : MUX2L
      port map(A => \I3.VDBil29r_net_1\, B => \I3.VDBi_57l29r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_369_net_1\);
    
    \I2.FID_7_IVL4R_1723\ : AND2
      port map(A => \I2.STATE3L2R_413\, B => \I2.DTOSl4r_net_1\, 
        Y => \I2.FID_7l4r_adt_net_93151_\);
    
    \I2.PIPE1_DT_735\ : MUX2L
      port map(A => \I2.PIPE1_DTl8r_net_1\, B => 
        \I2.PIPE1_DT_42l8r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854580__net_1\, 
        Y => \I2.PIPE1_DT_735_net_1\);
    
    \I2.RAMDT4L5R_3067\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_821\);
    
    \I1.REG_74_0_iv_0l275r\ : AO21
      port map(A => \REGl275r\, B => 
        \I1.N_145_adt_net_854768__net_1\, C => 
        \I1.REG_74l275r_adt_net_123388_\, Y => \I1.REG_74l275r\);
    
    \I3.PIPEA1l28r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEA1_326_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l28r_net_1\);
    
    \I1.REG_74_0_iv_0l180r\ : AO21
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_2_sqmuxa_adt_net_855392__net_1\, C => 
        \I1.REG_74l180r_adt_net_132338_\, Y => 
        \I1.REG_74l180r_net_1\);
    
    \I5.COMMANDl15r\ : DFFC
      port map(CLK => CLK_c, D => \I5.COMMAND_52_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.COMMANDl15r_net_1\);
    
    \I2.L2TYPE_4_IL8R_1627\ : OR2FT
      port map(A => \I2.N_4458\, B => \I2.N_4459\, Y => 
        \I2.N_4444_adt_net_67711_\);
    
    \I2.MIC_ERR_REGSl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_356_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl27r_net_1\);
    
    \I2.DTO_16_1_IV_1L1R_1210\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855692__net_1\, B => 
        \I2.DTO_9_ivl1r_net_1\, C => 
        \I2.DTO_16_1_iv_1l1r_adt_net_35122_\, Y => 
        \I2.DTO_16_1_iv_1l1r_adt_net_35128_\);
    
    \I2.DTO_16_1_IV_0L13R_1152\ : AND2
      port map(A => \I2.N_4671_adt_net_854596__net_1\, B => 
        \I2.DT_TEMPl13r_net_1\, Y => 
        \I2.DTO_16_1l13r_adt_net_32384_\);
    
    LED_R_pad : OB33PH
      port map(PAD => LED_R, A => LED_R_i_a3);
    
    TDCDA_padl7r : IB33
      port map(PAD => TDCDA(7), Y => TDCDA_cl7r);
    
    REGl304r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_205_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl304r\);
    
    \I2.MTDCRESA_378\ : OR3
      port map(A => MTDCRESA_c, B => \I2.TOKENA_TIMOUT_net_1\, C
         => PULSEl8r, Y => \I2.MTDCRESA_378_net_1\);
    
    \I3.DSS_0_1611\ : DFFS
      port map(CLK => CLK_c, D => \I3.DSSF1_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.DSS_718\);
    
    \I2.PIPE8_DT_21_0L29R_1672\ : AO21FTT
      port map(A => \I2.PIPE7_DTl31r_net_1\, B => 
        \I2.PIPE7_DTl29r_net_1\, C => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l29r_adt_net_82644_\);
    
    \I5.sstate1se_2_0\ : AO21FTT
      port map(A => TICKl0r, B => \I5.sstate1l10r_net_1\, C => 
        \I5.sstate1_ns_el3r_adt_net_9195_\, Y => 
        \I5.sstate1_ns_el3r\);
    
    \I3.VDBI_29L3R_2718\ : MUX2L
      port map(A => \I3.REGl94r\, B => 
        \I3.VDBi_20l3r_adt_net_144750_\, S => \I3.REGMAPL14R_734\, 
        Y => \I3.VDBi_29l3r_adt_net_618363_\);
    
    \I2.PIPE4_DTL10R_3086\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL10R_850\);
    
    \I2.L2SERVl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_921_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEl13r\);
    
    \I5.DATAl14r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l14r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl131r);
    
    \I3.VADm_0_a3l14r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl14r_net_1\, Y => \I3.VADml14r\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I142_Y_0_A2_3_1557\ : OR2
      port map(A => \I2.PIPE4_DTL8R_483\, B => 
        \I2.PIPE4_DTL7R_482\, Y => \I2.N_139_0_adt_net_55124_\);
    
    \I3.MBLTCYC\ : DFFC
      port map(CLK => CLK_c, D => \I3.MBLTCYC_114_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.MBLTCYC_net_1\);
    
    \I1.REG_74_0_ivl193r\ : AO21
      port map(A => \REGl193r\, B => \I1.N_65\, C => 
        \I1.REG_74l193r_adt_net_131183_\, Y => \I1.REG_74l193r\);
    
    \I2.PIPE10_DT_17_il13r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l0r_net_1\, C => \I2.PIPE10_DT_17_i_0l13r_net_1\, 
        Y => \I2.N_3799\);
    
    \I2.BNCID_VECTrff_5_260_0\ : AO21
      port map(A => \I2.BNCID_VECTwa13_1_net_1\, B => 
        \I2.BNCID_VECTrff_7_258_0_a2_0\, C => \I2.BNCID_VECTro_5\, 
        Y => \I2.BNCID_VECTrff_5_260_0_net_1\);
    
    \I1.REG_74_0_iv_0_0l249r\ : AO21
      port map(A => \REGl249r\, B => 
        \I1.REG_74_0_iv_0_o2_245_N_9_i_0\, C => 
        \I1.REG_74l249r_adt_net_125863_\, Y => \I1.REG_74l249r\);
    
    REGl226r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_127_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl226r\);
    
    \I3.REG_1_185\ : MUX2L
      port map(A => VDB_inl4r, B => \I3.REGl137r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855308__net_1\, Y => 
        \I3.REG_1_185_0\);
    
    \I3.REGMAPL47R_2931\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un216_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL47R_448\);
    
    \I2.ROFFSETl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_912_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl6r_net_1\);
    
    \I5.AIR_WDATA_58\ : MUX2H
      port map(A => \I5.N_463\, B => \I5.AIR_WDATAl8r_net_1\, S
         => \I5.N_461\, Y => \I5.AIR_WDATA_58_net_1\);
    
    \I1.REG_74_0l356r\ : NOR3FFT
      port map(A => \I1.N_273_10\, B => 
        \I1.REG_74_12_348_m9_i_net_1\, C => \I1.N_273_11_i\, Y
         => \I1.REG_74_0l348r\);
    
    \I2.DTOSl15r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl15r, Q => 
        \I2.DTOSl15r_net_1\);
    
    AMB_padl2r : IB33
      port map(PAD => AMB(2), Y => AMB_cl2r);
    
    \I2.un3_hwres\ : OR2
      port map(A => \HWRES_3_ADT_NET_738__17\, B => PULSEL5R_16, 
        Y => \I2.un3_hwres_i\);
    
    \I3.REGMAPl35r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un156_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl35r_net_1\);
    
    \I2.BNCID_VECTrff_4_261_0\ : AO21
      port map(A => \I2.BNCID_VECTwa12_1_net_1\, B => 
        \I2.BNCID_VECTrff_7_258_0_a2_0\, C => \I2.BNCID_VECTro_4\, 
        Y => \I2.BNCID_VECTrff_4_261_0_net_1\);
    
    \I2.FID_7_IVL2R_1730\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl50r, C => 
        \I2.STATE3l9r_net_1\, Y => \I2.FID_7l2r_adt_net_93358_\);
    
    \I2.PIPE1_DT_42_1_IVL1R_1515\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        B => \I2.PIPE1_DT_12l1r_net_1\, Y => 
        \I2.PIPE1_DT_42l1r_adt_net_52031_\);
    
    \I2.DTO_9_ivl30r\ : OA21TTF
      port map(A => \I2.N_4283_i_0_adt_net_854972__net_1\, B => 
        \I2.DT_TEMPl30r_net_1\, C => \I2.DT_SRAM_i_ml30r_net_1\, 
        Y => \I2.DTO_9_ivl30r_net_1\);
    
    \I2.DTESl9r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl9r, Q => 
        \I2.DTESl9r_net_1\);
    
    \I2.STATE2l4r_adt_net_855684_\ : BFR
      port map(A => \I2.STATE2l4r_net_1\, Y => 
        \I2.STATE2l4r_adt_net_855684__net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I190_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl20r_net_1\, Y => 
        \I2.ADD_21x21_fast_I190_Y_0\);
    
    \I2.DTO_16_1_iv_0l21r\ : OR2
      port map(A => \I2.DTO_16_1l21r_adt_net_30547_\, B => 
        \I2.DTO_16_1l21r_adt_net_30548_\, Y => \I2.DTO_16_1l21r\);
    
    \I3.UN1_REGMAP_30_0_A2_0_2082\ : NOR2
      port map(A => \I3.REGMAP_I_0_IL32R_774\, B => 
        \I3.REGMAPL31R_773\, Y => 
        \I3.un1_REGMAP_30_0_a2_0_adt_net_134424_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I153_Y_i_a4_0\ : OR2
      port map(A => \I2.N519\, B => \I2.N_86_i_adt_net_57123_\, Y
         => \I2.N_86_i\);
    
    \I1.BYTECNT_n1_i_0_x2\ : XOR2FT
      port map(A => \I1.BYTECNT_i_0_il1r_net_1\, B => 
        \I1.BYTECNTl0r_net_1\, Y => \I1.N_386_i_i_0\);
    
    \I0.EV_RESi_1462\ : DFFC
      port map(CLK => CLK_c, D => \I0.EV_RESi_1_net_1\, CLR => 
        \I0.un4_hwresi_i\, Q => EV_RES_C_569);
    
    \I2.PIPE5_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_698_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl22r_net_1\);
    
    \I1.N_41_9_adt_net_854784_\ : BFR
      port map(A => \I1.N_41_9\, Y => 
        \I1.N_41_9_adt_net_854784__net_1\);
    
    \I2.DTO_16_1_IVL14R_1150\ : AO21
      port map(A => \I2.N_182_adt_net_1007__net_1\, B => 
        \I2.DT_SRAMl14r_net_1\, C => 
        \I2.DTO_16_1l14r_adt_net_32208_\, Y => 
        \I2.DTO_16_1l14r_adt_net_32209_\);
    
    \I2.I_1338_ca_0_and2\ : NOR2FT
      port map(A => \I2.SUB8l6r_net_1\, B => \I2.OFFSETl3r_net_1\, 
        Y => \I2.N_3539_i_i\);
    
    \I2.PIPE8_DT_21l11r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl11r\, B => \I2.N_577\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l11r_net_1\);
    
    \I2.PIPE2_DTl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl14r_net_1\);
    
    \I3.PIPEB_94_2329\ : NOR2FT
      port map(A => \I3.PIPEBl15r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_94_adt_net_160083_\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I180_UN1_Y_2660\ : AO21
      port map(A => \I2.N301_2\, B => \I2.N479_adt_net_642225_\, 
        C => \I2.N300_0\, Y => \I2.I180_un1_Y_adt_net_252355_\);
    
    \I1.REG_74l332r\ : NAND2FT
      port map(A => \I1.REG_22_sqmuxa\, B => \I1.REG_74_0l332r\, 
        Y => \I1.N_201\);
    
    \I2.FID_7_0_ivl6r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl6r_net_1\, 
        C => \I2.FID_7l6r_adt_net_92935_\, Y => \I2.FID_7l6r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I120_Y_0\ : AO21
      port map(A => \I2.N_61_0\, B => \I2.N531_0_adt_net_60059_\, 
        C => \I2.N_140_0\, Y => \I2.N531_0\);
    
    \I2.DTO_16_1_IV_0L31R_1067\ : AO21
      port map(A => \I2.DTO_1l31r_net_1\, B => \I2.N_196_52\, C
         => \I2.DTO_16_1l31r_adt_net_28246_\, Y => 
        \I2.DTO_16_1l31r_adt_net_28256_\);
    
    \I2.un21_sram_empty_0\ : XOR2
      port map(A => \I2.RPAGEL12R_608\, B => \I2.L2ARRL0R_602\, Y
         => \I2.un21_sram_empty_0_net_1\);
    
    \I1.REG_1_278\ : MUX2H
      port map(A => \REGl377r\, B => \I1.REG_74l377r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_278_net_1\);
    
    \REG_i_il5r_adt_net_855556_\ : BFR
      port map(A => \REG_i_il5r_adt_net_855560__net_1\, Y => 
        \REG_i_il5r_adt_net_855556__net_1\);
    
    \I1.REG_1_260\ : MUX2H
      port map(A => \REGl359r\, B => \I1.REG_74l359r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_260_net_1\);
    
    \I1.REG_29_sqmuxa_0_a2_1_a2\ : OR3
      port map(A => \I1.REG_74_12_300_N_15_adt_net_3731__net_1\, 
        B => \I1.N_1169_adt_net_854812__net_1\, C => 
        \I1.N_260_220\, Y => \I1.REG_29_sqmuxa\);
    
    FID_padl10r : OB33PH
      port map(PAD => FID(10), A => FID_cl10r);
    
    \I3.VDBil13r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_353_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil13r_net_1\);
    
    \I2.N_3277_i_i_o3\ : OR2
      port map(A => \I2.STATE1l10r_net_1\, B => 
        \I2.STATE1l5r_net_1\, Y => \I2.N_3277\);
    
    \I2.DT_TEMP_7l27r\ : NOR2
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854232__net_1\, B => 
        \I2.N_4647\, Y => \I2.DT_TEMP_7l27r_net_1\);
    
    \I3.un1_evrdy_1_i_s_i_o2l0r\ : AND2
      port map(A => \I3.N_268_259\, B => \I3.REGMAPL0R_722\, Y
         => \I3.N_258\);
    
    \I3.REG_1l60r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_161_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl60r);
    
    \I2.MIC_REG2L3R_ADT_NET_834020_RD1__2974\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.MIC_REG2_312_adt_net_855644__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG2L3R_ADT_NET_834020_RD1__491\);
    
    \I2.BNC_ID_il0r\ : INV
      port map(A => \I2.BNC_IDl0r_net_1\, Y => \I2.BNC_ID_i_0l0r\);
    
    \I3.STATE1_NS_0_IV_0_0L8R_2119\ : NOR2FT
      port map(A => \I3.STATE1_IPL2R_886\, B => 
        \I3.N_57_i_0_0_adt_net_854688__net_1\, Y => 
        \I3.STATE1_nsl8r_adt_net_136092_\);
    
    \I1.REG_74_0_iv_0l215r\ : AO21
      port map(A => \FBOUTl2r\, B => \I1.REG_7_sqmuxa\, C => 
        \I1.REG_74l215r_adt_net_129206_\, Y => \I1.REG_74l215r\);
    
    \I1.REG_23_sqmuxa_0_a2_m2_e\ : AND3FFT
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__adt_net_855536__net_1\, 
        B => \I1.N_127_i\, C => \I1.REG_74_9_0_o4_a0_2l372r\, Y
         => \I1.REG_23_sqmuxa\);
    
    \I3.REG_1_224\ : MUX2L
      port map(A => VDB_inl11r, B => REGl417r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_224_0\);
    
    \I2.PIPE7_DTL27R_2774\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_67\);
    
    \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1_\ : 
        DFFC
      port map(CLK => CLK_c, D => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Ra1__net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__net_1\);
    
    \I2.REG_1_n1\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => \I2.REG_1_n1_0_net_1\, Y => \I2.REG_1_n1_net_1\);
    
    \I2.PIPE8_DT_544\ : MUX2L
      port map(A => \I2.PIPE8_DTl16r_net_1\, B => 
        \I2.PIPE8_DT_21l16r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_544_net_1\);
    
    ADE_padl7r : OB33PH
      port map(PAD => ADE(7), A => ADE_cl7r);
    
    REGl212r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_113_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl212r\);
    
    \I3.REG_1l160r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG_1_208_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl160r\);
    
    \I2.DTO_1_876\ : MUX2L
      port map(A => \I2.DTO_1l2r_net_1\, B => \I2.DTO_16_1_ivl2r\, 
        S => \I2.DTE_0_sqmuxa_i_0_N_3_1\, Y => 
        \I2.DTO_1_876_net_1\);
    
    \I5.REG_1l117r\ : DFFS
      port map(CLK => CLK_c, D => \I5.REG_1_54_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl117r);
    
    TDCDB_padl17r : IB33
      port map(PAD => TDCDB(17), Y => TDCDB_cl17r);
    
    \I2.DTO_16_1_iv_0l5r\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855676__net_1\, B => 
        \I2.DTO_9l5r\, C => \I2.DTO_16_1l5r_adt_net_34200_\, Y
         => \I2.DTO_16_1l5r\);
    
    \I1.REG_74_0_IVL320R_1896\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l320r_adt_net_119045_\);
    
    \I2.DTO_16_1l14r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l14r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l14r_Rd1__net_1\);
    
    \I3.PIPEBl19r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_98_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl19r_net_1\);
    
    \I3.VDBi_55l11r\ : MUX2H
      port map(A => \I3.VDBil11r_net_1\, B => 
        \I3.RAMDTSl11r_net_1\, S => 
        \I3.N_57_i_0_0_adt_net_854692__net_1\, Y => 
        \I3.VDBi_55l11r_net_1\);
    
    \I2.FIFO_END_EVNT_1472\ : DFFC
      port map(CLK => CLK_c, D => \I2.FIFO_END_EVNT_489_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.FIFO_END_EVNT_579\);
    
    \I2.MTDCRESB_379\ : OR3
      port map(A => MTDCRESB_c, B => \I2.TOKENB_TIMOUT_i_i\, C
         => PULSEl9r, Y => \I2.MTDCRESB_379_net_1\);
    
    \I1.REG_1_192\ : MUX2H
      port map(A => \REGl291r\, B => \I1.REG_74l291r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855468__net_1\, Y => 
        \I1.REG_1_192_net_1\);
    
    \I1.ISI\ : DFFC
      port map(CLK => CLK_c, D => \I1.ISI_54_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => F_SI_c);
    
    \I2.SUB9_1_ADD_18X18_FAST_I124_Y_1652\ : OA21TTF
      port map(A => \I2.N_3562_i\, B => \I2.SUB8l19r_net_1\, C
         => \I2.SUB8l20r_net_1\, Y => \I2.N434_adt_net_69831_\);
    
    \I2.PIPE7_DTl1r_1596\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL1R_703\);
    
    \I2.un1_STATE1_38_0_o2\ : AO21
      port map(A => \I2.N_3272\, B => \I2.N_3277\, C => 
        \I2.N_3292_adt_net_52393_\, Y => \I2.N_3292\);
    
    \I2.STATE1l18r_1520\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_o2_0l0r_net_1\, SET => CLEAR_STAT_i_0, Q
         => \I2.STATE1L18R_627\);
    
    \I1.REG_1_263\ : MUX2H
      port map(A => \REGl362r\, B => \I1.REG_74l362r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_263_net_1\);
    
    \I2.WPAGEl15r\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_948_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEl15r_net_1\);
    
    \I2.WOFFSETl0r_adt_net_854636_\ : BFR
      port map(A => \I2.WOFFSETl0r_adt_net_854640__net_1\, Y => 
        \I2.WOFFSETl0r_adt_net_854636__net_1\);
    
    \I5.AIR_WDATA_3_sqmuxa_i\ : NAND2FT
      port map(A => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\, B => 
        \I5.sstate2l1r_net_1\, Y => \I5.N_443\);
    
    \I2.STATE3l3r_1154\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl10r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3L3R_416\);
    
    \I1.SSTATE_NS_1_IV_0_0L7R_1768\ : NOR3
      port map(A => \I1.N_604\, B => \I1.COMMAND_net_1\, C => 
        \I1.LUT_net_1\, Y => \I1.sstate_nsl7r_adt_net_107573_\);
    
    \I3.VDBi_367\ : MUX2L
      port map(A => \I3.VDBil27r_net_1\, B => \I3.VDBi_57l27r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_367_net_1\);
    
    \I2.PIPE8_DT_557\ : MUX2L
      port map(A => \I2.PIPE8_DTl29r_net_1\, B => 
        \I2.PIPE8_DT_21l29r\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_557_net_1\);
    
    \I3.VDBI_29L3R_2719\ : AO21
      port map(A => \I3.VDBi_29l3r_adt_net_510711_\, B => 
        \I3.VDBi_29l3r_adt_net_510792_\, C => 
        \I3.VDBi_29l3r_adt_net_618363_\, Y => 
        \I3.VDBi_29l3r_net_1\);
    
    \I2.PIPE1_DT_42_1_IV_1L25R_1371\ : NOR2
      port map(A => REGl429r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855816__net_1\, Y => 
        \I2.PIPE1_DT_42_1_iv_1_il25r_adt_net_46307_\);
    
    \I2.DTE_21_1_IV_0L9R_1307\ : AO21
      port map(A => \I2.DT_TEMPl9r_net_1\, B => \I2.N_4038\, C
         => \I2.DTE_21_1l9r_adt_net_38621_\, Y => 
        \I2.DTE_21_1l9r_adt_net_38635_\);
    
    \I1.REG_74_i_o2_1_0_364_m5\ : MUX2L
      port map(A => \I1.REG_74_i_o2_1_0_364_N_5\, B => 
        \I1.REG_74_i_o2_1_0_364_N_2\, S => \I1.PAGECNTl9r_net_1\, 
        Y => \I1.REG_74_i_o2_1_0_364_N_6\);
    
    \I2.STATEE_NSL3R_1025\ : AND3FFT
      port map(A => \I2.CHAIN_ERRS_net_1\, B => 
        \I2.INT_ERRS_net_1\, C => \I2.STATEel4r_net_1\, Y => 
        \I2.STATEe_nsl3r_adt_net_22967_\);
    
    REGl319r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_220_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl319r\);
    
    \I3.VDBOFFB_30_IV_0L7R_2351\ : AND2
      port map(A => \REGl292r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161756_\);
    
    \I3.VDBOFFB_30_IV_0L2R_2442\ : AND2
      port map(A => \REGl351r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162710_\);
    
    \I2.un2_evnt_word_I_20\ : XOR2
      port map(A => \I2.N_42\, B => 
        \I2.WOFFSETl4r_adt_net_854980__net_1\, Y => \I2.I_20\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I142_Y_0_a2_1_1006\ : OA21
      port map(A => \I2.N_140_0_ADT_NET_947__328\, B => 
        \I2.N_139_0_adt_net_55124_\, C => \I2.RAMDT4L5R_136\, Y
         => \I2.N_107_ADT_NET_256840__384\);
    
    \I2.DTE_21_1_IV_0L8R_1309\ : AND2
      port map(A => \I2.STATE2l3r_net_1\, B => \I2.N_3967\, Y => 
        \I2.DTE_21_1l8r_adt_net_38735_\);
    
    \I2.resyn_0_I2_FID_428\ : MUX2H
      port map(A => FID_cl12r, B => \I2.FID_7l12r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\, 
        Y => \I2.FID_428\);
    
    \I2.PIPE6_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_478_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl24r_net_1\);
    
    \I2.PIPE8_DT_21l21r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl21r\, B => 
        \I2.PIPE7_DTl21r_net_1\, S => \I2.NWPIPE7_net_1\, Y => 
        \I2.PIPE8_DT_21l21r_net_1\);
    
    \I2.STATE2l4r_adt_net_855680_\ : BFR
      port map(A => \I2.STATE2l4r_adt_net_855684__net_1\, Y => 
        \I2.STATE2l4r_adt_net_855680__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I53_Y\ : NAND2
      port map(A => \I2.N273_546\, B => \I2.N270_0_544\, Y => 
        \I2.N303_0\);
    
    \I2.STATE3l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_nsl8r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3l5r_net_1\);
    
    \I2.L2RF2_i\ : INV
      port map(A => \I2.L2RF2_net_1\, Y => \I2.L2RF2_i_net_1\);
    
    \I3.VDBI_57_0_IV_0_0L8R_2220\ : AO21
      port map(A => REGl125r, B => \I3.N_2058\, C => 
        \I3.VDBi_57l8r_adt_net_142723_\, Y => 
        \I3.VDBi_57l8r_adt_net_142678_\);
    
    \I2.OFFSET_37_20l6r\ : MUX2L
      port map(A => \I2.N_785\, B => \I2.N_777\, S => 
        \I2.PIPE7_DTL26R_356\, Y => \I2.N_793\);
    
    \I2.STATE4_ns_a3_il0r\ : NOR2
      port map(A => \I2.STATE4l1r_net_1\, B => \I2.N_3376_1\, Y
         => \I2.STATE4_ns_a3_il0r_net_1\);
    
    \I2.DTESl1r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl1r, Q => 
        \I2.DTESl1r_net_1\);
    
    \I2.DT_TEMPl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_782_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl21r_net_1\);
    
    \I2.L2TYPEl9r_1551\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_598_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPE_I_0_IL9R_658\);
    
    \I2.TDCDBSl3r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl3r, Q => 
        \I2.TDCDBSl3r_net_1\);
    
    \I2.PIPE10_DT_17_il20r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l7r_net_1\, C => \I2.PIPE10_DT_17_i_0l20r_net_1\, 
        Y => \I2.N_3806\);
    
    \I2.PIPE1_DT_42_1_IV_1L25R_1372\ : OAI21TTF
      port map(A => REGl445r, B => \I2.N_3234\, C => 
        \I2.PIPE1_DT_42_1_iv_1_il25r_adt_net_46307_\, Y => 
        \I2.PIPE1_DT_42_1_iv_1_il25r_adt_net_46311_\);
    
    \I2.DTO_16_1l9r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l9r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l9r_Rd1__net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__2993\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__540\);
    
    \I2.L2TYPE_4_i_o2l7r\ : AND2FT
      port map(A => \I2.N_4454\, B => \I2.N_4460\, Y => 
        \I2.N_4466\);
    
    \I2.STOP_RDSRAM_1488\ : DFFC
      port map(CLK => CLK_c, D => \I2.STOP_RDSRAM_453_i_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.STOP_RDSRAM_595\);
    
    \I2.PIPE8_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_558_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl30r_net_1\);
    
    EF_pad : IB33
      port map(PAD => EF, Y => EF_c);
    
    \I3.PIPEA_237\ : MUX2L
      port map(A => \I3.PIPEAl6r_net_1\, B => 
        \I3.PIPEA_8l6r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854676__net_1\, Y
         => \I3.PIPEA_237_net_1\);
    
    \I3.VDBOFFB_30_IV_0L2R_2453\ : OR2
      port map(A => \I3.VDBoffb_30l2r_adt_net_162741_\, B => 
        \I3.VDBoffb_30l2r_adt_net_162742_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162747_\);
    
    \I2.OFFSETl1r_1572\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_561_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL1R_679\);
    
    \I2.SUB9_1_ADD_18x18_fast_I60_Y\ : OAI21TTF
      port map(A => \I2.SUB8l15r_adt_net_855572__net_1\, B => 
        \I2.N296_adt_net_69573_\, C => \I2.N328_adt_net_70573_\, 
        Y => \I2.N328\);
    
    \I1.PAGECNTlde_0_o2_2_1238\ : NAND2FT
      port map(A => \I1.N_310_RD1__335\, B => 
        \I1.N_311_i_i_Rd1__net_1\, Y => \I1.N_325_500\);
    
    \I2.OFFSET_37_16l4r\ : MUX2L
      port map(A => \REGl265r\, B => \REGl201r\, S => 
        \I2.PIPE7_DTL27R_80\, Y => \I2.N_759\);
    
    \I2.PIPE7_DTL27R_2796\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_89\);
    
    \I3.un6_tcnt1_i\ : INV
      port map(A => \I3.TCNT1l0r_net_1\, Y => \I3.TCNT1_i_0l0r\);
    
    \I3.REG_1_159\ : MUX2L
      port map(A => VDB_inl10r, B => REGl58r, S => 
        \I3.N_1935_adt_net_855328__net_1\, Y => \I3.REG_1_159_0\);
    
    \I2.TDCDRYBS\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDRYB_c, Q => 
        \I2.TDCDRYBS_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I43_Y\ : AND2
      port map(A => \I2.N235\, B => \I2.N238\, Y => \I2.N308\);
    
    \I3.un1_singcyc8_i_0_o3\ : OR2
      port map(A => \I3.ASBS_net_1\, B => 
        \I3.N_80_adt_net_159051_\, Y => \I3.N_80\);
    
    \I2.PIPE1_DT_42_1_ivl18r\ : OR3
      port map(A => \I2.PIPE1_DT_42l18r_adt_net_47443_\, B => 
        \I2.PIPE1_DT_42l18r_adt_net_47455_\, C => 
        \I2.PIPE1_DT_42l18r_adt_net_47456_\, Y => 
        \I2.PIPE1_DT_42l18r\);
    
    VDB_padl3r : IOB33PH
      port map(PAD => VDB(3), A => \I3.VDBml3r_net_1\, EN => 
        \I3.un1_vdb_0\, Y => VDB_inl3r);
    
    RAMDT_padl4r : IOB33PH
      port map(PAD => RAMDT(4), A => \I1.RAMDT_SPI_1l4r_net_1\, 
        EN => \I1.RAMDT_SPI_e_net_1\, Y => RAMDT_inl4r);
    
    \I2.TOKINAi\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKINAi_325_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => TOKINA_c);
    
    \I1.REG_17_sqmuxa_0_a2_0_a3_0_a2_843\ : NAND2
      port map(A => \I1.N_590_230\, B => 
        \I1.PAGECNTl9r_adt_net_854816__net_1\, Y => 
        \I1.N_260_221\);
    
    \I1.sstatel10r\ : DFFS
      port map(CLK => CLK_c, D => \I1.N_43_i_0\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.sstatel10r_net_1\);
    
    PAF_pad : IB33
      port map(PAD => PAF, Y => PAF_c);
    
    \I2.un2_evnt_word_I_45\ : XOR2
      port map(A => \I2.WOFFSETl8r\, B => \I2.DWACT_FINC_E_0l4r\, 
        Y => \I2.I_45\);
    
    \I2.RAMDT4l9r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl9r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l9r_net_1\);
    
    \I3.PIPEA_8l30r\ : OR2FT
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854484__net_1\, B => 
        \I3.N_239\, Y => \I3.PIPEA_8l30r_net_1\);
    
    \I2.L2TYPE_590\ : MUX2L
      port map(A => \I2.L2TYPE_i_0_il1r\, B => \I2.N_4451\, S => 
        \I2.N_4482_0\, Y => \I2.L2TYPE_590_net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__3091\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854732__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__861\);
    
    \I3.N_1906_i_0_0_adt_net_855636_\ : BFR
      port map(A => \I3.N_1906_i_0_0\, Y => 
        \I3.N_1906_i_0_0_adt_net_855636__net_1\);
    
    \I1.REG_74_0_IVL349R_1864\ : NOR2FT
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_24_sqmuxa_adt_net_854780__net_1\, Y => 
        \I1.REG_74l349r_adt_net_116203_\);
    
    \I2.N_4250_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_4250\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.N_4250_Rd1__net_1\);
    
    REGl230r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_131_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl230r\);
    
    \I2.RAMAD_4l13r\ : MUX2L
      port map(A => \I2.N_540\, B => 
        \I1.PAGECNTl5r_adt_net_855548__net_1\, S => LOAD_RES_1, Y
         => \I2.RAMAD_4l13r_net_1\);
    
    \I2.L2TYPE_4_IL10R_1623\ : OR2FT
      port map(A => \I2.N_4456\, B => \I2.N_4459\, Y => 
        \I2.N_4442_adt_net_67433_\);
    
    \I2.resyn_0_I2_FID_432\ : MUX2H
      port map(A => FID_cl16r, B => \I2.FID_7l16r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\, 
        Y => \I2.FID_432\);
    
    REGl197r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_98_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl197r\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854484_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854492__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854484__net_1\);
    
    \I2.N_4283_i_0_a2_m1_e_0_667\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__48\, B => 
        \I2.TEMPF_net_1\, Y => \I2.N_4283_I_0_45\);
    
    \I3.VDBOFFB_30_IV_0L0R_2479\ : AND2
      port map(A => \REGl341r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        Y => \I3.VDBoffb_30l0r_adt_net_163094_\);
    
    \I2.PIPE1_DT_42_1_IVL16R_1415\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\, B => 
        \I2.PIPE1_DT_30l16r_net_1\, C => 
        \I2.PIPE1_DT_42l16r_adt_net_47835_\, Y => 
        \I2.PIPE1_DT_42l16r_adt_net_47852_\);
    
    \I2.PIPE1_DT_42_1_IVL11R_1455\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855044__net_1\, 
        B => \I2.PIPE1_DT_12l11r_net_1\, Y => 
        \I2.PIPE1_DT_42l11r_adt_net_49689_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I147_Y\ : AO21FTF
      port map(A => \I2.N325_0\, B => 
        \I2.N411_adt_net_4092__net_1\, C => \I2.N324\, Y => 
        \I2.N411\);
    
    \I2.BNCID_VECT_tile_DOUTl5r\ : MUX2L
      port map(A => \I2.DIN_REG1l5r\, B => \I2.DOUT_TMPl5r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl5r\);
    
    \I2.UN1_CHAIN_RDY_1_SQMUXA_I_1707\ : NOR3
      port map(A => \I2.STATEe_ipl1r\, B => \I2.STATEe_ipl2r\, C
         => \I2.INT_ERRS_net_1\, Y => \I2.N_3494_adt_net_90556_\);
    
    \I2.un1_NWPIPE7_2_946\ : OAI21TTF
      port map(A => \I2.CHA_DATA8_net_1\, B => 
        \I2.CHB_DATA8_net_1\, C => 
        \I2.un1_NWPIPE7_2_adt_net_73600_\, Y => 
        \I2.UN1_NWPIPE7_2_ADT_NET_73606__324\);
    
    \I3.STATE1_NS_0_IV_0_0L7R_2121\ : NOR3
      port map(A => \I3.N_1641\, B => 
        \I3.STATE1_tr24_i_0_o2_1_i_adt_net_135386_\, C => 
        \I3.TCNT_0_sqmuxa\, Y => 
        \I3.STATE1_nsl7r_adt_net_136177_\);
    
    \I2.PIPE1_DT_42_1_IVL8R_1473\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        B => \I2.PIPE1_DT_12l8r_net_1\, Y => 
        \I2.PIPE1_DT_42l8r_adt_net_50430_\);
    
    \I2.DT_TEMPl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_791_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl30r_net_1\);
    
    \I3.TCNTl2r_1168\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT_382_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TCNTL2R_430\);
    
    DPR_padl2r : IB33
      port map(PAD => DPR(2), Y => DPR_cl2r);
    
    \I2.STATE2l5r_1245\ : DFFS
      port map(CLK => CLK_c, D => \I2.N_2796_i_0\, SET => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L5R_507\);
    
    \I2.PIPE6_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_463_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl9r_net_1\);
    
    \I2.DTESl10r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl10r, Q => 
        \I2.DTESl10r_net_1\);
    
    \I3.N_57_i_0_o2\ : OR2
      port map(A => \I3.N_1912\, B => \I3.TCNTL3R_878\, Y => 
        \I3.N_1919\);
    
    \I2.un1_reg80_i\ : AND3
      port map(A => \I2.N_3824_adt_net_90293_\, B => 
        \I2.N_3824_adt_net_90294_\, C => 
        \I2.N_3824_adt_net_90298_\, Y => 
        \I2.N_3824_adt_net_90281_\);
    
    \I2.PIPE10_DT_623\ : MUX2L
      port map(A => \I2.PIPE10_DTl18r_net_1\, B => \I2.N_3804\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_623_net_1\);
    
    \I1.REG_74_0_IVL395R_1795\ : NOR2FT
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_29_sqmuxa_adt_net_855520__net_1\, Y => 
        \I1.REG_74l395r_adt_net_110612_\);
    
    \I3.VDBi_31l29r\ : MUX2L
      port map(A => \I3.REGl162r\, B => \I3.VDBi_20l29r\, S => 
        \I3.REGMAPl17r_adt_net_854280__net_1\, Y => 
        \I3.VDBi_31l29r_net_1\);
    
    \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668_\ : BFR
      port map(A => \I2.N_4646_1_ADT_NET_1645_RD1__489\, Y => 
        \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855668__net_1\);
    
    \I3.VDBi_57_0_iv_0_0l15r\ : OR2
      port map(A => \I3.VDBi_57l15r_adt_net_139971_\, B => 
        \I3.VDBi_57l15r_adt_net_139972_\, Y => \I3.VDBi_57l15r\);
    
    REGl384r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_285_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl384r\);
    
    \I2.PIPE5_DT_6l17r\ : MUX2L
      port map(A => \I2.PIPE5_DT_6_dl17r_net_1\, B => 
        \I2.un27_pipe5_dt0l17r\, S => \I2.PIPE5_DT_6_sl19r_net_1\, 
        Y => \I2.PIPE5_DT_6l17r_net_1\);
    
    \I1.REG_3_sqmuxa_0_a2_0_818_898\ : NAND2FT
      port map(A => \I1.PAGECNTL9R_244\, B => 
        \I1.N_238_Rd1__adt_net_854888__net_1\, Y => 
        \I1.N_254_276\);
    
    \I2.PIPE1_DT_42_1_IVL15R_1435\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\, B => 
        \I2.PIPE1_DT_30l15r_net_1\, C => 
        \I2.PIPE1_DT_42l15r_adt_net_48701_\, Y => 
        \I2.PIPE1_DT_42l15r_adt_net_48717_\);
    
    \I2.BNCID_VECTROR_10_TZ_0_1421\ : AND2
      port map(A => \I2.BNCID_VECTra12_1_net_1\, B => 
        \I2.BNCID_VECTro_4\, Y => 
        \I2.BNCID_VECTror_10_tz_0_adt_net_48139_\);
    
    \I2.STATE2_NS_4_0L2R_1049\ : NOR2
      port map(A => \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__158\, B
         => \I2.N_237\, Y => \I2.STATE2_nsl2r_adt_net_24911_\);
    
    \I2.MIC_ERR_REGS_335\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl7r_net_1\, B => 
        \I2.MIC_ERR_REGSl6r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855840__net_1\, Y => 
        \I2.MIC_ERR_REGS_335_net_1\);
    
    \I3.REG_1_202\ : MUX2L
      port map(A => VDB_inl21r, B => \I3.REGl154r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855296__net_1\, Y => 
        \I3.REG_1_202_0\);
    
    \I3.VDBil5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_345_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil5r_net_1\);
    
    \I2.DTOSl22r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl22r, Q => 
        \I2.DTOSl22r_net_1\);
    
    \I2.OFFSET_37_6l0r\ : MUX2L
      port map(A => \I2.N_667\, B => \I2.N_659\, S => 
        \I2.PIPE7_DTL26R_351\, Y => \I2.N_675\);
    
    \I3.PIPEBl7r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_86_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl7r_net_1\);
    
    \I2.WPAGE_950\ : MUX2H
      port map(A => \I2.WPAGEl13r_net_1\, B => 
        \I2.WPAGE_n1_net_1\, S => 
        \I2.WPAGEe_adt_net_855056__net_1\, Y => 
        \I2.WPAGE_950_net_1\);
    
    \I2.PIPE8_DT_555\ : MUX2L
      port map(A => \I2.PIPE8_DTl27r_net_1\, B => 
        \I2.PIPE8_DT_21l27r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_555_net_1\);
    
    \I1.REG_1_212\ : MUX2H
      port map(A => \REGl311r\, B => \I1.REG_74l311r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_212_net_1\);
    
    \I2.DTO_16_1l13r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l13r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l13r_Rd1__net_1\);
    
    \I2.DTE_2_1_0l10r\ : XOR2
      port map(A => \I2.CRC32l18r_net_1\, B => 
        \I2.CRC32l6r_net_1\, Y => \I2.DTE_2_1_0l10r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I54_Y_1683\ : AND2FT
      port map(A => \I2.LSRAM_OUTl13r\, B => 
        \I2.PIPE7_DTL13R_692\, Y => \I2.N304_0_adt_net_86999_\);
    
    \I2.PIPE7_DTl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl9r_net_1\);
    
    \I2.EVNT_NUM_962\ : MUX2L
      port map(A => \I2.EVNT_NUMl1r_net_1\, B => 
        \I2.EVNT_NUM_n1_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_962_net_1\);
    
    \I2.UN5_TDCGDA1_1011\ : NOR3FTT
      port map(A => \I2.un5_tdcgda1_adt_net_21626_\, B => 
        \I2.un7_tdcgda1_3_i_i\, C => \I2.un7_tdcgda1_2_i_i\, Y
         => \I2.un5_tdcgda1_adt_net_21623_\);
    
    \I2.DTE_21_1_iv_0l8r\ : OR3
      port map(A => \I2.DTE_21_1l8r_adt_net_38739_\, B => 
        \I2.DTE_21_1l8r_adt_net_38753_\, C => 
        \I2.DTE_21_1l8r_adt_net_38754_\, Y => \I2.DTE_21_1l8r\);
    
    \I2.ENDF_1511\ : DFFC
      port map(CLK => CLK_c, D => \I2.ENDF_712_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ENDF_618\);
    
    \I2.STATE1l9r_1524\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3208_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1L9R_631\);
    
    \I5.sstate1l3r\ : DFFC
      port map(CLK => CLK_c, D => \I5.N_96\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l3r_net_1\);
    
    \I3.VADm_0_a3l1r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl1r_net_1\, Y => \I3.VADml1r\);
    
    \I2.PIPE1_DT_42_1_IVL13R_1442\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl29r_net_1\, Y => 
        \I2.PIPE1_DT_42l13r_adt_net_49191_\);
    
    \I2.PIPE10_DT_630\ : MUX2L
      port map(A => \I2.PIPE10_DTl25r_net_1\, B => 
        \I2.PIPE9_DTl25r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_630_net_1\);
    
    \I1.REG_1_214\ : MUX2H
      port map(A => \REGl313r\, B => \I1.REG_74l313r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_214_net_1\);
    
    \I3.REG3l1r_1637\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG3_126_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3L1R_744\);
    
    \I2.RAMDT4L12R_2816\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_144\);
    
    \I5.sstate1se_8_0_0_m2\ : MUX2H
      port map(A => \I5.sstate1l4r_net_1\, B => 
        \I5.sstate1l5r_net_1\, S => TICKl0r, Y => 
        \I5.sstate1_ns_el9r\);
    
    \I2.STATE2_ns_a6_0_a2l3r\ : NOR2
      port map(A => \I2.N_176_i_adt_net_855708__net_1\, B => 
        \I2.DTE_cl_0_sqmuxa_2_adt_net_904__net_1\, Y => 
        \I2.STATE2_nsl3r\);
    
    \I1.REG_74_0_ivl263r\ : AO21
      port map(A => \REGl263r\, B => 
        \I1.N_137_adt_net_854760__net_1\, C => 
        \I1.REG_74l263r_adt_net_124457_\, Y => \I1.REG_74l263r\);
    
    \I2.MAJORITY_REG_I_IL7R_1214\ : OA21
      port map(A => \I2.MIC_REG3l7r_net_1\, B => 
        \I2.MIC_REG1l7r_net_1\, C => \I2.MIC_REG2l7r_net_1\, Y
         => \REGl29r_adt_net_35602_\);
    
    \I0.CLEAR\ : OR2FT
      port map(A => REGl18r, B => \I0.CLEAR_adt_net_15818_\, Y
         => \I0.CLEAR_net_1\);
    
    ADE_padl11r : OB33PH
      port map(PAD => ADE(11), A => ADE_cl11r);
    
    \I1.REG_1_229\ : MUX2H
      port map(A => \REGl328r\, B => \I1.REG_74l328r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y => 
        \I1.REG_1_229_net_1\);
    
    \I2.PIPE8_DT_21l4r\ : MUX2L
      port map(A => \I2.LSRAM_OUTl4r\, B => \I2.N_570\, S => 
        \I2.N_4707_i_0\, Y => \I2.PIPE8_DT_21l4r_net_1\);
    
    \I2.UN1_REG80_I_1704\ : AND3
      port map(A => \I2.N_3824_adt_net_90295_\, B => 
        \I2.N_3824_adt_net_90291_\, C => 
        \I2.N_3824_adt_net_90292_\, Y => 
        \I2.N_3824_adt_net_90298_\);
    
    \I2.TRGSERVl2r_1474\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TRGSERV_2l2r\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TRGSERVL2R_581\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I180_UN1_Y_2670\ : NOR3FFT
      port map(A => \I2.N309_0\, B => 
        \I2.I180_un1_Y_adt_net_309337_\, C => 
        \I2.N495_i_adt_net_202144_\, Y => 
        \I2.I180_un1_Y_adt_net_215260_\);
    
    \I2.PIPE10_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_636_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl31r_net_1\);
    
    REGl270r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_171_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl270r\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I141_Y_0_O4_2676\ : 
        NAND2FT
      port map(A => 
        \I2.N_3_0_adt_net_1070__adt_net_855604__net_1\, B => 
        \I2.N_13_1\, Y => \I2.N522_0_adt_net_329219_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I74_Y\ : AOI21
      port map(A => \I2.N236\, B => \I2.N240_0\, C => \I2.N239\, 
        Y => \I2.N324\);
    
    \I2.SRAM_EVNT_c1_i_o2\ : AND2
      port map(A => \I2.SRAM_EVNTl0r_net_1\, B => 
        \I2.SRAM_EVNTl1r_net_1\, Y => \I2.N_3855\);
    
    \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014_\ : NAND3FFT
      port map(A => \I2.ENDF_402\, B => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_20149__183\, C => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_60\, Y => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__net_1\);
    
    DTE_padl2r : IOB33PH
      port map(PAD => DTE(2), A => \I2.DTE_1l2r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl2r);
    
    \I2.CRC32_809\ : MUX2L
      port map(A => \I2.CRC32l14r_net_1\, B => \I2.N_3931\, S => 
        \I2.N_2826_1_ADT_NET_794__331\, Y => \I2.CRC32_809_net_1\);
    
    \I3.STATE2l2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE2l3r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.STATE2l2r_net_1\);
    
    \I2.TDCl1r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TDC_651_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.TDCl1r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL20R_1393\ : OAI21FTF
      port map(A => REGl440r, B => 
        \I2.N_3234_adt_net_855648__net_1\, C => 
        \I2.PIPE1_DT_42l20r_adt_net_47061_\, Y => 
        \I2.PIPE1_DT_42l20r_adt_net_47067_\);
    
    \I1.REG_1_185\ : MUX2H
      port map(A => \REGl284r\, B => \I1.REG_74l284r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\, Y
         => \I1.REG_1_185_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I182_Y\ : XOR2FT
      port map(A => \I2.N_42_0\, B => 
        \I2.ADD_21x21_fast_I182_Y_0\, Y => 
        \I2.un27_pipe5_dt0l12r\);
    
    \I2.EVNT_NUM_c8\ : AND2
      port map(A => \I2.EVNT_NUMl8r_net_1\, B => 
        \I2.EVNT_NUM_c7_net_1\, Y => \I2.EVNT_NUM_c8_net_1\);
    
    \I2.PIPE2_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl12r_net_1\);
    
    DTE_padl23r : IOB33PH
      port map(PAD => DTE(23), A => \I2.DTE_1l23r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl23r);
    
    \I1.SBYTE_8_0_a2_i_o4l0r\ : NOR2
      port map(A => \I1.sstatel6r_net_1\, B => \I1.N_362\, Y => 
        \I1.N_371_i\);
    
    \I3.REGMAPl34r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un151_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl34r_net_1\);
    
    \I2.FIDl28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_444\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl28r);
    
    \I3.REG_1l151r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_199_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl151r\);
    
    \I2.PIPE7_DTL27R_2775\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_68\);
    
    \I2.OFFSET_37_5l3r\ : MUX2L
      port map(A => \REGl400r\, B => \REGl336r\, S => 
        \I2.PIPE7_DTL27R_81\, Y => \I2.N_670\);
    
    \I5.AIR_WDATAl15r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_62_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl15r_net_1\);
    
    \I2.FID_7_0_IVL13R_966\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl61r, C => 
        \I2.FID_7l13r_adt_net_18081_\, Y => 
        \I2.FID_7l13r_adt_net_18089_\);
    
    \I2.SRAM_EVNTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SRAM_EVNT_n3_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.SRAM_EVNTl3r_net_1\);
    
    \I1.REG_1_187\ : MUX2H
      port map(A => \REGl286r\, B => \I1.REG_74l286r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\, Y => 
        \I1.REG_1_187_net_1\);
    
    \I3.VDBm_0l2r\ : MUX2L
      port map(A => \I3.PIPEAl2r_net_1\, B => \I3.PIPEBl2r_net_1\, 
        S => \I3.BLTCYC_net_1\, Y => \I3.N_144\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I184_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_801\, B => 
        \I2.PIPE4_DTl14r_net_1\, Y => 
        \I2.ADD_21x21_fast_I184_Y_0_0\);
    
    \I3.STATE1_ipl0r_adt_net_854356_\ : BFR
      port map(A => \I3.STATE1_ipl0r_adt_net_854360__net_1\, Y
         => \I3.STATE1_ipl0r_adt_net_854356__net_1\);
    
    \I3.un10_tcnt2_i\ : NOR3FTT
      port map(A => \I3.un6_tcnt1_net_1\, B => 
        \I3.un10_tcnt2_adt_net_135290_\, C => 
        \I3.un10_tcnt2_adt_net_135291_\, Y => 
        \I3.un10_tcnt2_i_net_1\);
    
    \I2.STATE1l18r_1521\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.STATE1_ns_o2_0l0r_net_1\, SET => CLEAR_STAT_i_0, Q
         => \I2.STATE1L18R_628\);
    
    \I2.PIPE1_DT_30l20r\ : MUX2L
      port map(A => \I2.TDCDBSl20r_net_1\, B => 
        \I2.TDCDBSl18r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855084__net_1\, Y
         => \I2.PIPE1_DT_30l20r_net_1\);
    
    DTO_padl18r : IOB33PH
      port map(PAD => DTO(18), A => \I2.DTO_1l18r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl18r);
    
    \I2.OFFSET_37_26l4r\ : MUX2L
      port map(A => \REGl225r\, B => \I2.N_831\, S => 
        \I2.PIPE7_DTL26R_360\, Y => \I2.N_839\);
    
    \I2.G_EVNT_NUM_930\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl4r_net_1\, B => \I2.N_4344\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_930_net_1\);
    
    \I2.REG_1_n6\ : XOR2FT
      port map(A => \I2.N_3834_i_0\, B => \I2.REG_1_n6_0_net_1\, 
        Y => \I2.REG_1_n6_net_1\);
    
    \I2.TDCDASl31r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl31r, Q => 
        \I2.TDCDASl31r_net_1\);
    
    \I5.un1_sstate2_1_i_a2\ : OR2
      port map(A => \I5.sstate2l1r_net_1\, B => 
        \I5.sstate2l2r_net_1\, Y => \I5.N_480\);
    
    \I2.CRC32_7_0_x2l9r\ : XOR2
      port map(A => \I2.CRC32l9r_net_1\, B => 
        \I2.DT_TEMPl9r_net_1\, Y => \I2.N_57_i_0\);
    
    REGl392r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_293_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl392r\);
    
    \I1.PAGECNT_319_adt_net_854864_\ : BFR
      port map(A => \I1.PAGECNT_319_net_1\, Y => 
        \I1.PAGECNT_319_adt_net_854864__net_1\);
    
    \I2.DTO_16_1_IVL23R_1101\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854612__net_1\, 
        B => \I2.DT_TEMPl23r_net_1\, C => 
        \I2.DTO_16_1l23r_adt_net_30106_\, Y => 
        \I2.DTO_16_1l23r_adt_net_30114_\);
    
    \I2.BNCID_VECT_tile_0_DOUTl2r\ : MUX2L
      port map(A => \I2.DIN_REG1l2r\, B => \I2.DOUT_TMPl2r\, S
         => \I2.N_13\, Y => \I2.BNCID_VECTrxl10r\);
    
    \I2.CRC32_12_0_0_m2l25r\ : MUX2L
      port map(A => \I2.DT_TEMPl25r_net_1\, B => 
        \I2.DT_SRAMl25r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854192__net_1\, Y => 
        \I2.N_4349_i_i\);
    
    \I3.PIPEA1_12l7r\ : AND2
      port map(A => DPR_cl7r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854508__net_1\, Y => 
        \I3.PIPEA1_12l7r_net_1\);
    
    \I0.BNC_RESerr_1\ : AND2FT
      port map(A => \I0.BNC_RESF2_net_1\, B => 
        \I0.BNC_RESF1_net_1\, Y => \I0.BNC_RESerr_1_net_1\);
    
    \I5.DATAl12r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l12r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl129r);
    
    \I1.REG_1_226\ : MUX2H
      port map(A => \REGl325r\, B => \I1.REG_74l325r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y => 
        \I1.REG_1_226_net_1\);
    
    \I1.REG_74_0_IVL270R_1953\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, Y => 
        \I1.REG_74l270r_adt_net_123818_\);
    
    \I1.REG_74_2_4L228R_1851\ : AND2FT
      port map(A => \I1.N_299_adt_net_833868_Rd1__net_1\, B => 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__363\, Y => 
        \I1.REG_74_2_4_il228r_adt_net_115250_\);
    
    REGl348r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_249_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl348r\);
    
    \I3.VDBi_57l6r_adt_net_143327_\ : AO21
      port map(A => \I3.N_2045\, B => \I3.REGl97r\, C => 
        \I3.VDBi_57l6r_adt_net_143326__net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143327__net_1\);
    
    \I2.ROFFSET_n6_tz\ : XOR2
      port map(A => \I2.ROFFSETl6r_net_1\, B => 
        \I2.ROFFSET_c5_net_1\, Y => \I2.ROFFSET_n6_tz_i\);
    
    \I2.LSRAM_INl25r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_409_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl25r_net_1\);
    
    \I2.REG_1_n9_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855788__net_1\, B
         => REGl41r, Y => \I2.REG_1_n9_0_net_1\);
    
    \I1.REG_8_sqmuxa_0_a2_788\ : NOR2
      port map(A => \I1.N_268_Rd1__adt_net_854800__net_1\, B => 
        \I1.N_243_167\, Y => \I1.N_12233_I_166\);
    
    \I1.REG_74_12_0l188r_895\ : NAND3
      port map(A => \I1.N_347_adt_net_854788__net_1\, B => 
        \I1.REG_74_i_o2_i_0l364r_net_1\, C => \I1.N_57_9_i\, Y
         => \I1.N_65_12_273\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2698\ : 
        AND3FFT
      port map(A => \I2.N_128_0_adt_net_55238_\, B => 
        \I2.N_3_0_adt_net_1070__adt_net_855604__net_1\, C => 
        \I2.N_152_i_0_adt_net_502321_\, Y => 
        \I2.N_152_i_0_adt_net_502544_\);
    
    \I2.REG_1l37r_1459\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n5_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL37R_566);
    
    \I0.CLEARF2\ : DFFS
      port map(CLK => CLK_c, D => \I0.CLEARF1_i_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I0.CLEARF2_i\);
    
    \I5.sstate1_0l13r_1464\ : DFFS
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el0r\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SSTATE1L13R_571\);
    
    \I3.REGMAPl17r_adt_net_854300_\ : BFR
      port map(A => \I3.REGMAPl17r_net_1\, Y => 
        \I3.REGMAPl17r_adt_net_854300__net_1\);
    
    \I2.DTE_21_1_IVL11R_1297\ : OR3
      port map(A => \I2.DTO_16_1l11r_adt_net_32872_\, B => 
        \I2.DTE_21_1l11r_adt_net_38407_\, C => 
        \I2.DTE_21_1l11r_adt_net_38414_\, Y => 
        \I2.DTE_21_1l11r_adt_net_38416_\);
    
    \I2.CHAIN_RDY\ : DFFS
      port map(CLK => CLK_c, D => \I2.CHAIN_RDY_490_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.CHAIN_RDY_net_1\);
    
    \I1.REG_10_sqmuxa_adt_net_854716_\ : BFR
      port map(A => \I1.REG_10_sqmuxa\, Y => 
        \I1.REG_10_sqmuxa_adt_net_854716__net_1\);
    
    \I2.MIC_REG3l5r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_322_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l5r_net_1\);
    
    \I2.PIPE8_DT_553\ : MUX2L
      port map(A => \I2.PIPE8_DTl25r_net_1\, B => 
        \I2.PIPE8_DT_21l25r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_553_net_1\);
    
    \I2.RAMAD1_12l10r\ : MUX2L
      port map(A => \I2.TDCDASl21r_net_1\, B => 
        \I2.TDCDBSl21r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855180__net_1\, Y => 
        \I2.RAMAD1_12l10r_net_1\);
    
    \I3.TICKl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.un12_tcnt3_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.TICKl2r_net_1\);
    
    \I2.DTO_16_1_IVL23R_1099\ : AND2
      port map(A => \I2.STATE2l4r_adt_net_855676__net_1\, B => 
        \I2.DTO_9l23r\, Y => \I2.DTO_16_1l23r_adt_net_30100_\);
    
    \I2.PIPE5_DT_700\ : MUX2L
      port map(A => \I2.PIPE5_DTl24r_net_1\, B => 
        \I2.PIPE4_DTl24r_net_1\, S => \I2.NWPIPE4_576\, Y => 
        \I2.PIPE5_DT_700_net_1\);
    
    \I2.STATE3l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE3_ns_il11r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.STATE3l2r_net_1\);
    
    \I2.resyn_0_I2_BITCNT_n4_i_o3\ : AND2
      port map(A => \I2.N_4329\, B => \I2.BITCNT_i_0_il4r\, Y => 
        \I2.N_4330\);
    
    \I3.VDBi_57l2r_adt_net_145303_\ : AO21
      port map(A => \I3.N_2037\, B => \I3.N_134\, C => 
        \I3.VDBi_57l2r_adt_net_145285__net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145303__net_1\);
    
    \I2.L2TYPE_4_IL6R_1631\ : AND2
      port map(A => \I2.L2TYPEl6r_net_1\, B => 
        \I2.N_4446_adt_net_67934_\, Y => 
        \I2.N_4446_adt_net_67977_\);
    
    \I2.TDCDASl11r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl11r, Q => 
        \I2.TDCDASl11r_net_1\);
    
    \I2.PIPE4_DTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl2r_net_1\);
    
    \I2.L2TYPE_4_IL2R_1638\ : AND2
      port map(A => \I2.L2TYPEl2r_net_1\, B => 
        \I2.N_4450_adt_net_68435_\, Y => 
        \I2.N_4450_adt_net_68478_\);
    
    \I2.WPAGE_n2\ : XOR2
      port map(A => \I2.WPAGEl14r_net_1\, B => 
        \I2.WPAGE_c1_net_1\, Y => \I2.WPAGE_n2_net_1\);
    
    VAD_padl1r : IOB33PH
      port map(PAD => VAD(1), A => \I3.VADml1r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl1r);
    
    \I1.REG_1_132\ : MUX2H
      port map(A => \REGl231r\, B => \I1.REG_74l231r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855428__net_1\, Y => 
        \I1.REG_1_132_net_1\);
    
    \I3.VDBI_57_IV_0_0L6R_2236\ : AO21
      port map(A => \I3.PIPEAl6r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l6r_adt_net_143384_\, Y => 
        \I3.VDBi_57l6r_adt_net_143401_\);
    
    \I2.PIPE10_DT_17_il19r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l6r_net_1\, C => \I2.PIPE10_DT_17_i_0l19r_net_1\, 
        Y => \I2.N_3805\);
    
    \I2.PIPE7_DTl14r_1584\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl14r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL14R_691\);
    
    \I2.TRGARR_3_I_17\ : XOR2
      port map(A => \I2.DWACT_ADD_CI_0_g_array_12l0r\, B => 
        \I2.TRGARRl3r_net_1\, Y => \I2.TRGARR_3l3r\);
    
    \I3.VDBil25r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_365_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil25r_net_1\);
    
    \I2.PIPE10_DT_629\ : MUX2L
      port map(A => \I2.PIPE10_DTl24r_net_1\, B => 
        \I2.PIPE9_DTl24r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_629_net_1\);
    
    \I2.REG_1_n11_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855788__net_1\, B
         => REGl43r, Y => \I2.REG_1_n11_0_net_1\);
    
    \I2.STATE1_ns_il4r\ : NOR2
      port map(A => \I2.N_3287_i_0\, B => 
        \I2.N_3283_adt_net_855064__net_1\, Y => 
        \I2.STATE1_ns_il4r_net_1\);
    
    \I3.REG_44_IL84R_2307\ : AOI21FTT
      port map(A => REGl84r, B => \I3.N_98_0\, C => \I3.N_1663\, 
        Y => \I3.N_1630_adt_net_150503_\);
    
    \I1.REG_1_183\ : MUX2H
      port map(A => \REGl282r\, B => \I1.REG_74l282r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855444__net_1\, Y => 
        \I1.REG_1_183_net_1\);
    
    \I2.EVNT_NUM_n8\ : NOR2
      port map(A => EV_RES_c, B => \I2.EVNT_NUM_n8_tz_i\, Y => 
        \I2.EVNT_NUM_n8_net_1\);
    
    \I2.DTO_16_1_IVL15R_1142\ : AO21FTT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854616__net_1\, 
        B => \I2.DT_TEMPl15r_net_1\, C => 
        \I2.DTO_16_1l15r_adt_net_31956_\, Y => 
        \I2.DTO_16_1l15r_adt_net_31962_\);
    
    \I2.INT_ERRBS_527\ : MUX2L
      port map(A => \I2.INT_ERRBS_i_i\, B => 
        \I2.INT_ERRBF1_net_1\, S => 
        \I2.N_3876_adt_net_855252__net_1\, Y => 
        \I2.INT_ERRBS_527_net_1\);
    
    FID_padl26r : OB33PH
      port map(PAD => FID(26), A => FID_cl26r);
    
    \I2.NWPIPE1\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.NWPIPE1_726_net_1\, 
        SET => CLEAR_STAT_i_0, Q => \I2.NWPIPE1_net_1\);
    
    \I3.REGMAP_i_0_il40r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un181_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il40r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I176_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_800\, B => 
        \I2.PIPE4_DTl6r_net_1\, Y => 
        \I2.ADD_21x21_fast_I176_Y_0_0\);
    
    \I2.RAMDT4l12r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l12r_net_1\);
    
    DTE_padl1r : IOB33PH
      port map(PAD => DTE(1), A => \I2.DTE_1l1r_net_1\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl1r);
    
    \I1.REG_74_0_IV_0L359R_1848\ : AND2
      port map(A => \FBOUTl2r\, B => \I1.REG_25_sqmuxa\, Y => 
        \I1.REG_74l359r_adt_net_114955_\);
    
    \I3.VDBOFFB_55_2438\ : AND2FT
      port map(A => \I3.N_178_adt_net_1360__net_1\, B => 
        \I3.VDBoffbl3r_net_1\, Y => 
        \I3.VDBoffb_55_adt_net_162600_\);
    
    \I2.PIPE5_DT_6_dl18r\ : MUX2L
      port map(A => \I2.PIPE4_DTl18r_net_1\, B => 
        \I2.un27_pipe5_dt1l18r\, S => 
        \I2.N_4547_1_adt_net_1209__adt_net_855616__net_1\, Y => 
        \I2.PIPE5_DT_6_dl18r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L2R_2449\ : AO21
      port map(A => \REGl359r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        C => \I3.VDBoffb_30l2r_adt_net_162710_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162742_\);
    
    \I2.CRC32_12_i_0_x2l17r\ : XOR2FT
      port map(A => \I2.CRC32l17r_net_1\, B => \I2.N_224_i_i\, Y
         => \I2.N_252_i_i_0\);
    
    \I3.VDBi_57_0_ivl23r\ : AO21FTT
      port map(A => \I3.N_1905\, B => \I3.VDBi_31l23r_net_1\, C
         => \I3.VDBi_57l23r_adt_net_138951_\, Y => 
        \I3.VDBi_57l23r\);
    
    \I2.OFFSET_37_4l6r\ : MUX2L
      port map(A => \REGl371r\, B => \REGl307r\, S => 
        \I2.PIPE7_DTL27R_68\, Y => \I2.N_665\);
    
    \I1.REG_1_228\ : MUX2H
      port map(A => \REGl327r\, B => \I1.REG_74l327r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855508__net_1\, Y => 
        \I1.REG_1_228_net_1\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854584_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854584__net_1\);
    
    \I2.REG_1l34r_1766\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n2_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL34R_872);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I172_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l9r_net_1\, B => 
        \I2.PIPE4_DTl2r_net_1\, Y => 
        \I2.ADD_21x21_fast_I172_Y_0_0\);
    
    \I2.PIPE1_DT_42_1_IVL9R_1468\ : AND2
      port map(A => \I2.PIPE1_DT_42l15r_adt_net_48714_\, B => 
        \I2.BNCID_VECTrxl5r\, Y => 
        \I2.PIPE1_DT_42l9r_adt_net_50189_\);
    
    \I3.PIPEA1l31r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_329_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l31r_net_1\);
    
    \I1.REG_74_3_4l380r\ : OR3
      port map(A => \I1.REG_74_2_4_il228r_adt_net_115250_\, B => 
        \I1.REG_74_3_4_il380r_adt_net_123086_\, C => 
        \I1.REG_74_3_4_il380r_adt_net_123085_\, Y => 
        \I1.REG_74_3_4_il380r\);
    
    \I1.REG_74_0_iv_0l217r\ : AO21
      port map(A => \REGl217r\, B => \I1.N_89\, C => 
        \I1.REG_74l217r_adt_net_129034_\, Y => \I1.REG_74l217r\);
    
    REGl314r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_215_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl314r\);
    
    \I3.REG_44_i_a2_1_0_a3l83r\ : OR2FT
      port map(A => \I3.REGMAPl13r_net_1\, B => \I3.N_303\, Y => 
        \I3.REG_1_sqmuxa_3\);
    
    \I2.ADE_4l3r\ : MUX2H
      port map(A => \I2.WOFFSETl4r_adt_net_854980__net_1\, B => 
        \I2.ROFFSETl4r_net_1\, S => NOESRAME_c, Y => 
        \I2.ADE_4l3r_net_1\);
    
    \I2.CRC32_2l3r\ : XOR2
      port map(A => \I2.CRC32l3r_net_1\, B => 
        \I2.DT_SRAMl3r_net_1\, Y => \I2.CRC32_2l3r_net_1\);
    
    \I2.DTO_16_1_ivl30r\ : OA21FTF
      port map(A => \I2.N_182_ADT_NET_1007__386\, B => 
        \I2.DT_SRAMl30r_adt_net_854200__net_1\, C => 
        \I2.DTO_16_1_iv_1l30r_net_1\, Y => 
        \I2.DTO_16_1_ivl30r_net_1\);
    
    \I3.REGMAP_I_0_IL58R_3049\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un235_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL58R_803\);
    
    \I1.REG_15_sqmuxa_adt_net_855460_\ : BFR
      port map(A => \I1.REG_15_sqmuxa\, Y => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I151_Y_i_a2_2\ : AO21
      port map(A => \I2.RAMDT4L12R_829\, B => 
        \I2.PIPE4_DTL19R_634\, C => 
        \I2.N_152_i_0_adt_net_4117__net_1\, Y => 
        \I2.N_152_i_0_adt_net_55873_\);
    
    \I3.TCNT2_n4\ : XOR2
      port map(A => \I3.TCNT2_i_0_il4r_net_1\, B => \I3.TCNT2_c3\, 
        Y => \I3.TCNT2_n4_net_1\);
    
    \I2.DTO_16_1_IV_0L20R_1120\ : AO21
      port map(A => \I2.N_182_adt_net_1007__net_1\, B => 
        \I2.DT_SRAMl20r_net_1\, C => 
        \I2.DTO_16_1l20r_adt_net_30792_\, Y => 
        \I2.DTO_16_1l20r_adt_net_30793_\);
    
    \I2.PIPE10_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_605_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl0r_net_1\);
    
    \I3.VDBi_368\ : MUX2L
      port map(A => \I3.VDBil28r_net_1\, B => \I3.VDBi_57l28r\, S
         => \I3.UN1_STATE1_13_1_ADT_NET_1351__114\, Y => 
        \I3.VDBi_368_net_1\);
    
    \I2.G_EVNT_NUM_933\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl1r_net_1\, B => \I2.N_4637\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_933_net_1\);
    
    \I3.PIPEA_233\ : MUX2L
      port map(A => \I3.PIPEAl2r_net_1\, B => 
        \I3.PIPEA_8l2r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854680__net_1\, Y
         => \I3.PIPEA_233_net_1\);
    
    \I2.DTOSl17r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl17r, Q => 
        \I2.DTOSl17r_net_1\);
    
    \I2.DTO_16_1l21r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l21r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l21r_Rd1__net_1\);
    
    \I2.DTE_1_844\ : MUX2L
      port map(A => \I2.DTE_1l4r_Rd1__net_1\, B => 
        \I2.DTE_21_1l4r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836004_Rd1__net_1\, Y => 
        \I2.DTE_1l4r\);
    
    \I3.VDBI_57_IV_0L5R_2248\ : AO21
      port map(A => \I3.VDBil5r_net_1\, B => \I3.N_2048\, C => 
        \I3.VDBi_57l5r_adt_net_143861_\, Y => 
        \I3.VDBi_57l5r_adt_net_143862_\);
    
    \I2.PIPE1_DT_42_1_IVL17R_1406\ : AND2FT
      port map(A => \I2.PIPE1_DT_42_3_0L28R_342\, B => 
        \I2.EVNT_NUMl1r_net_1\, Y => 
        \I2.PIPE1_DT_42l17r_adt_net_47637_\);
    
    VAD_padl19r : OTB33PH
      port map(PAD => VAD(19), A => \I3.VADml19r\, EN => 
        NOEAD_c_i_0);
    
    \I3.REG1l0r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG1_133_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG1l0r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I211_Y\ : XOR2
      port map(A => \I2.N486_i\, B => 
        \I2.SUB_21x21_fast_I211_Y_0\, Y => \I2.SUB8_2l15r\);
    
    \I2.PIPE7_DTl2r_1595\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL2R_702\);
    
    \I2.DTO_16_1_IV_0L24R_1095\ : AO21
      port map(A => \I2.N_182_adt_net_1007__net_1\, B => 
        \I2.N_4194\, C => \I2.DTO_16_1l24r_adt_net_29868_\, Y => 
        \I2.DTO_16_1l24r_adt_net_29869_\);
    
    \I2.DT_TEMPl10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_771_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl10r_net_1\);
    
    REGl368r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_269_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl368r\);
    
    \I3.VDBOFFA_31_IV_0L5R_2529\ : AND2
      port map(A => \REGl234r\, B => \I3.REGMAPl26r_net_1\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163648_\);
    
    \I2.FIDl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.FID_419_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => FID_cl3r);
    
    \I2.CRC32_819\ : MUX2L
      port map(A => \I2.CRC32l24r_net_1\, B => \I2.N_3941\, S => 
        \I2.N_2826_1_ADT_NET_794__329\, Y => \I2.CRC32_819_net_1\);
    
    \I1.REG_1_186\ : MUX2H
      port map(A => \REGl285r\, B => \I1.REG_74l285r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\, Y => 
        \I1.REG_1_186_net_1\);
    
    \I3.un25_reg_ads_0_a2_0_a3\ : NOR3
      port map(A => \I3.WRITES_8\, B => \I3.N_578\, C => 
        \I3.N_573\, Y => \I3.un25_reg_ads_0_a2_0_a3_net_1\);
    
    \I3.VDBi_43l3r\ : MUX2L
      port map(A => REGl409r, B => \I3.VDBi_40l3r_net_1\, S => 
        \I3.REGMAPl55r_net_1\, Y => \I3.VDBi_43l3r_net_1\);
    
    \I2.L2ARR_941\ : MUX2L
      port map(A => \I2.L2ARRl3r_net_1\, B => \I2.L2ARR_n3_net_1\, 
        S => \I2.N_4482_0\, Y => \I2.L2ARR_941_net_1\);
    
    \I2.DTO_16_1_IV_0_0L6R_1191\ : AND2
      port map(A => \I2.DTO_1l6r\, B => \I2.N_196_52\, Y => 
        \I2.DTO_16_1l6r_adt_net_33912_\);
    
    \I2.NWPIPE8_1_sqmuxa_0_0\ : AND3
      port map(A => \I2.TRAIL_MIS7_i_net_1\, B => 
        \I2.NWPIPE7_688\, C => \I2.LSRAM_FL_RD7_net_1\, Y => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\);
    
    \I2.N_3876_adt_net_855252_\ : BFR
      port map(A => \I2.N_3876_adt_net_855256__net_1\, Y => 
        \I2.N_3876_adt_net_855252__net_1\);
    
    \I3.VDBI_57_0_IV_0L21R_2166\ : AO21
      port map(A => \I3.VDBil21r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l21r_adt_net_139179_\, Y => 
        \I3.VDBi_57l21r_adt_net_139189_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I14_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L5R_814\, B => 
        \I2.PIPE4_DTL14R_638\, Y => \I2.N_57\);
    
    \I3.VDBOFFB_30_IV_0L4R_2410\ : AO21
      port map(A => \REGl321r\, B => \I3.REGMAPl37r_net_1\, C => 
        \I3.VDBoffb_30l4r_adt_net_162318_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162359_\);
    
    \I3.N_1463_i_1_adt_net_855364_\ : BFR
      port map(A => \I3.N_1463_i_1\, Y => 
        \I3.N_1463_i_1_adt_net_855364__net_1\);
    
    \I3.REG_1L7R_901\ : OA21
      port map(A => \I3.REG1l7r_net_1\, B => \I3.REG2l7r_net_1\, 
        C => \I3.REG3l7r_net_1\, Y => \REGl7r_adt_net_8466_\);
    
    \I2.END_TDC2\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_TDC1_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_TDC2_net_1\);
    
    FBOUTl6r : DFFC
      port map(CLK => CLK_c, D => \I1.SBYTE_64_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \FBOUTl6r\);
    
    \I2.un1_DTO_cl_1_sqmuxa_2_0_o2\ : OR2FT
      port map(A => \I2.N_2870\, B => 
        \I2.un1_DTO_cl_1_sqmuxa_2_adt_net_22202_\, Y => 
        \I2.un1_DTO_cl_1_sqmuxa_2\);
    
    \I3.REG3l0r\ : DFFS
      port map(CLK => CLK_c, D => \I3.REG3_125_net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG3l0r_net_1\);
    
    \I1.REG_1_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_242\, B => \I1.N_255\, Y => 
        \I1.REG_1_sqmuxa\);
    
    \I1.PAGECNT_321_adt_net_854880_\ : BFR
      port map(A => \I1.PAGECNT_321_net_1\, Y => 
        \I1.PAGECNT_321_adt_net_854880__net_1\);
    
    \I1.REG_74_2l404r\ : OR3FFT
      port map(A => \I1.REG_74_2_0l404r_Rd1__net_1\, B => 
        \I1.REG_74_11_a0l404r_net_1\, C => 
        \I1.N_1169_adt_net_854828__net_1\, Y => \I1.N_273_9\);
    
    \I2.PIPE10_DT_17_il15r\ : OA21TTF
      port map(A => \I2.N_3822_adt_net_855588__net_1\, B => 
        \I2.SUB9l2r_net_1\, C => \I2.PIPE10_DT_17_i_0l15r_net_1\, 
        Y => \I2.N_3801\);
    
    \I1.REG_1_297\ : MUX2H
      port map(A => \REGl396r\, B => \I1.REG_74l396r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855528__net_1\, Y
         => \I1.REG_1_297_net_1\);
    
    \I5.SENS_ADDR_1_SQMUXA_927\ : NAND3FFT
      port map(A => \I5.SENS_ADDRl0r_net_1\, B => 
        \I5.SENS_ADDRl1r_net_1\, C => \I5.SENS_ADDRl2r_net_1\, Y
         => \I5.SENS_ADDR_1_sqmuxa_adt_net_14344_\);
    
    \I3.VDBi_57_iv_0_0l0r\ : OR3
      port map(A => \I3.VDBi_57l0r_adt_net_146655_\, B => 
        \I3.VDBi_57l0r_adt_net_146660_\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_4066__net_1\, Y
         => \I3.VDBi_57l0r\);
    
    \I2.SUB8l14r_adt_net_855568_\ : BFR
      port map(A => \I2.SUB8l14r_net_1\, Y => 
        \I2.SUB8l14r_adt_net_855568__net_1\);
    
    \I3.TCNT_n4_0_0_x2\ : XOR2
      port map(A => \I3.N_1919\, B => \I3.TCNTl4r_net_1\, Y => 
        \I3.N_263_i\);
    
    \I1.REG_1_262\ : MUX2H
      port map(A => \REGl361r\, B => \I1.REG_74l361r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_262_net_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I38_Y_1646\ : AO21
      port map(A => \I2.N_3543_i_i\, B => \I2.G_1_0\, C => 
        \I2.N_3545_i_i\, Y => \I2.N303_adt_net_69116_\);
    
    \I3.VDBi_40_1l12r\ : MUX2L
      port map(A => REGl129r, B => \I3.VDBi_31l12r_net_1\, S => 
        \I3.REGMAPl16r_net_1\, Y => \I3.N_350\);
    
    \I3.PIPEA1_317\ : MUX2L
      port map(A => \I3.PIPEA1l19r_net_1\, B => 
        \I3.PIPEA1_12l19r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__252\, Y => 
        \I3.PIPEA1_317_net_1\);
    
    \I3.un54_reg_ads_0_a2_1_a2\ : OR2
      port map(A => \I3.N_546\, B => \I3.N_551\, Y => \I3.N_573\);
    
    \I2.resyn_0_I2_FID_431\ : MUX2H
      port map(A => FID_cl15r, B => \I2.FID_7l15r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\, 
        Y => \I2.FID_431\);
    
    \I2.PIPE10_DT_605\ : MUX2L
      port map(A => \I2.PIPE10_DTl0r_net_1\, B => 
        \I2.PIPE9_DTl0r_net_1\, S => \I2.NWPIPE9_0_7\, Y => 
        \I2.PIPE10_DT_605_net_1\);
    
    \I2.PIPE9_DT_284\ : MUX2L
      port map(A => \I2.PIPE9_DTl15r_net_1\, B => 
        \I2.PIPE8_DTl15r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_284_net_1\);
    
    \I2.OFFSET_37_6l7r\ : MUX2L
      port map(A => \I2.N_674\, B => \I2.N_666\, S => 
        \I2.PIPE7_DTL26R_350\, Y => \I2.N_682\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I164_Y_2652\ : NOR3
      port map(A => \I2.N312_0_adt_net_86445_\, B => 
        \I2.N312_0_adt_net_86450_\, C => \I2.N316_i_i\, Y => 
        \I2.N495_i_adt_net_202032_\);
    
    \I2.MIC_REG2_314\ : MUX2H
      port map(A => \I2.MIC_REG2_i_0_il5r_net_1\, B => 
        \I2.MIC_REG2l6r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855768__net_1\, Y => 
        \I2.MIC_REG2_314_net_1\);
    
    \I2.OFFSET_37_16l2r\ : MUX2L
      port map(A => \REGl263r\, B => \REGl199r\, S => 
        \I2.PIPE7_DTL27R_83\, Y => \I2.N_757\);
    
    \I3.PIPEA1_12l3r\ : AND2
      port map(A => DPR_cl3r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854452__net_1\, Y => 
        \I3.PIPEA1_12l3r_net_1\);
    
    \I3.N_1935_adt_net_855316_\ : BFR
      port map(A => \I3.N_1935\, Y => 
        \I3.N_1935_adt_net_855316__net_1\);
    
    \I5.SDAin_i_m4\ : MUX2L
      port map(A => SDAB_in, B => SDAA_in, S => 
        \I5.CHAIN_SELECT_net_1\, Y => \I5.N_101\);
    
    \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854444_\ : 
        BFR
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__46\, Y => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854444__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I208_Y_0\ : XOR2
      port map(A => \I2.LSRAM_OUTl12r\, B => 
        \I2.PIPE7_DTl12r_net_1\, Y => 
        \I2.SUB_21x21_fast_I208_Y_0\);
    
    \I1.REG_74l388r\ : OR3FTT
      port map(A => \I1.REG_74_13_388_N_11\, B => 
        \I1.N_257_adt_net_111276_\, C => 
        \I1.N_257_adt_net_111279_\, Y => \I1.N_257\);
    
    \I3.BLTCYC\ : DFFC
      port map(CLK => CLK_c, D => \I3.BLTCYC_113_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.BLTCYC_net_1\);
    
    \I1.REG_1_264\ : MUX2H
      port map(A => \REGl363r\, B => \I1.REG_74l363r\, S => 
        \I1.N_50_0_ADT_NET_1409__282\, Y => \I1.REG_1_264_net_1\);
    
    \PULSE_0L0R_ADT_NET_834380_RD1__2841\ : DFFC
      port map(CLK => CLK_c, D => 
        \I3.PULSE_330_adt_net_854736__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \PULSE_0L0R_ADT_NET_834380_RD1__199\);
    
    \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__2752\ : OAI21TTF
      port map(A => \I2.N_176_i_adt_net_855708__net_1\, B => 
        \I2.DTE_CL_0_SQMUXA_2_ADT_NET_904__159\, C => 
        \I2.N_4667_1_ADT_NET_1046__32\, Y => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\);
    
    \I2.resyn_0_I2_FID_427\ : MUX2H
      port map(A => FID_cl11r, B => \I2.FID_7l11r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855824__net_1\, 
        Y => \I2.FID_427\);
    
    \I2.DTESl29r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl29r, Q => 
        \I2.DTESl29r_net_1\);
    
    \I2.N475_adt_net_460353_\ : OR3
      port map(A => \I2.N475_adt_net_87328__net_1\, B => 
        \I2.N475_adt_net_442369__net_1\, C => 
        \I2.N475_adt_net_442371__net_1\, Y => 
        \I2.N475_adt_net_460353__net_1\);
    
    \I2.PIPE3_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl7r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl7r_net_1\);
    
    \I1.SBYTE_0_sqmuxa_0_0\ : NAND2FT
      port map(A => \I1.SBYTE_0_sqmuxa_adt_net_105487_\, B => 
        \I1.N_457\, Y => \I1.SBYTE_0_sqmuxa\);
    
    \I2.ADOl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADO_3l6r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADO_cl6r);
    
    \I2.SUB8_518\ : MUX2H
      port map(A => \I2.SUB8l15r_adt_net_855572__net_1\, B => 
        \I2.SUB8_2l15r\, S => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855140__net_1\, Y => 
        \I2.SUB8_518_net_1\);
    
    \I3.REG_1l51r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_152_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl51r);
    
    \I2.PIPE10_DT_628\ : MUX2L
      port map(A => \I2.PIPE10_DTl23r_net_1\, B => 
        \I2.PIPE9_DTl23r_net_1\, S => \I2.NWPIPE9_0_net_1\, Y => 
        \I2.PIPE10_DT_628_net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2459\ : AND2
      port map(A => \REGl286r\, B => \I3.REGMAPl33r_net_1\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162896_\);
    
    \I3.REGMAPL9R_3031\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un41_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL9R_785\);
    
    \I2.MIC_REG3l1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_318_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l1r_net_1\);
    
    \I2.STATE3l4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_12254_i\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE3l4r_net_1\);
    
    \I2.DTOSl20r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl20r, Q => 
        \I2.DTOSl20r_net_1\);
    
    \I3.PIPEA_8_0l31r\ : MUX2L
      port map(A => DPR_cl31r, B => \I3.PIPEA1l31r_net_1\, S => 
        \I3.N_1463_i_1_adt_net_855356__net_1\, Y => \I3.N_240\);
    
    \I5.AIR_WDATA_57\ : MUX2H
      port map(A => \I5.sstate2l1r_net_1\, B => 
        \I5.AIR_WDATAl2r_net_1\, S => \I5.N_461\, Y => 
        \I5.AIR_WDATA_57_net_1\);
    
    \I2.resyn_0_I2_BITCNT_n3_i_o3\ : AND2
      port map(A => \I2.N_4328\, B => \I2.BITCNTl3r_net_1\, Y => 
        \I2.N_4329\);
    
    \I2.DT_TEMP_7l3r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854256__net_1\, B => 
        \I2.DT_SRAMl3r_net_1\, Y => \I2.DT_TEMP_7l3r_net_1\);
    
    \I2.OFFSET_37_9l5r\ : MUX2L
      port map(A => \REGl394r\, B => \REGl330r\, S => 
        \I2.PIPE7_DTL27R_78\, Y => \I2.N_704\);
    
    \I2.OFFSETl3r_1570\ : DFFC
      port map(CLK => CLK_c, D => \I2.OFFSET_563_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.OFFSETL3R_677\);
    
    \I3.REG_1l111r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_292_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl111r);
    
    \I2.STATE1l8r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3234_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1l8r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I174_Y\ : XOR2
      port map(A => \I2.N394_0\, B => 
        \I2.ADD_21x21_fast_I174_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l4r\);
    
    \I2.PIPE3_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl24r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl24r_net_1\);
    
    \I2.L_LUT\ : DFFC
      port map(CLK => CLK_c, D => \I2.L_LUT_498_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L_LUT_net_1\);
    
    \I1.REG_74_0_IVL228R_1999\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => \I1.N_12233_i\, Y
         => \I1.REG_74l228r_adt_net_127964_\);
    
    \I2.L2SERVl2r_1507\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_920_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL14R_614\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I0_S_0_x2\ : XOR2
      port map(A => \I2.RAMDT4l7r_net_1\, B => 
        \I2.PIPE4_DTl0r_net_1\, Y => \I2.un27_pipe5_dt1l0r\);
    
    \I3.VDBi_57_iv_0_0_a2_2l2r\ : NAND2
      port map(A => \I3.STATE1_ipl3r_adt_net_854364__net_1\, B
         => \I3.N_57_i_0_0_adt_net_854700__net_1\, Y => 
        \I3.N_2047\);
    
    \I3.PIPEA1l0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA1_298_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l0r_net_1\);
    
    \I3.VDBil30r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_370_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil30r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL20R_1392\ : NOR2FT
      port map(A => REGl424r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, Y => 
        \I2.PIPE1_DT_42l20r_adt_net_47061_\);
    
    \I3.TCNT2_i_0_il6r\ : DFFC
      port map(CLK => CLK_c, D => TCNT2_390, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT2_i_0_il6r_net_1\);
    
    \I3.STATE1_NS_1_IV_0L2R_2097\ : AO21FTT
      port map(A => \I3.N_1904\, B => 
        \I3.N_57_i_0_0_adt_net_854692__net_1\, C => 
        \I3.STATE1_ipl0r_adt_net_854356__net_1\, Y => 
        \I3.STATE1_nsl2r_adt_net_134789_\);
    
    \I3.un106_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_580\, B => \I3.N_551\, Y => 
        \I3.un106_reg_ads_0_a2_0_a3_net_1\);
    
    RAMAD_padl11r : OB33PH
      port map(PAD => RAMAD(11), A => RAMAD_cl11r);
    
    \I2.PIPE1_DT_42_1_IVL14R_1441\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855748__net_1\, B => 
        \I2.PIPE1_DT_30l14r_net_1\, C => 
        \I2.PIPE1_DT_42l14r_adt_net_48948_\, Y => 
        \I2.PIPE1_DT_42l14r_adt_net_48964_\);
    
    \I2.PIPE10_DT_624\ : MUX2L
      port map(A => \I2.PIPE10_DTl19r_net_1\, B => \I2.N_3805\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_624_net_1\);
    
    \I1.N_65_ADT_NET_1433__2847\ : OR3
      port map(A => \I1.N_65_12_272\, B => 
        \I1.N_193_adt_net_118653__net_1\, C => \I1.N_97_6\, Y => 
        \I1.N_65_ADT_NET_1433__217\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I75_Y\ : NAND2
      port map(A => \I2.N240_0\, B => \I2.N237_0\, Y => 
        \I2.N325_0\);
    
    \I2.L2SERV_n1\ : XOR2
      port map(A => \I2.RPAGEl13r\, B => \I2.RPAGEl12r\, Y => 
        \I2.L2SERV_n1_net_1\);
    
    \I1.REG_74_0_IVL400R_1789\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_30_sqmuxa_adt_net_854376__net_1\, Y => 
        \I1.REG_74l400r_adt_net_110100_\);
    
    \I2.OFFSET_37_7l4r\ : MUX2L
      port map(A => \I2.N_679\, B => \I2.N_655\, S => 
        \I2.PIPE7_DTL25R_682\, Y => \I2.N_687\);
    
    \I2.N_2868_1_adt_net_835992_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2868_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\);
    
    \I2.PIPE8_DT_548\ : MUX2L
      port map(A => \I2.PIPE8_DTl20r_net_1\, B => 
        \I2.PIPE8_DT_21l20r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_548_net_1\);
    
    REGl356r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_257_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl356r\);
    
    \I3.REG_1l414r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_221_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl414r);
    
    \I3.TCNT3_n2\ : XOR2
      port map(A => \I3.TCNT3_i_0_il2r_net_1\, B => \I3.TCNT3_c1\, 
        Y => \I3.TCNT3_n2_net_1\);
    
    \I2.SUB8l12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_515_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l12r_net_1\);
    
    BNC_RES_pad : OB33PH
      port map(PAD => BNC_RES, A => BNC_RES_c);
    
    \I2.PIPE10_DTl8r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE10_DT_613_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE10_DTl8r_net_1\);
    
    \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__3095\ : OAI21
      port map(A => \I2.REG_0l3r_adt_net_19771_Rd1__net_1\, B => 
        \I2.REG_0l3r_adt_net_19773_Rd1__net_1\, C => 
        \I2.END_EVNT10_407\, Y => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__871\);
    
    \I1.REG_74_0_IVL344R_1869\ : AND2
      port map(A => \FBOUTl3r\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l344r_adt_net_116670_\);
    
    \I1.BITCNTL0R_2745\ : DFFC
      port map(CLK => CLK_c, D => \I1.BITCNT_317_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.BITCNTL0R_18\);
    
    RMIC_pad : OB33PH
      port map(PAD => RMIC, A => RMIC_c);
    
    \I2.N_1174_i_i_a2\ : AND2FT
      port map(A => \I2.FIFO_END_EVNT_392\, B => EVREAD_387, Y
         => \I2.N_119\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I40_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl19r\, B => 
        \I2.PIPE7_DTl19r_net_1\, Y => \I2.N288_0\);
    
    \I1.REG_74_0_IVL231R_1995\ : AND2
      port map(A => \FBOUTl2r\, B => 
        \I1.REG_9_sqmuxa_adt_net_854728__net_1\, Y => 
        \I1.REG_74l231r_adt_net_127538_\);
    
    \I2.RAMAD_4l2r\ : MUX2L
      port map(A => \I2.N_529\, B => 
        \I1.BYTECNTl2r_adt_net_855020__net_1\, S => LOAD_RES, Y
         => \I2.RAMAD_4l2r_net_1\);
    
    \I5.SBYTEl2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_67_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl2r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I121_Y_i_o4\ : OAI21
      port map(A => \I2.N_29_i_0\, B => 
        \I2.ADD_21x21_fast_I121_Y_i_a3_0_i_0\, C => \I2.N_89_0\, 
        Y => \I2.N_31_0\);
    
    \I2.DT_TEMP_7l5r\ : AND2FT
      port map(A => \I2.WR_SRAM_2_adt_net_748__net_1\, B => 
        \I2.DT_SRAMl5r_net_1\, Y => \I2.DT_TEMP_7l5r_net_1\);
    
    \I2.DTO_16_1_iv_0_o2_0_i_o2l21r_773\ : OAI21FTF
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.CRC32_1_SQMUXA_0_38\, C => 
        \I2.N_182_ADT_NET_1007__155\, Y => \I2.N_197_151\);
    
    \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__3094\ : OAI21
      port map(A => \I2.REG_0l3r_adt_net_19771_Rd1__net_1\, B => 
        \I2.REG_0l3r_adt_net_19773_Rd1__net_1\, C => 
        \I2.END_EVNT10_407\, Y => 
        \I2.DTE_0_SQMUXA_I_O2_M6_I_A5_2_I_ADT_NET_2404__870\);
    
    \I1.PAGECNTL9R_2852\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_318_adt_net_854856__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL9R_246\);
    
    RAMDT_padl12r : IOB33PH
      port map(PAD => RAMDT(12), A => \I1.RAMDT_SPI_1l5r_net_1\, 
        EN => \I1.RAMDT_SPI_E_0\, Y => RAMDT_inl12r);
    
    \I2.un2_tdcgdb1_0_adt_net_830_\ : OR3FTT
      port map(A => \I2.TDCDBSl30r_net_1\, B => 
        \I2.TDCDBSL31R_503\, C => \I2.TDCDBSl29r_net_1\, Y => 
        \I2.un2_tdcgdb1_0_adt_net_830__net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I35_P0N_1284\ : OR2FT
      port map(A => \I2.LSRAM_OUTl14r_adt_net_854944__net_1\, B
         => \I2.PIPE7_DTl14r_net_1\, Y => \I2.N273_546\);
    
    \I3.TCNT_N3_0_0_2138\ : XOR2FT
      port map(A => \I3.N_1912\, B => \I3.TCNTl3r_net_1\, Y => 
        \I3.TCNT_n3_adt_net_137329_\);
    
    N_1_I3_TCNT3_c5 : AND2
      port map(A => \I3.TCNT3l5r_net_1\, B => \I3.TCNT3_c4\, Y
         => \N_1.I3.TCNT3_c5\);
    
    \I5.REG_1l444r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_27_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl444r);
    
    \I1.BYTECNT_n3_0_x2\ : XOR2FT
      port map(A => \I1.BYTECNTl3r_net_1\, B => \I1.N_323\, Y => 
        \I1.N_392_i\);
    
    DTO_padl12r : IOB33PH
      port map(PAD => DTO(12), A => \I2.DTO_1l12r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl12r);
    
    \I2.FID_7_0_IVL24R_988\ : AO21
      port map(A => \I2.STATE3l7r_net_1\, B => REGl72r, C => 
        \I2.FID_7l24r_adt_net_19115_\, Y => 
        \I2.FID_7l24r_adt_net_19123_\);
    
    \I2.ROFFSET_248\ : NAND2FT
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855704__net_1\, B => 
        \I2.ROFFSETl12r_net_1\, Y => \I2.N_1379\);
    
    \I2.MIC_REG1_304\ : MUX2H
      port map(A => \I2.MIC_REG1l3r_adt_net_834596_Rd1__net_1\, B
         => \I2.MIC_REG1l4r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_net_1\, Y => 
        \I2.MIC_REG1_304_net_1\);
    
    \I3.VDBi_29l9r_adt_net_142020_\ : AO21
      port map(A => REGl57r, B => 
        \I3.REGMAPl9r_adt_net_854320__net_1\, C => 
        \I3.VDBi_29l9r_adt_net_142014__net_1\, Y => 
        \I3.VDBi_29l9r_adt_net_142020__net_1\);
    
    NOE32W_pad : OB33PH
      port map(PAD => NOE32W, A => NOE32W_c);
    
    REGl234r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_135_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl234r\);
    
    \I3.UN1_STATE2_15_1_ADT_NET_1342__2860\ : OR2
      port map(A => \I3.STATE2_nsl0r_adt_net_136048_\, B => 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\, Y => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__254\);
    
    \I1.PAGECNT_322_adt_net_854384_\ : BFR
      port map(A => \I1.PAGECNT_322_net_1\, Y => 
        \I1.PAGECNT_322_adt_net_854384__net_1\);
    
    \I1.REG_1_200\ : MUX2H
      port map(A => \REGl299r\, B => \I1.REG_74l299r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855464__net_1\, Y => 
        \I1.REG_1_200_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I147_Y\ : XOR2
      port map(A => \I2.N463\, B => \I2.ADD_18x18_fast_I147_Y_0\, 
        Y => \I2.SUB9_1l10r\);
    
    \I2.PIPE3_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE2_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE3_DTl27r_net_1\);
    
    \I5.REG_1l446r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_29_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl446r);
    
    \I3.VDBI_20_IVL4R_2683\ : NOR3FFT
      port map(A => REGl36r, B => \I3.REGMAPL7R_460\, C => 
        \I3.N_1907_266\, Y => \I3.VDBi_20l4r_adt_net_414879_\);
    
    \I2.ADE_4l7r\ : MUX2H
      port map(A => \I2.WOFFSETl8r\, B => \I2.ROFFSETl8r_net_1\, 
        S => NOESRAME_c, Y => \I2.ADE_4l7r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL22R_1384\ : AO21
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_1_1_adt_net_855764__net_1\, B => 
        \I2.TDCDBSl22r_net_1\, C => 
        \I2.PIPE1_DT_42l22r_adt_net_46749_\, Y => 
        \I2.PIPE1_DT_42l22r_adt_net_46764_\);
    
    \I1.REG_74_0_IVL187R_2047\ : AND2
      port map(A => \FBOUTl6r\, B => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\, Y => 
        \I1.REG_74l187r_adt_net_131699_\);
    
    \I2.PIPE1_DTl17r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_744_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl17r_net_1\);
    
    \I1.N_50_0_ADT_NET_1409__2873\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__200\, B => 
        \I1.N_50_0_ADT_NET_109751__257\, Y => 
        \I1.N_50_0_ADT_NET_1409__295\);
    
    \I2.PIPE7_DTL27R_2782\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_75\);
    
    \I3.PULSE_339\ : MUX2L
      port map(A => PULSEl9r, B => \I3.PULSE_46l9r\, S => 
        \I3.N_1409_adt_net_854740__net_1\, Y => 
        \I3.PULSE_339_net_1\);
    
    \I2.NWPIPE1_726\ : MUX2L
      port map(A => \I2.un1_STATE1_39_i_0\, B => 
        \I2.NWPIPE1_net_1\, S => \I2.un1_STATE1_38\, Y => 
        \I2.NWPIPE1_726_net_1\);
    
    \I3.EVREADi_225\ : MUX2L
      port map(A => EVREAD, B => \I3.N_1860_2\, S => 
        \I3.un1_STATE2_9_net_1\, Y => \I3.EVREADi_225_net_1\);
    
    \I2.END_EVNT10_1145\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT9_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT10_407\);
    
    \I2.DT_TEMP_7l10r\ : AND2FT
      port map(A => 
        \I2.WR_SRAM_2_adt_net_748__adt_net_854252__net_1\, B => 
        \I2.DT_SRAMl10r_net_1\, Y => \I2.DT_TEMP_7l10r_net_1\);
    
    \I2.N_3876_adt_net_855256_\ : BFR
      port map(A => \I2.N_3876\, Y => 
        \I2.N_3876_adt_net_855256__net_1\);
    
    \I1.REG_74_2_i_a2_0_0l404r\ : OR2
      port map(A => \I1.PAGECNT_319_adt_net_854864__net_1\, B => 
        \I1.PAGECNT_320_adt_net_854868__net_1\, Y => 
        \I1.REG_74_12_300_N_13_Ra1_\);
    
    \I1.REG_74l180r\ : OR3
      port map(A => \I1.N_41_8\, B => 
        \I1.N_113_ADT_NET_3714__270\, C => \I1.REG_1_sqmuxa\, Y
         => \I1.N_49\);
    
    \I2.DT_TEMPl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DT_TEMP_773_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DT_TEMPl12r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I49_Y\ : AND2
      port map(A => \I2.N279\, B => \I2.N276\, Y => \I2.N299_0\);
    
    \I1.SBYTE_0_SQMUXA_0_0_1751\ : NOR3
      port map(A => \I1.N_366\, B => \I1.sstatel2r_net_1\, C => 
        \I1.N_362\, Y => \I1.SBYTE_0_sqmuxa_adt_net_105487_\);
    
    REGl393r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_294_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl393r\);
    
    VAD_padl13r : IOB33PH
      port map(PAD => VAD(13), A => \I3.VADml13r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl13r);
    
    TDCDA_padl17r : IB33
      port map(PAD => TDCDA(17), Y => TDCDA_cl17r);
    
    \I3.STATE1_IPL2R_3100\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl8r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_IPL2R_886\);
    
    \I2.PIPE5_DTl7r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_683_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl7r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L3R_2437\ : OR3
      port map(A => \I3.VDBoffb_30l3r_adt_net_162557_\, B => 
        \I3.VDBoffb_30l3r_adt_net_162553_\, C => 
        \I3.VDBoffb_30l3r_adt_net_162554_\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162560_\);
    
    \I2.DTE_21_1_iv_0_o2_0_a2_0l12r\ : AO21TTF
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855000__net_1\, 
        B => \I2.STATE2L3R_439\, C => \I2.N_223_156\, Y => 
        \I2.N_3965_0\);
    
    \I2.PIPE1_DT_42_1_IVL18R_1402\ : NOR2FT
      port map(A => REGl422r, B => 
        \I2.STATE1_ns_0l5r_adt_net_855812__net_1\, Y => 
        \I2.PIPE1_DT_42l18r_adt_net_47449_\);
    
    \I1.N_50_0_adt_net_109760_\ : AND3
      port map(A => \I1.N_304_Rd1__net_1\, B => 
        \I1.N_50_0_adt_net_109757__net_1\, C => 
        \I1.N_50_0_adt_net_109756__net_1\, Y => 
        \I1.N_50_0_adt_net_109760__net_1\);
    
    \I1.REG_1_203\ : MUX2H
      port map(A => \REGl302r\, B => \I1.REG_74l302r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_203_net_1\);
    
    \I2.RAMDT4L5R_3061\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_815\);
    
    \I3.N_354_0_adt_net_855372_\ : BFR
      port map(A => \I3.N_354_0\, Y => 
        \I3.N_354_0_adt_net_855372__net_1\);
    
    \I2.DTE_21_1_IVL14R_1280\ : AO21FTT
      port map(A => \I2.DTO_cl_0_sqmuxa_0_adt_net_855204__net_1\, 
        B => \I2.DT_TEMPl14r_net_1\, C => 
        \I2.DTE_21_1l14r_adt_net_38053_\, Y => 
        \I2.DTE_21_1l14r_adt_net_38068_\);
    
    \I1.REG_74_0_IVL284R_1935\ : NOR2FT
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_15_sqmuxa_adt_net_855460__net_1\, Y => 
        \I1.REG_74l284r_adt_net_122377_\);
    
    \I2.CRC32_12_i_0l7r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_250_i_i_0\, Y => 
        \I2.N_3924\);
    
    \I2.RAMAD1l8r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_662_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l8r_net_1\);
    
    \I2.SUB9_582\ : MUX2H
      port map(A => \I2.SUB9l14r_net_1\, B => \I2.SUB9_1l14r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_582_net_1\);
    
    \I1.N_50_0_ADT_NET_1409__2885\ : OR2
      port map(A => \PULSE_0L0R_ADT_NET_834380_RD1__200\, B => 
        \I1.N_50_0_adt_net_109751__net_1\, Y => 
        \I1.N_50_0_ADT_NET_1409__321\);
    
    REGl328r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_229_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl328r\);
    
    \I2.PIPE4_DTl2r_1252_1752\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl2r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL2R_859\);
    
    \I2.OFFSET_37_26l2r\ : MUX2L
      port map(A => \REGl223r\, B => \I2.N_829\, S => 
        \I2.PIPE7_DTl26r_net_1\, Y => \I2.N_837\);
    
    \I1.REG_74_2l340r\ : NOR3FFT
      port map(A => \I1.N_232_1\, B => \I1.REG_74_12_300_N_15\, C
         => \I1.REG_74_2_2_il340r\, Y => \I1.N_73_10\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I180_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_801\, B => 
        \I2.PIPE4_DTl10r_net_1\, Y => 
        \I2.ADD_21x21_fast_I180_Y_0_0\);
    
    \I2.CRC32_2_0_x2l9r\ : XOR2
      port map(A => \I2.CRC32l9r_net_1\, B => \I2.N_4047\, Y => 
        \I2.N_56_i_0\);
    
    \I3.VDBI_29L3R_2701\ : AO21
      port map(A => 
        \I2.REG_0l3r_adt_net_848__adt_net_854204__net_1\, B => 
        \I3.REGMAPl1r_net_1\, C => \I3.N_2031\, Y => 
        \I3.VDBi_29l3r_adt_net_510792_\);
    
    \I2.OFFSET_37_4l5r\ : MUX2L
      port map(A => \REGl370r\, B => \REGl306r\, S => 
        \I2.PIPE7_DTL27R_69\, Y => \I2.N_664\);
    
    \I5.sstate2se_2_i\ : MUX2L
      port map(A => \I5.sstate2l1r_net_1\, B => 
        \I5.sstate2l2r_net_1\, S => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\, Y => 
        \I5.sstate2se_2_i_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2603\ : AND2
      port map(A => \REGl214r\, B => \I3.REGMAP_i_0_il24r_net_1\, 
        Y => \I3.VDBoffa_31l1r_adt_net_164416_\);
    
    \I3.VDBi_52l4r\ : MUX2H
      port map(A => \I3.VDBil4r_net_1\, B => \FBOUTl4r\, S => 
        \I3.N_57_i_0_0_adt_net_854696__net_1\, Y => 
        \I3.VDBi_52l4r_net_1\);
    
    FID_padl27r : OB33PH
      port map(PAD => FID(27), A => FID_cl27r);
    
    \I2.LSRAM_IN_401\ : MUX2L
      port map(A => \I2.PIPE5_DTl17r_net_1\, B => 
        \I2.LSRAM_INl17r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_401_net_1\);
    
    \I2.N_2828_adt_net_1062__adt_net_835304_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.N_2828_adt_net_1062__net_1\, 
        CLR => CLEAR_STAT_i_0, Q => 
        \I2.N_2828_adt_net_1062__adt_net_835304_Rd1__net_1\);
    
    \I2.PIPE5_DT_6l19r\ : MUX2L
      port map(A => \I2.PIPE5_DT_6_dl19r_net_1\, B => 
        \I2.un27_pipe5_dt0l19r\, S => \I2.PIPE5_DT_6_sl19r_net_1\, 
        Y => \I2.PIPE5_DT_6l19r_net_1\);
    
    \I2.DTE_21_1_IV_0L8R_1311\ : AND2
      port map(A => \I2.DTE_1l8r\, B => 
        \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__175\, Y => 
        \I2.DTE_21_1l8r_adt_net_38739_\);
    
    REGl274r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_175_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl274r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I120_Y_0_76_tz_tz\ : AO21
      port map(A => \I2.N_52_0\, B => \I2.N357_0\, C => 
        \I2.N_2358_tz_tz_adt_net_55567_\, Y => \I2.N_2358_tz_tz\);
    
    \I2.SUB9_573\ : MUX2H
      port map(A => \I2.SUB9l5r_net_1\, B => \I2.SUB9_1l5r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_573_net_1\);
    
    \I2.REG_0l3r_adt_net_848__adt_net_854220_\ : BFR
      port map(A => 
        \I2.REG_0l3r_adt_net_848__adt_net_854228__net_1\, Y => 
        \I2.REG_0l3r_adt_net_848__adt_net_854220__net_1\);
    
    \I1.REG_29_sqmuxa_0_a2_1_a2_841\ : OR3
      port map(A => \I1.REG_74_12_300_N_15_adt_net_3731__net_1\, 
        B => \I1.N_1169_adt_net_854812__net_1\, C => 
        \I1.N_260_221\, Y => \I1.REG_29_SQMUXA_219\);
    
    \I2.N_4646_1_adt_net_1645_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => 
        \I2.N_4646_1_adt_net_1645_Ra1__net_1\, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.N_4646_1_adt_net_1645_Rd1__net_1\);
    
    \I5.REG_1_43\ : MUX2L
      port map(A => \I5.SENS_ADDRl2r_net_1\, B => REGl430r, S => 
        \I5.REG_1_sqmuxa_0_net_1\, Y => \I5.REG_1_43_net_1\);
    
    \I3.REG_1l143r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_191_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl143r\);
    
    \I2.STATE1_ns_a3_i_o3l12r_800\ : NAND2
      port map(A => \I2.STATE1L7R_632\, B => \I2.N_3883\, Y => 
        \I2.N_3889_178\);
    
    \I2.MIC_ERR_REGSl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_359_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl30r_net_1\);
    
    \I1.REG_74_i_o2_1_0_364_m4_0\ : AND2FT
      port map(A => \I1.PAGECNT_322_net_1\, B => 
        \I1.PAGECNT_321_net_1\, Y => \I1.N_238_Ra1_\);
    
    \I1.REG_74_0_IVL301R_1917\ : AND2
      port map(A => \FBOUTl0r\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l301r_adt_net_120782_\);
    
    \I2.DTE_21_1_iv_0_0l4r\ : OR3
      port map(A => \I2.DTE_21_1l4r_adt_net_39201_\, B => 
        \I2.DTE_21_1l4r_adt_net_39209_\, C => 
        \I2.DTE_21_1l4r_adt_net_39210_\, Y => \I2.DTE_21_1l4r\);
    
    \I2.DTO_16_1l12r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l12r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l12r_Rd1__net_1\);
    
    \I2.un23_nwpipe4_i_a4\ : NOR2
      port map(A => \I2.dataout_0_adt_net_855800__net_1\, B => 
        \I2.dataout_1\, Y => \I2.N_4595\);
    
    \I3.STATE1_ns_1_iv_0l2r\ : OR2
      port map(A => \I3.STATE1_nsl2r_adt_net_134784_\, B => 
        \I3.STATE1_nsl2r_adt_net_134789_\, Y => \I3.STATE1_nsl2r\);
    
    \I3.VADm_0_a3l31r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl31r_net_1\, Y => \I3.VADml31r\);
    
    \I3.VDBOFFB_30_IV_0L7R_2352\ : AND2
      port map(A => \REGl364r\, B => \I3.REGMAP_i_0_il42r_net_1\, 
        Y => \I3.VDBoffb_30l7r_adt_net_161760_\);
    
    \I1.REG_74_0_ivl239r\ : AO21
      port map(A => \REGl239r\, B => \I1.N_113\, C => 
        \I1.REG_74l239r_adt_net_126813_\, Y => \I1.REG_74l239r\);
    
    VAD_padl6r : IOB33PH
      port map(PAD => VAD(6), A => \I3.VADml6r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl6r);
    
    \I3.VDBI_57_IV_0L5R_2244\ : AND2
      port map(A => \I3.N_2034\, B => \I3.RAMDTSl5r_net_1\, Y => 
        \I3.VDBi_57l5r_adt_net_143846_\);
    
    \I3.VDBOFFA_31_IV_0L7R_2500\ : AO21
      port map(A => \REGl196r\, B => \I3.REGMAPl21r_net_1\, C => 
        \I3.VDBoffa_31l7r_adt_net_163268_\, Y => 
        \I3.VDBoffa_31l7r_adt_net_163309_\);
    
    \I2.OFFSET_37_14l0r\ : MUX2L
      port map(A => \I2.N_731\, B => \I2.N_683\, S => 
        \I2.PIPE7_DTl24r_net_1\, Y => \I2.N_739\);
    
    \I2.CRC32_797\ : MUX2L
      port map(A => \I2.CRC32l2r_net_1\, B => \I2.N_3919\, S => 
        \I2.N_2826_1_adt_net_794__net_1\, Y => 
        \I2.CRC32_797_net_1\);
    
    NPWON_c_i : INV
      port map(A => NPWON_c, Y => NPWON_c_i_0);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I4_G0N_0_o2\ : NAND2
      port map(A => \I2.RAMDT4L11R_441\, B => 
        \I2.PIPE4_DTL4R_477\, Y => \I2.N_67\);
    
    \I2.DTE_21_1_IV_0_0L17R_1225\ : AO21
      port map(A => \I2.N_3965_0\, B => \I2.G_EVNT_NUMl1r_net_1\, 
        C => \I2.DTE_21_1l17r_adt_net_36140_\, Y => 
        \I2.DTE_21_1l17r_adt_net_36154_\);
    
    \I3.VDBml10r\ : MUX2L
      port map(A => \I3.VDBil10r_net_1\, B => \I3.N_152\, S => 
        \I3.SINGCYC_881\, Y => \I3.VDBml10r_net_1\);
    
    \I2.MIC_ERR_REGS_366\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl38r_net_1\, B => 
        \I2.MIC_ERR_REGSl37r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_366_net_1\);
    
    \I3.PIPEA1_12l9r\ : AND2
      port map(A => DPR_cl9r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854504__net_1\, Y => 
        \I3.PIPEA1_12l9r_net_1\);
    
    \I2.BNCID_VECT_tile_0_DIN_REG1l1r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl9r_net_1\, Q => 
        \I2.DIN_REG1l1r\);
    
    \I2.G_EVNT_NUMl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_923_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl11r_net_1\);
    
    \I2.PIPE1_DT_30l16r\ : MUX2L
      port map(A => \I2.TDCDBSl16r_net_1\, B => 
        \I2.TDCDBSl14r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855072__net_1\, Y
         => \I2.PIPE1_DT_30l16r_net_1\);
    
    \I2.LEAD_FLAG6_638\ : AO21
      port map(A => \I2.N_4534_adt_net_1171__net_1\, B => 
        \I2.N_4534_adt_net_64476_\, C => 
        \I2.LEAD_FLAG6_638_adt_net_64516_\, Y => 
        \I2.LEAD_FLAG6_638_net_1\);
    
    \I2.PIPE4_DTL4R_3088\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL4R_852\);
    
    \I2.resyn_0_I2_TRAIL_MIS6_491\ : MUX2L
      port map(A => \I2.TRAIL_MIS6_net_1\, B => \I2.N_4643\, S
         => END_FLUSH_560, Y => \I2.TRAIL_MIS6_491\);
    
    \I2.DTO_16_1l25r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTO_16_1l25r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTO_16_1l25r_Rd1__net_1\);
    
    DTO_padl2r : IOB33PH
      port map(PAD => DTO(2), A => \I2.DTO_1l2r_net_1\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl2r);
    
    \I3.PIPEB_94\ : AO21
      port map(A => DPR_cl15r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_94_adt_net_160083_\, Y => 
        \I3.PIPEB_94_net_1\);
    
    \I1.REG_1_88\ : MUX2H
      port map(A => \REGl187r\, B => \I1.REG_74l187r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855420__net_1\, Y => 
        \I1.REG_1_88_net_1\);
    
    \I3.PIPEA_236\ : MUX2L
      port map(A => \I3.PIPEAl5r_net_1\, B => 
        \I3.PIPEA_8l5r_net_1\, S => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854676__net_1\, Y
         => \I3.PIPEA_236_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I144_Y_2657\ : AO21
      port map(A => \I2.N319_0\, B => \I2.N322\, C => \I2.N318\, 
        Y => \I2.N510_adt_net_232425_\);
    
    \I2.REG_1_C7_I_1741\ : NOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855784__net_1\, B
         => \I2.N_126\, Y => \I2.N_3836_i_0_adt_net_101388_\);
    
    \I5.sstate1se_1_i_0_m4\ : MUX2L
      port map(A => \I5.sstate1l12r_net_1\, B => 
        \I5.sstate1l11r_net_1\, S => TICKL0R_558, Y => \I5.N_100\);
    
    \I3.PIPEB_85_2338\ : NOR2FT
      port map(A => \I3.PIPEBl6r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_85_adt_net_160461_\);
    
    \I2.PIPE8_DT_554\ : MUX2L
      port map(A => \I2.PIPE8_DTl26r_net_1\, B => 
        \I2.PIPE8_DT_21l26r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_554_net_1\);
    
    \I2.PIPE9_DTl24r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_293_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl24r_net_1\);
    
    \I3.REG1_138\ : MUX2L
      port map(A => VDB_inl5r, B => \I3.REG1l5r_net_1\, S => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\, Y => 
        \I3.REG1_138_net_1\);
    
    \I3.VASl14r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_76_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VAS_i_0_il14r\);
    
    \I2.PIPE8_DT_21_0l29r\ : AO21FTT
      port map(A => \I2.N_565_0_adt_net_855732__net_1\, B => 
        \I2.PIPE8_DTl29r_net_1\, C => 
        \I2.PIPE8_DT_21l29r_adt_net_82644_\, Y => 
        \I2.PIPE8_DT_21l29r\);
    
    \I2.N_4667_1_adt_net_1046__adt_net_854424_\ : BFR
      port map(A => \I2.N_4667_1_adt_net_1046__net_1\, Y => 
        \I2.N_4667_1_adt_net_1046__adt_net_854424__net_1\);
    
    \I1.N_193_adt_net_1425_\ : OR3FFT
      port map(A => \I1.N_179\, B => \I1.N_185_9\, C => 
        \I1.N_193_adt_net_118660__net_1\, Y => 
        \I1.N_193_adt_net_1425__net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I188_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L12R_800\, B => 
        \I2.PIPE4_DTl18r_net_1\, Y => 
        \I2.ADD_21x21_fast_I188_Y_0_0\);
    
    \I3.REG_1_164\ : MUX2L
      port map(A => VDB_inl15r, B => REGl63r, S => 
        \I3.N_1935_adt_net_855324__net_1\, Y => \I3.REG_1_164_0\);
    
    \I2.PIPE4_DTl12r_1250\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl12r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL12R_512\);
    
    \I2.OFFSET_37_9l4r\ : MUX2L
      port map(A => \REGl393r\, B => \REGl329r\, S => 
        \I2.PIPE7_DTL27R_79\, Y => \I2.N_703\);
    
    \I3.VDBOFFB_30_IV_0L4R_2412\ : AO21
      port map(A => \REGl297r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l4r_adt_net_162326_\, Y => 
        \I3.VDBoffb_30l4r_adt_net_162361_\);
    
    \I2.L2TYPE_4_0_o2l15r\ : OR2
      port map(A => \I2.N_4454\, B => \I2.N_4455\, Y => 
        \I2.N_4468\);
    
    \I2.PIPE1_DT_30l30r\ : OA21
      port map(A => \I2.un2_tdcgdb1_0_adt_net_21805__net_1\, B
         => \I2.TDCDBSl28r_net_1\, C => \I2.TDCDBSl30r_net_1\, Y
         => \I2.PIPE1_DT_30l30r_net_1\);
    
    \I2.BNCID_VECTror_adt_net_48219_\ : AND2
      port map(A => \I2.BNCID_VECTra14_1_net_1\, B => 
        \I2.BNCID_VECTro_2\, Y => 
        \I2.BNCID_VECTror_adt_net_48219__net_1\);
    
    ADE_padl10r : OB33PH
      port map(PAD => ADE(10), A => ADE_cl10r);
    
    \I5.sstate1l10r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el3r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l10r_net_1\);
    
    \I2.LEAD_FLAG6_7_I_0_O2L7R_1593\ : NAND2FT
      port map(A => END_FLUSH_560, B => \I2.PIPE5_DTl31r_net_1\, 
        Y => \I2.N_222_adt_net_63455_\);
    
    \I2.L2TYPE_601\ : MUX2L
      port map(A => \I2.L2TYPEl12r_net_1\, B => \I2.N_4440\, S
         => \I2.N_4482_0\, Y => \I2.L2TYPE_601_net_1\);
    
    \I2.OFFSET_37_6l6r\ : MUX2L
      port map(A => \I2.N_673\, B => \I2.N_665\, S => 
        \I2.PIPE7_DTL26R_351\, Y => \I2.N_681\);
    
    \I1.REG_74_0_IVL324R_1892\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_20_sqmuxa_adt_net_855484__net_1\, Y => 
        \I1.REG_74l324r_adt_net_118701_\);
    
    \I2.PIPE1_DT_2_sqmuxa_1_1_799\ : NOR2FT
      port map(A => \I2.TDCGDB1_net_1\, B => \I2.N_3889_179\, Y
         => \I2.PIPE1_DT_2_SQMUXA_1_1_177\);
    
    \I3.PIPEB_97_2326\ : NOR2FT
      port map(A => \I3.PIPEBl18r_net_1\, B => 
        \I3.un1_STATE2_6_1_adt_net_1481__net_1\, Y => 
        \I3.PIPEB_97_adt_net_159957_\);
    
    \I2.STATE1l10r_1483\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3206_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1L10R_590\);
    
    \I2.un2_chain_errs_i_a2\ : NOR2FT
      port map(A => \I2.CHAIN_ERRS_net_1\, B => 
        \I2.INT_ERRS_net_1\, Y => \I2.N_3510\);
    
    \I2.RAMAD_4l11r\ : MUX2L
      port map(A => \I2.N_538\, B => 
        \I1.PAGECNTl3r_adt_net_835116_Rd1__net_1\, S => 
        LOAD_RES_1, Y => \I2.RAMAD_4l11r_net_1\);
    
    \I2.DTO_16_1_IVL22R_1110\ : AO21
      port map(A => \I2.DTO_1l22r\, B => \I2.N_196_53\, C => 
        \I2.DTO_16_1l22r_adt_net_30346_\, Y => 
        \I2.DTO_16_1l22r_adt_net_30362_\);
    
    \I1.PAGECNTL6R_2854\ : DFFC
      port map(CLK => CLK_c, D => 
        \I1.PAGECNT_321_adt_net_854880__net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.PAGECNTL6R_248\);
    
    \I5.SDAnoe_8_adt_net_991_\ : OAI21FTF
      port map(A => \I5.sstate1l7r_net_1\, B => \I5.N_67\, C => 
        \I5.N_71\, Y => \I5.SDAnoe_8_adt_net_991__net_1\);
    
    \I2.un1_tdc_res_35_i\ : AND2FT
      port map(A => \I2.N_4680_0\, B => REGl416r, Y => 
        \I2.N_4616_i_0\);
    
    \I2.N_2828_adt_net_1062_\ : OAI21FTF
      port map(A => \I2.N_4261\, B => \I2.N_2838_i_0\, C => 
        \I2.N_2828_adt_net_39957__net_1\, Y => 
        \I2.N_2828_adt_net_1062__net_1\);
    
    \I1.REG_74_0_ivl390r\ : AO21
      port map(A => \REGl390r\, B => \I1.N_265\, C => 
        \I1.REG_74l390r_adt_net_111042_\, Y => \I1.REG_74l390r\);
    
    \I3.RAMDTSl0r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl0r, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.RAMDTSl0r_net_1\);
    
    \I3.VDBi_40_0_i_m2l8r\ : MUX2L
      port map(A => REGl426r, B => REGl442r, S => 
        \I3.REGMAPl57r_net_1\, Y => \I3.N_2271\);
    
    \I3.PIPEB_90\ : AO21
      port map(A => DPR_cl11r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855284__net_1\, 
        C => \I3.PIPEB_90_adt_net_160251_\, Y => 
        \I3.PIPEB_90_net_1\);
    
    \I1.REG_74_0_IVL224R_2003\ : AND2
      port map(A => \FBOUTl3r\, B => \I1.N_12233_i\, Y => 
        \I1.REG_74l224r_adt_net_128308_\);
    
    \I3.REG_1_ml70r\ : AND2
      port map(A => REGl70r, B => 
        \I3.REGMAPl9r_adt_net_854312__net_1\, Y => 
        \I3.VDBi_20l22r\);
    
    \I3.VDBml1r\ : MUX2L
      port map(A => \I3.VDBil1r_net_1\, B => \I3.N_143\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml1r_net_1\);
    
    \I5.sstate1l2r\ : DFFC
      port map(CLK => CLK_c, D => \I5.sstate1_ns_el11r\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.sstate1l2r_net_1\);
    
    \I1.REG_1_237\ : MUX2H
      port map(A => \REGl336r\, B => \I1.REG_74l336r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855504__net_1\, Y => 
        \I1.REG_1_237_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I164_Y_2654\ : NOR2
      port map(A => \I2.N255_0\, B => \I2.N312_0_adt_net_86445_\, 
        Y => \I2.N495_i_adt_net_202144_\);
    
    \I2.DTO_9_iv_0_o2l0r\ : OAI21TTF
      port map(A => \I2.N_4283_i_0_adt_net_854972__net_1\, B => 
        \I2.DT_TEMPl0r_net_1\, C => 
        \I2.DTO_9_ivl0r_adt_net_35332_\, Y => \I2.DTO_9_ivl0r\);
    
    \I2.DTE_1l16r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1l16r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l16r_Rd1__net_1\);
    
    \I2.REG_1_c12_i\ : OAI21FTF
      port map(A => \I2.un8_evread_1_adt_net_855788__net_1\, B
         => \I2.N_136_1\, C => \I2.N_3841_i_0_adt_net_101174_\, Y
         => \I2.N_3841_i_0\);
    
    \I2.DTO_16_1_IV_0L5R_1196\ : AO21
      port map(A => \I2.N_182_ADT_NET_1007__385\, B => 
        \I2.DT_SRAMl5r_net_1\, C => 
        \I2.DTO_16_1l5r_adt_net_34198_\, Y => 
        \I2.DTO_16_1l5r_adt_net_34199_\);
    
    \I2.DTOSl28r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl28r, Q => 
        \I2.DTOSl28r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L7R_2355\ : AO21
      port map(A => \REGl404r\, B => \I3.REGMAPl47r_net_1\, C => 
        \I3.VDBoffb_30l7r_adt_net_161744_\, Y => 
        \I3.VDBoffb_30l7r_adt_net_161788_\);
    
    \I3.VDBoff_4_i_il4r\ : MUX2L
      port map(A => \I3.VDBoffbl4r_net_1\, B => 
        \I3.VDBoffal4r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_2068\);
    
    \I3.RAMAD_VME_36\ : MUX2H
      port map(A => RAMAD_VMEl12r, B => \I3.REGl95r\, S => 
        \I3.TCNT_0_sqmuxa_0\, Y => \I3.RAMAD_VME_36_net_1\);
    
    \I2.un5_tdcgda1\ : OR2
      port map(A => \I2.un5_tdcgda1_adt_net_21623_\, B => 
        \I2.FIRST_TDC_i_0_i\, Y => \I2.un5_tdcgda1_net_1\);
    
    \I5.SBYTEl4r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_69_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl4r_net_1\);
    
    ADO_padl1r : OB33PH
      port map(PAD => ADO(1), A => ADO_cl1r);
    
    \I1.REG_74_0_ivl296r\ : AO21
      port map(A => \REGl296r\, B => \I1.N_169\, C => 
        \I1.REG_74l296r_adt_net_121212_\, Y => \I1.REG_74l296r\);
    
    \I3.VDBOFFB_30_IV_0L1R_2466\ : AO21
      port map(A => \REGl294r\, B => \I3.REGMAPl34r_net_1\, C => 
        \I3.VDBoffb_30l1r_adt_net_162896_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162931_\);
    
    \I1.REG_74L388R_1803\ : AO21FTF
      port map(A => 
        \I1.REG_74_1_396_m7_i_3_adt_net_854840__net_1\, B => 
        \I1.REG_74_24_404_N_6_i_i\, C => \I1.REG_29_SQMUXA_219\, 
        Y => \I1.N_257_adt_net_111276_\);
    
    DTO_padl16r : IOB33PH
      port map(PAD => DTO(16), A => \I2.DTO_1l16r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl16r);
    
    \I5.COMMAND_4l15r\ : MUX2L
      port map(A => \I5.AIR_WDATAl15r_net_1\, B => REGl116r, S
         => REGl7r, Y => \I5.COMMAND_4l15r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I210_Y\ : XOR2
      port map(A => \I2.N489_i\, B => 
        \I2.SUB_21x21_fast_I210_Y_0\, Y => \I2.SUB8_2l14r\);
    
    \I2.PIPE8_DT_530\ : MUX2L
      port map(A => \I2.PIPE8_DTl2r_net_1\, B => 
        \I2.PIPE8_DT_21l2r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_530_net_1\);
    
    \I3.TCNT2_n1\ : XOR2
      port map(A => \I3.TCNT2_i_0_il0r_net_1\, B => 
        \I3.TCNT2l1r_net_1\, Y => \I3.TCNT2_n1_net_1\);
    
    \I2.PIPE9_DTl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_282_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl13r_net_1\);
    
    \I2.PIPE6_DT_483\ : MUX2H
      port map(A => \I2.PIPE5_DTl29r_net_1\, B => 
        \I2.PIPE6_DTl29r_net_1\, S => 
        \I2.un1_end_flush_9_1_adt_net_1193__net_1\, Y => 
        \I2.PIPE6_DT_483_net_1\);
    
    \I2.un1_TOKENB_CNT_I_10\ : XOR2
      port map(A => \I2.TOKENB_CNTl1r_net_1\, B => 
        \I2.DWACT_ADD_CI_0_TMP_1l0r\, Y => \I2.I_10\);
    
    \I2.RAMDT4L5R_3059\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl5r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L5R_813\);
    
    \I2.PIPE1_DTl11r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_738_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl11r_net_1\);
    
    \I2.PIPE9_DTl6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_275_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl6r_net_1\);
    
    \I2.BNCID_VECTwa15_1\ : AND2
      port map(A => \I2.TRGARRl0r_net_1\, B => 
        \I2.TRGARRl1r_net_1\, Y => \I2.BNCID_VECTwa15_1_net_1\);
    
    \I2.PIPE2_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl21r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl21r_net_1\);
    
    \I2.DT_SRAM_0l25r\ : MUX2L
      port map(A => \I2.PIPE10_DTl25r_net_1\, B => 
        \I2.PIPE5_DTl25r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854220__net_1\, Y => 
        \I2.N_893\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I154_Y_0_o2\ : OAI21FTT
      port map(A => \I2.N_32_0\, B => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4\, C => \I2.N_8_0\, Y
         => \I2.N_82_0\);
    
    \I2.BITCNTl2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.BITCNT_938\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.BITCNTl2r_net_1\);
    
    VAD_padl26r : OTB33PH
      port map(PAD => VAD(26), A => \I3.VADml26r\, EN => 
        NOEAD_c_i_0);
    
    \I1.REG_1_250\ : MUX2H
      port map(A => \REGl349r\, B => \I1.REG_74l349r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_250_net_1\);
    
    \I3.VDBOFFA_31_IV_0L5R_2537\ : AO21
      port map(A => \REGl186r\, B => \I3.REGMAPl20r_net_1\, C => 
        \I3.VDBoffa_31l5r_adt_net_163652_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163690_\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I40_Y_1654\ : AO21
      port map(A => \I2.N_3541_i_i\, B => \I2.G_1_1\, C => 
        \I2.N_3543_i_i\, Y => \I2.N305_adt_net_70150_\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2277\ : AND2
      port map(A => \I3.N_2036\, B => 
        \I3.VDBi_57_iv_0_0_o2_0_8_tzl0r_net_1\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146426_\);
    
    \I2.BNCID_VECT_tile_0_WADDR_REG1l0r\ : DFF
      port map(CLK => CLK_c, D => \I2.TRGARRl0r_net_1\, Q => 
        \I2.WADDR_REG1l0r\);
    
    \I2.resyn_0_I2_FID_435\ : MUX2H
      port map(A => FID_cl19r, B => \I2.FID_7l19r\, S => 
        \I2.un1_STATE3_10_1_adt_net_999__adt_net_855820__net_1\, 
        Y => \I2.FID_435\);
    
    \I1.REG_74_3_i_a2_i_0l172r\ : NAND3FFT
      port map(A => \I1.N_1169_168\, B => 
        \I1.REG_74_4_i_a2_404_N_4_i_adt_net_1465__net_1\, C => 
        \I1.REG_74_5_404_M1_E_0_279\, Y => \I1.N_273_6_i_0\);
    
    \I2.RAMAD_4_0l12r\ : MUX2H
      port map(A => \I2.RAMAD1l12r_net_1\, B => RAMAD_VMEl12r, S
         => \REG_i_il5r_adt_net_855552__net_1\, Y => \I2.N_539\);
    
    \I3.REG3_0_sqmuxa_adt_net_855632_\ : BFR
      port map(A => \I3.REG3_0_sqmuxa\, Y => 
        \I3.REG3_0_sqmuxa_adt_net_855632__net_1\);
    
    \I2.PIPE10_DT_17_I_A3_2L13R_1610\ : OR3
      port map(A => \I2.N_3822_adt_net_64757_\, B => 
        \I2.SUB9_i_0_il15r\, C => \I2.SUB9l14r_net_1\, Y => 
        \I2.N_3822_adt_net_64763_\);
    
    \I3.un161_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_554\, B => \I3.N_582\, Y => 
        \I3.un161_reg_ads_0_a2_0_a3_net_1\);
    
    \I3.REG_1l102r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_283_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl102r);
    
    \I2.STATE3_ns_a7l9r\ : AND2FT
      port map(A => \I2.N_3012\, B => 
        \I2.N_12254_i_adt_net_24491_\, Y => \I2.N_12254_i\);
    
    \I2.DTE_1_863\ : MUX2L
      port map(A => \I2.DTE_1l25r_Rd1__net_1\, B => 
        \I2.N_4644_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835992_Rd1__net_1\, Y => 
        \I2.DTE_1l25r\);
    
    \I2.SUB8l14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB8_517_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB8l14r_net_1\);
    
    \I3.REGMAPL16R_2927\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un64_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPL16R_444\);
    
    \I2.PIPE7_DTL27R_2784\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_77\);
    
    \I3.VDBOFFA_31_IV_0L5R_2544\ : OR3
      port map(A => \I3.VDBoffa_31l5r_adt_net_163695_\, B => 
        \I3.VDBoffa_31l5r_adt_net_163689_\, C => 
        \I3.VDBoffa_31l5r_adt_net_163690_\, Y => 
        \I3.VDBoffa_31l5r_adt_net_163699_\);
    
    \I0.COM_SERF1\ : DFFC
      port map(CLK => CLK_c, D => COM_SER_c, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I0.COM_SERF1_net_1\);
    
    \I3.REG_1_270\ : MUX2H
      port map(A => REGl89r, B => \I3.N_1635\, S => 
        \I3.N_127_adt_net_855312__net_1\, Y => \I3.REG_1_270_0\);
    
    \I2.DTE_21_1_IV_0L9R_1305\ : AND2
      port map(A => \I2.N_4047\, B => 
        \I2.N_199_0_ADT_NET_1054__36\, Y => 
        \I2.DTE_21_1l9r_adt_net_38625_\);
    
    \I2.majority_reg_i_il7r\ : AO21
      port map(A => \I2.MIC_REG3l7r_net_1\, B => 
        \I2.MIC_REG1l7r_net_1\, C => \REGl29r_adt_net_35602_\, Y
         => REGl29r);
    
    \I2.un28_sram_empty_15_0\ : MUX2L
      port map(A => \I2.N_633\, B => \I2.N_626\, S => 
        \I2.RPAGEL12R_608\, Y => \I2.un28_sram_empty\);
    
    \I2.CRC32_2l1r\ : XOR2FT
      port map(A => \I2.CRC32l1r_net_1\, B => 
        \I2.DT_SRAMl1r_net_1\, Y => \I2.CRC32_2_il1r\);
    
    \I2.DTE_2_1l5r\ : XOR2
      port map(A => \I2.CRC32l1r_net_1\, B => 
        \I2.DTE_2_1_0l5r_net_1\, Y => \I2.DTE_2_1l5r_net_1\);
    
    \I3.PIPEA1_301\ : MUX2L
      port map(A => \I3.PIPEA1l3r_net_1\, B => 
        \I3.PIPEA1_12l3r_net_1\, S => 
        \I3.un1_STATE2_15_1_adt_net_1342__net_1\, Y => 
        \I3.PIPEA1_301_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2613\ : AO21
      port map(A => \REGl166r\, B => \I3.REGMAPl18r_net_1\, C => 
        \I3.VDBoffa_31l1r_adt_net_164428_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164454_\);
    
    \I2.SUB8_1_sqmuxa_0_adt_net_855136_\ : BFR
      port map(A => \I2.SUB8_1_sqmuxa_0\, Y => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855136__net_1\);
    
    TDC_RESB_pad : OB33PH
      port map(PAD => TDC_RESB, A => TDC_RES_c_c);
    
    \I2.END_EVNT1\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.END_EVNT1_710_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.END_EVNT1_net_1\);
    
    \I2.un1_STATE2_15_i_0_a2_1_i_677\ : NAND2
      port map(A => \I2.STATE2L5R_508\, B => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__58\, Y => 
        \I2.N_4641_55\);
    
    \I3.VDBI_57_0_IV_0L19R_2172\ : AND2
      port map(A => \I3.PIPEAl19r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l19r_adt_net_139387_\);
    
    \I1.REG_1_253\ : MUX2H
      port map(A => \REGl352r\, B => \I1.REG_74l352r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_253_net_1\);
    
    \I2.ADEl4r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l4r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl4r);
    
    \I3.VDBOFFA_31_IV_0L1R_2605\ : AND2
      port map(A => \REGl270r\, B => \I3.REGMAPl31r_net_1\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164424_\);
    
    \I3.REG_1l159r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_207_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl159r\);
    
    \I2.STATE2l4r_adt_net_855688_\ : BFR
      port map(A => \I2.STATE2l4r_net_1\, Y => 
        \I2.STATE2l4r_adt_net_855688__net_1\);
    
    \I3.REG2l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG2_146_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REG2l5r_net_1\);
    
    \I3.PIPEAl27r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEA_258_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl27r_net_1\);
    
    \I2.REG_1_n0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => \I2.REG_1_n0_0_net_1\, Y => \I2.REG_1_n0_net_1\);
    
    \I2.I_1338_G_1\ : XOR2FT
      port map(A => \I2.SUB8L6R_706\, B => \I2.OFFSETL3R_677\, Y
         => \I2.G_1_3\);
    
    \I2.SUB8l11r_adt_net_855580_\ : BFR
      port map(A => \I2.SUB8l11r_net_1\, Y => 
        \I2.SUB8l11r_adt_net_855580__net_1\);
    
    \I2.L2TYPE_599\ : MUX2L
      port map(A => \I2.L2TYPEl10r_net_1\, B => \I2.N_4442\, S
         => \I2.N_4482_0\, Y => \I2.L2TYPE_599_net_1\);
    
    \I2.PIPE7_DTl8r_1590\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl8r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL8R_697\);
    
    \I2.OFFSET_37_24l0r\ : MUX2L
      port map(A => \I2.N_811\, B => \I2.N_803\, S => 
        \I2.PIPE7_DTL26R_356\, Y => \I2.N_819\);
    
    \I2.BNCID_VECTria_7_0\ : AND2
      port map(A => \I2.BNCID_VECTra15_1_net_1\, B => 
        \I2.BNCID_VECTro_7\, Y => \I2.BNCID_VECTria_7_0_net_1\);
    
    \I2.PIPE9_DT_273\ : MUX2L
      port map(A => \I2.PIPE9_DTl4r_net_1\, B => 
        \I2.PIPE8_DTl4r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_6\, Y
         => \I2.PIPE9_DT_273_net_1\);
    
    VAD_padl17r : OTB33PH
      port map(PAD => VAD(17), A => \I3.VADml17r\, EN => 
        NOEAD_c_i_0);
    
    \I2.DTE_1_855\ : MUX2L
      port map(A => \I2.DTE_1l15r_Rd1__net_1\, B => 
        \I2.DTE_21_1l15r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_835996_Rd1__net_1\, Y => 
        \I2.DTE_1l15r\);
    
    \I5.SBYTE_9_1L0R_922\ : AND2
      port map(A => \I5.sstate1l5r_net_1\, B => \I5.N_101\, Y => 
        \I5.SBYTE_9l0r_adt_net_11050_\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I153_Y_i_a4_0_1\ : OA21
      port map(A => \I2.PIPE4_DTL11R_408\, B => 
        \I2.PIPE4_DTL12R_510\, C => \I2.RAMDT4L12R_823\, Y => 
        \I2.N_112_1\);
    
    \I2.N_2864_0_adt_net_835284_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.N_2864_0_adt_net_854268__net_1\, CLR => 
        CLEAR_STAT_i_0, Q => 
        \I2.N_2864_0_adt_net_835284_Rd1__net_1\);
    
    \I2.DT_SRAMl0r_998\ : MUX2L
      port map(A => \I2.N_868\, B => \I2.PIPE2_DTl0r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAML0R_376\);
    
    \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_28083_\ : OAI21FTF
      port map(A => \I2.NWPIPE2_net_1\, B => 
        \I2.DTO_16_1_iv_0_o2_2tt_21_m3_net_1\, C => 
        \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_1085__net_1\, Y
         => \I2.DTO_16_1_iv_0_a2_5_0_0l21r_adt_net_28083__net_1\);
    
    \I1.PAGECNT_n6_i_i_o2_1\ : NOR2FT
      port map(A => \I1.PAGECNT_324_net_1\, B => \I1.N_305_Ra1_\, 
        Y => \I1.N_308_Ra1_\);
    
    \I3.VDBI_57_0_IV_0_0L8R_2223\ : AND2FT
      port map(A => \I3.N_1905_1_adt_net_855384__net_1\, B => 
        \I3.VDBi_57l8r_adt_net_1606__net_1\, Y => 
        \I3.VDBi_57l8r_adt_net_142784_\);
    
    \I2.STATE1l17r_1467\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_3798\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1L17R_574\);
    
    \I2.RAMAD_4l15r\ : MUX2L
      port map(A => \I2.N_542\, B => \I1.PAGECNTl7r_net_1\, S => 
        LOAD_RES_1, Y => \I2.RAMAD_4l15r_net_1\);
    
    \I2.RAMAD1l0r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.RAMAD1_654_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.RAMAD1l0r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2462\ : AND2
      port map(A => \REGl342r\, B => \I3.REGMAP_i_0_il40r_net_1\, 
        Y => \I3.VDBoffb_30l1r_adt_net_162908_\);
    
    \I2.UN1_PIPE1_DT_1_SQMUXA_2_0_A3_998\ : AND2
      port map(A => \I2.STATE1L7R_633\, B => \I2.N_3879\, Y => 
        \I2.N_3902_adt_net_20437_\);
    
    \I3.REG_1_188\ : MUX2L
      port map(A => VDB_inl7r, B => \I3.REGl140r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855304__net_1\, Y => 
        \I3.REG_1_188_0\);
    
    \I1.REG_74_i_o2_1_0_364_m1\ : NAND2FT
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854400__net_1\, 
        B => \I1.REG_74_i_o2_1_0tt_364_m2_e_net_1\, Y => 
        \I1.REG_74_i_o2_1_0_364_N_2\);
    
    TDCDA_padl9r : IB33
      port map(PAD => TDCDA(9), Y => TDCDA_cl9r);
    
    \I2.PIPE4_DTL9R_3036\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTL9R_790\);
    
    \I1.N_50_0_adt_net_109751_\ : NOR3FFT
      port map(A => \I1.N_232_1_296\, B => 
        \I1.N_50_0_adt_net_109760__net_1\, C => \I1.N_435_1\, Y
         => \I1.N_50_0_adt_net_109751__net_1\);
    
    \I2.L2TYPEl2r_1546\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2TYPE_591_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2TYPEL2R_653\);
    
    \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_1085_\ : AO21FTT
      port map(A => \I2.N_4030\, B => 
        \I2.DTO_16_1_iv_0_o2_2tt_21_m3_net_1\, C => 
        \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_28030__net_1\, Y
         => \I2.DTO_16_1_iv_0_o2_2_21_b0_0_1_adt_net_1085__net_1\);
    
    \I2.DTE_1l31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_1_869_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_1l31r_net_1\);
    
    \I5.AIR_WDATAl11r\ : DFFC
      port map(CLK => CLK_c, D => \I5.AIR_WDATA_61_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.AIR_WDATAl11r_net_1\);
    
    \I1.REG_3_sqmuxa_adt_net_855408_\ : BFR
      port map(A => \I1.REG_3_sqmuxa\, Y => 
        \I1.REG_3_sqmuxa_adt_net_855408__net_1\);
    
    \I1.ISI_0_SQMUXA_1_0_I_2075\ : AO21
      port map(A => \I1.N_366\, B => \I1.N_463_1\, C => 
        \PULSE_0l0r_adt_net_834380_Rd1__adt_net_854908__net_1\, Y
         => \I1.N_1375_adt_net_134070_\);
    
    REGl194r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_95_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl194r\);
    
    \I2.OFFSET_37_1l0r\ : MUX2L
      port map(A => \REGl349r\, B => \REGl285r\, S => 
        \I2.PIPE7_DTL27R_66\, Y => \I2.N_635\);
    
    FID_padl3r : OB33PH
      port map(PAD => FID(3), A => FID_cl3r);
    
    \I2.W_ERR_WORDS\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.W_ERR_WORDS_327_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.W_ERR_WORDS_net_1\);
    
    \I3.REG_1_I_IL18R_934\ : OA21
      port map(A => \I3.REG3l405r_net_1\, B => 
        \I3.REG2l405r_net_1\, C => \I3.REG1l405r_net_1\, Y => 
        \REGl18r_adt_net_15773_\);
    
    \I1.N_1367_i_adt_net_854516_\ : BFR
      port map(A => \I1.N_1367_i\, Y => 
        \I1.N_1367_i_adt_net_854516__net_1\);
    
    \I2.CRC32_12_il0r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_4027_i_0\, Y => 
        \I2.N_3917\);
    
    \I2.FID_7_0_IVL7R_1718\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl7r_net_1\, 
        Y => \I2.FID_7l7r_adt_net_92833_\);
    
    \I3.VDBI_57_0_IVL26R_2151\ : AND2
      port map(A => \I3.PIPEAl26r_net_1\, B => \I3.N_90_i_0_1\, Y
         => \I3.VDBi_57l26r_adt_net_138571_\);
    
    \I3.REG_1l161r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_209_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.REGl161r\);
    
    \I3.un1_noe64ri\ : OR2FT
      port map(A => \I3.MBLTCYC_844\, B => \I3.ADACKCYC_727\, Y
         => NOEAD_c);
    
    \I2.UN1_STATE1_39_6_1527\ : NAND2FT
      port map(A => \I2.N_3277\, B => \I2.PIPE1_DT_42_1l29r\, Y
         => \I2.un1_STATE1_39_6_i_adt_net_52470_\);
    
    \I1.REG_74_0_iv_0l221r\ : AO21
      port map(A => \FBOUTl0r\, B => \I1.N_12233_i\, C => 
        \I1.REG_74l221r_adt_net_128566_\, Y => \I1.REG_74l221r\);
    
    \I3.VAS_67\ : MUX2L
      port map(A => VAD_inl5r, B => \I3.VASl5r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_67_net_1\);
    
    \I2.N_4283_i_0_a2_m1_e_0_665\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__47\, B => 
        \I2.TEMPF_adt_net_855740__net_1\, Y => \I2.N_4283_I_0_43\);
    
    \I2.STATE2L3R_2923\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl2r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L3R_440\);
    
    \I2.L2TYPE_4_i_o2_0l13r\ : NAND2FT
      port map(A => \I2.L2ARRl1r_net_1\, B => \I2.L2ARRl0r_net_1\, 
        Y => \I2.N_4457\);
    
    \I3.PULSE_46_0_iv_0_0_o2l5r\ : NAND2FT
      port map(A => \I3.STATE1_ipl3r_adt_net_854368__net_1\, B
         => \I3.N_291\, Y => \I3.N_311\);
    
    \I5.SBYTEl3r\ : DFFC
      port map(CLK => CLK_c, D => \I5.SBYTE_68_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I5.SBYTEl3r_net_1\);
    
    \I3.VASl6r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VAS_68_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VASl6r_net_1\);
    
    \I2.MIC_ERR_REGSl14r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_343_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl14r_net_1\);
    
    \I2.BNCID_VECTrff_4_261_0_a2_0\ : NOR3FFT
      port map(A => TDCTRG_c, B => \I2.TRGARRl2r_net_1\, C => 
        \I2.TRGARRl3r_net_1\, Y => 
        \I2.BNCID_VECTrff_7_258_0_a2_0\);
    
    \I2.STATE2L4R_2869\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl1r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2L4R_291\);
    
    \I1.REG_74_0_IV_0L179R_2055\ : AND2
      port map(A => \REGl179r\, B => \I1.N_49_267\, Y => 
        \I1.REG_74l179r_adt_net_132424_\);
    
    \I2.PIPE8_DT_541\ : MUX2L
      port map(A => \I2.PIPE8_DTl13r_net_1\, B => 
        \I2.PIPE8_DT_21l13r_net_1\, S => 
        \I2.NWPIPE8_1_sqmuxa_0_0_net_1\, Y => 
        \I2.PIPE8_DT_541_net_1\);
    
    \I3.REGMAPl8r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un37_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPl8r_net_1\);
    
    \I2.SUB9_1_ADD_18X18_FAST_I31_Y_1650\ : NOR2
      port map(A => \I2.SUB8l14r_net_1\, B => \I2.SUB8l13r_net_1\, 
        Y => \I2.N296_adt_net_69573_\);
    
    FID_padl7r : OB33PH
      port map(PAD => FID(7), A => FID_cl7r);
    
    \I2.PIPE9_DTl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_281_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl12r_net_1\);
    
    \I2.OFFSET_37_3l1r\ : MUX2L
      port map(A => \I2.N_644\, B => \I2.N_636\, S => 
        \I2.PIPE7_DTL26R_350\, Y => \I2.N_652\);
    
    \I2.DTO_16_1_iv_1l30r\ : AO21FTT
      port map(A => \I2.DTO_1l30r_net_1\, B => \I2.N_196_53\, C
         => \I2.DTO_16_1_iv_1l30r_adt_net_28472_\, Y => 
        \I2.DTO_16_1_iv_1l30r_net_1\);
    
    \I2.un7_bnc_id_1_I_23\ : AND2
      port map(A => \I2.N_37\, B => \I2.BNC_IDL4R_712\, Y => 
        \I2.N_34_0\);
    
    \I2.PIPE8_DTl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE8_DT_531_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE8_DTl3r_net_1\);
    
    \I1.REG_74_12_0l188r\ : NAND3
      port map(A => \I1.N_347_adt_net_854788__net_1\, B => 
        \I1.REG_74_i_o2_i_0l364r_net_1\, C => \I1.N_57_9_i\, Y
         => \I1.N_65_12\);
    
    \I2.CRC32_1_sqmuxa_1_i_o2_926\ : OR2
      port map(A => \I2.STATE2L4R_291\, B => \I2.STATE2L3R_438\, 
        Y => \I2.N_4261_304\);
    
    \I2.G_EVNT_NUM_928\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl6r_net_1\, B => \I2.N_4638\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_928_net_1\);
    
    \I2.ADD_18x18_fast_I110_Y_0_adt_net_3684_\ : OR3
      port map(A => \I2.N_3558_i_adt_net_855584__net_1\, B => 
        \I2.SUB8l13r_adt_net_855564__net_1\, C => 
        \I2.N291_adt_net_4302__net_1\, Y => 
        \I2.ADD_18x18_fast_I110_Y_0_adt_net_3684__net_1\);
    
    \I2.N411_adt_net_194981_\ : OR2FT
      port map(A => \I2.LSRAM_OUTl1r\, B => \I2.PIPE7_DTL1R_703\, 
        Y => \I2.N411_adt_net_194981__net_1\);
    
    \I2.DTE_21_1l13r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l13r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l13r_Rd1__net_1\);
    
    \I1.REG_74_0_ivl167r\ : AO21
      port map(A => \REGl167r\, B => \I1.N_41\, C => 
        \I1.REG_74l167r_adt_net_133493_\, Y => \I1.REG_74l167r\);
    
    \I2.PIPE1_DT_30l5r\ : MUX2L
      port map(A => \I2.TDCDBSl5r_net_1\, B => 
        \I2.TDCDBSl3r_net_1\, S => 
        \I2.un2_tdcgdb1_0_adt_net_830__adt_net_855080__net_1\, Y
         => \I2.PIPE1_DT_30l5r_net_1\);
    
    \I1.REG_74_0_ivl316r\ : AO21
      port map(A => \REGl316r\, B => \I1.N_185\, C => 
        \I1.REG_74l316r_adt_net_119389_\, Y => 
        \I1.REG_74l316r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I209_Y\ : XOR2
      port map(A => \I2.N492_i\, B => 
        \I2.SUB_21x21_fast_I209_Y_0\, Y => \I2.SUB8_2l13r\);
    
    \I1.REG_74_0_iv_0l191r\ : AO21
      port map(A => \FBOUTl2r\, B => \I1.REG_4_sqmuxa\, C => 
        \I1.REG_74l191r_adt_net_131355_\, Y => \I1.REG_74l191r\);
    
    \I2.STATE1_ns_i_a3l8r\ : OR2
      port map(A => \I2.STATE1l10r_net_1\, B => \I2.N_3275\, Y
         => \I2.N_3316\);
    
    \I1.RAMDT_SPI_e\ : DFFC
      port map(CLK => CLK_c, D => \I1.LOAD_RES_i_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.RAMDT_SPI_e_net_1\);
    
    \I2.MIC_ERR_REGSl36r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_365_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl36r_net_1\);
    
    \I2.NLD\ : DFFS
      port map(CLK => CLK_c, D => \I2.NLD_647_net_1\, SET => 
        CLEAR_STAT_i_0, Q => NLD_c);
    
    \I1.REG_74_2_0_i_0l188r\ : NAND3FFT
      port map(A => \I1.N_1169_168\, B => \I1.N_237\, C => 
        \I1.REG_74_5_404_M1_E_0_280\, Y => \I1.N_273_5_i\);
    
    \I3.STATE1_tr24_59_1_i_a2_0_a2_0_a2_1_a2\ : AND3FFT
      port map(A => \I3.REGMAPL18R_778\, B => 
        \I3.REGMAP_I_0_IL24R_777\, C => \I3.N_68_adt_net_134367_\, 
        Y => \I3.N_68\);
    
    \I3.VDBi_20_ivl11r\ : AO21
      port map(A => \I3.VDBi_20l12r_adt_net_140770_\, B => 
        \I3.N_278\, C => \I3.VDBi_20l11r_adt_net_141166_\, Y => 
        \I3.VDBi_20l11r\);
    
    \I2.ERR_WORDS_RDY_415\ : AO21FTT
      port map(A => \I2.ERR_WORDS_RDY_0_sqmuxa\, B => 
        \I2.ERR_WORDS_RDY_net_1\, C => 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1\, Y => 
        \I2.ERR_WORDS_RDY_415_net_1\);
    
    \I2.ROFFSETl3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_915_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl3r_net_1\);
    
    \I2.FIFO_END_EVNT_1130\ : DFFC
      port map(CLK => CLK_c, D => \I2.FIFO_END_EVNT_489_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.FIFO_END_EVNT_392\);
    
    \I3.VDBOFFA_31_IV_0L0R_2628\ : AO21
      port map(A => \REGl173r\, B => \I3.REGMAP_i_0_il19r_net_1\, 
        C => \I3.VDBoffa_31l0r_adt_net_164606_\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164641_\);
    
    \I3.VDBi_40l11r\ : MUX2L
      port map(A => \I3.N_349\, B => \I3.N_1856\, S => 
        \I3.N_354_0_adt_net_855368__net_1\, Y => 
        \I3.VDBi_40l11r_net_1\);
    
    \I2.RAMAD_4l7r\ : MUX2L
      port map(A => \I2.N_534\, B => \I1.BYTECNTl7r_net_1\, S => 
        LOAD_RES, Y => \I2.RAMAD_4l7r_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL20R_1390\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855040__net_1\, 
        B => \I2.PIPE1_DT_12l20r_net_1\, Y => 
        \I2.PIPE1_DT_42l20r_adt_net_47053_\);
    
    \I2.DTO_16_1_iv_0l24r\ : OR2
      port map(A => \I2.DTO_16_1l24r_adt_net_29869_\, B => 
        \I2.DTO_16_1l24r_adt_net_29870_\, Y => \I2.DTO_16_1l24r\);
    
    \I4.bcntl1r\ : DFFC
      port map(CLK => CLK_c, D => \I4.bcnt_6_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I4.bcntl1r_net_1\);
    
    \I2.OFFSET_37_5l7r\ : MUX2L
      port map(A => \REGl404r\, B => \REGl340r\, S => 
        \I2.PIPE7_DTL27R_74\, Y => \I2.N_674\);
    
    \I2.STATE5_ns_0l3r\ : AO21FTF
      port map(A => \I2.MSERCLKS_net_1\, B => 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1\, C => \I2.N_4332\, Y => 
        \I2.STATE5_nsl3r\);
    
    \I2.PIPE1_DT_745\ : MUX2L
      port map(A => \I2.PIPE1_DTl18r_net_1\, B => 
        \I2.PIPE1_DT_42l18r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854572__net_1\, 
        Y => \I2.PIPE1_DT_745_net_1\);
    
    REGl397r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_298_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl397r\);
    
    \I2.PIPE10_DT_17_I_A3_2L13R_1613\ : OR2FT
      port map(A => \I2.N_22_i_0\, B => 
        \I2.N_3822_adt_net_64763_\, Y => 
        \I2.N_3822_adt_net_64766_\);
    
    \I3.VDBi_57l2r_adt_net_145225_\ : AO21
      port map(A => REGl34r, B => \I3.REGMAPL7R_460\, C => 
        \I3.REGMAPl8r_net_1\, Y => 
        \I3.VDBi_57l2r_adt_net_145225__net_1\);
    
    \I3.VDBI_57_0_IVL28R_2146\ : AO21
      port map(A => \I3.VDBil28r_net_1\, B => 
        \I3.N_1910_0_adt_net_854340__net_1\, C => 
        \I3.VDBi_57l28r_adt_net_138305_\, Y => 
        \I3.VDBi_57l28r_adt_net_138311_\);
    
    \I2.PIPE5_DT_697\ : MUX2H
      port map(A => \I2.PIPE4_DTl21r_net_1\, B => 
        \I2.PIPE5_DTl21r_net_1\, S => \I2.NWPIPE4_net_1\, Y => 
        \I2.PIPE5_DT_697_net_1\);
    
    \I3.REGMAP_I_0_IL58R_2990\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un235_reg_ads_0_a2_2_a3_net_1\, Q => 
        \I3.REGMAP_I_0_IL58R_537\);
    
    \I5.SENS_ADDRl1r\ : DFFC
      port map(CLK => CLK_c, D => \I5.I_13\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I5.SENS_ADDRl1r_net_1\);
    
    \I2.un1_STATE2_7_0\ : OR3
      port map(A => \I2.STATE2l0r_net_1\, B => 
        \I2.STATE2l1r_adt_net_855124__net_1\, C => 
        \I2.un1_STATE2_7_adt_net_53240_\, Y => \I2.un1_STATE2_7\);
    
    \I2.NWPIPE6\ : DFFS
      port map(CLK => CLK_c, D => \I2.NWPIPE6_449_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I2.NWPIPE6_net_1\);
    
    \I1.REG_74_0_IV_I_A2L201R_2033\ : AND2
      port map(A => \REGl201r\, B => \I1.N_182_i\, Y => 
        \I1.N_1340_adt_net_130447_\);
    
    \I2.BNCID_VECTrff_5\ : DFFC
      port map(CLK => CLK_c, D => 
        \I2.BNCID_VECTrff_5_260_0_net_1\, CLR => CLEAR_STAT_i_0, 
        Q => \I2.BNCID_VECTro_5\);
    
    \I2.L2SERVl1r_1503\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2SERV_921_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RPAGEL13R_610\);
    
    \I2.DTE_1_849\ : MUX2L
      port map(A => \I2.DTE_1l9r_Rd1__net_1\, B => 
        \I2.DTE_21_1l9r_Rd1__net_1\, S => 
        \I2.N_2868_1_adt_net_836000_Rd1__net_1\, Y => 
        \I2.DTE_1l9r\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I205_Y\ : XOR2FT
      port map(A => \I2.N504\, B => \I2.SUB_21x21_fast_I205_Y_0\, 
        Y => \I2.SUB8_2l9r\);
    
    \I2.PIPE1_DT_42_1_IVL14R_1439\ : AO21
      port map(A => \I2.STATE1l0r_net_1\, B => 
        \I2.MIC_ERR_REGSl46r_net_1\, C => 
        \I2.PIPE1_DT_42l14r_adt_net_48944_\, Y => 
        \I2.PIPE1_DT_42l14r_adt_net_48962_\);
    
    \I5.DATA_12_IVL1R_926\ : OA21TTF
      port map(A => \I5.sstate1se_12_i_adt_net_8689_\, B => 
        REGl118r, C => \I5.SDAin_m_1_net_1\, Y => 
        \I5.DATA_12_ivl1r_adt_net_14302_\);
    
    \I2.PIPE5_DTl30r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_706_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl30r_net_1\);
    
    \I3.UN1_STATE2_15_1_ADT_NET_1342__2858\ : OR2
      port map(A => \I3.STATE2_nsl0r_adt_net_136048_\, B => 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\, Y => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__252\);
    
    \I2.DT_SRAMl6r\ : MUX2L
      port map(A => \I2.N_874\, B => \I2.PIPE2_DTl6r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__net_1\, Y => 
        \I2.DT_SRAMl6r_net_1\);
    
    \I2.CRC32_795\ : MUX2L
      port map(A => \I2.CRC32l0r_net_1\, B => \I2.N_3917\, S => 
        \I2.N_2826_1_adt_net_794__net_1\, Y => 
        \I2.CRC32_795_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I140_Y_0_o2_1_754\ : 
        OR3FFT
      port map(A => \I2.N_107\, B => \I2.N_128_134\, C => 
        \I2.N_74_i_0_i_adt_net_54331_\, Y => \I2.N_74_I_0_I_132\);
    
    \I1.REG_74_0_IVL386R_1807\ : AND2
      port map(A => \FBOUTl5r\, B => \I1.REG_28_sqmuxa\, Y => 
        \I1.REG_74l386r_adt_net_111491_\);
    
    \I3.PIPEB_86\ : AO21
      port map(A => DPR_cl7r, B => 
        \I3.un1_STATE2_7_1_adt_net_1473__adt_net_855288__net_1\, 
        C => \I3.PIPEB_86_adt_net_160419_\, Y => 
        \I3.PIPEB_86_net_1\);
    
    \I1.REG_74_0_IVL326R_1890\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_21_sqmuxa_adt_net_855496__net_1\, Y => 
        \I1.REG_74l326r_adt_net_118432_\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2523\ : AO21
      port map(A => \REGl171r\, B => \I3.REGMAPl18r_net_1\, C => 
        \I3.N_2070_adt_net_163478_\, Y => 
        \I3.N_2070_adt_net_163504_\);
    
    \I2.OFFSET_37_2l5r\ : MUX2L
      port map(A => \REGl386r\, B => \REGl322r\, S => 
        \I2.PIPE7_DTL27R_69\, Y => \I2.N_648\);
    
    \I2.L2ARR_n2\ : XOR2FT
      port map(A => \I2.L2ARRl2r_net_1\, B => \I2.N_4454\, Y => 
        \I2.L2ARR_n2_net_1\);
    
    \I2.PHASE_861\ : DFFC
      port map(CLK => CLK_c, D => \I2.NOESRAME_c_i_0\, CLR => 
        CLEAR_STAT_i_0, Q => NOESRAME_C_239);
    
    \I3.TCNT_380\ : MUX2H
      port map(A => \I3.TCNTl4r_net_1\, B => \I3.TCNT_n4\, S => 
        \I3.TCNTe\, Y => \I3.TCNT_380_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL3R_1506\ : AO21FTT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        B => \I2.PIPE1_DT_12l3r_net_1\, C => 
        \I2.PIPE1_DT_42l3r_adt_net_51627_\, Y => 
        \I2.PIPE1_DT_42l3r_adt_net_51636_\);
    
    \I2.OFFSET_566\ : MUX2L
      port map(A => \I2.OFFSETl6r_net_1\, B => \I2.OFFSET_37l6r\, 
        S => \I2.UN1_NWPIPE7_2_297\, Y => \I2.OFFSET_566_net_1\);
    
    \I1.REG_74_8_1_tzl340r\ : AND2
      port map(A => \I1.PAGECNTL5R_311\, B => 
        \I1.PAGECNT_0L7R_ADT_NET_835112_RD1__362\, Y => 
        \I1.REG_74_8_1_tzl340r_net_1\);
    
    \I2.MIC_ERR_REGSl18r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_347_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl18r_net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I48_Y\ : OR2
      port map(A => \I2.N346_adt_net_69448__net_1\, B => 
        \I2.N311_adt_net_69399_\, Y => \I2.N313_0\);
    
    \I2.OFFSET_37_5l4r\ : MUX2L
      port map(A => \REGl401r\, B => \REGl337r\, S => 
        \I2.PIPE7_DTL27R_79\, Y => \I2.N_671\);
    
    \I1.REG_20_sqmuxa_0_a2\ : NOR2
      port map(A => \I1.N_253\, B => \I1.N_243\, Y => 
        \I1.REG_20_sqmuxa\);
    
    \I3.REGMAPl12r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un51_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl12r_net_1\);
    
    \I2.RAMAD_4l10r\ : MUX2L
      port map(A => \I2.N_537\, B => 
        \I1.PAGECNTl2r_adt_net_834908_Rd1__net_1\, S => 
        LOAD_RES_1, Y => \I2.RAMAD_4l10r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I171_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l8r_net_1\, B => 
        \I2.PIPE4_DT_i_il1r_net_1\, Y => 
        \I2.ADD_21x21_fast_I171_Y_0_0\);
    
    \I5.DATAl8r\ : DFFC
      port map(CLK => CLK_c, D => \I5.DATA_12l8r_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl125r);
    
    \I3.N_1409_adt_net_854740_\ : BFR
      port map(A => \I3.N_1409_adt_net_854744__net_1\, Y => 
        \I3.N_1409_adt_net_854740__net_1\);
    
    \I3.PULSE_335\ : AO21
      port map(A => PULSEL5R_16, B => 
        \I3.N_1409_adt_net_854744__net_1\, C => \I3.PULSE_46l5r\, 
        Y => \I3.PULSE_335_net_1\);
    
    \I2.FCNT_c1_0_o3\ : OR2
      port map(A => \I2.FCNTL1R_504\, B => \I2.FCNT_C0_398\, Y
         => \I2.FCNT_c1\);
    
    \I3.PULSEl5r_638\ : DFFC
      port map(CLK => CLK_c, D => \I3.PULSE_335_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => PULSEL5R_16);
    
    \I2.L2ARRl3r_1498\ : DFFC
      port map(CLK => CLK_c, D => \I2.L2ARR_941_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.L2ARRL3R_605\);
    
    \I3.VDBm_0l12r\ : MUX2L
      port map(A => \I3.PIPEAl12r_net_1\, B => 
        \I3.PIPEBl12r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_154\);
    
    \I1.REG_1_202\ : MUX2H
      port map(A => \REGl301r\, B => \I1.REG_74l301r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_202_net_1\);
    
    \I3.VDBOFFA_31_IV_0L1R_2615\ : OR2
      port map(A => \I3.VDBoffa_31l1r_adt_net_164451_\, B => 
        \I3.VDBoffa_31l1r_adt_net_164452_\, Y => 
        \I3.VDBoffa_31l1r_adt_net_164457_\);
    
    \I2.DTO_1_893\ : MUX2L
      port map(A => \I2.DTO_1l19r_Rd1__net_1\, B => 
        \I2.DTO_16_1l19r_Rd1__net_1\, S => 
        \I2.DTE_0_sqmuxa_i_0_N_3_1_adt_net_834764_Rd1__net_1\, Y
         => \I2.DTO_1l19r\);
    
    \I2.un1_STATE1_40_1_adt_net_45389_\ : AOI21TTF
      port map(A => \I2.N_3882\, B => 
        \I2.N_3283_adt_net_855064__net_1\, C => 
        \I2.STATE1l18r_net_1\, Y => 
        \I2.un1_STATE1_40_1_adt_net_45389__net_1\);
    
    \I3.un33_reg_ads_0_a2_0_a3\ : NOR2
      port map(A => \I3.N_634\, B => \I3.N_637\, Y => 
        \I3.un33_reg_ads_0_a2_0_a3_net_1\);
    
    \I2.LSRAM_INl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.LSRAM_IN_385_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.LSRAM_INl1r_net_1\);
    
    \I5.SBYTE_71\ : MUX2H
      port map(A => \I5.SBYTEl6r_net_1\, B => \I5.N_26\, S => 
        \I5.N_406\, Y => \I5.SBYTE_71_net_1\);
    
    \I2.PIPE4_DTl22r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl22r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl22r_net_1\);
    
    \I2.PIPE1_DTl15r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_742_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl15r_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \I2.ROFFSETl1r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ROFFSET_917_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.ROFFSETl1r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I50_Y_1686\ : AND2FT
      port map(A => \I2.LSRAM_OUTl14r\, B => 
        \I2.PIPE7_DTL14R_691\, Y => \I2.N300_0_adt_net_87051_\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I18_G0N_0_a2\ : AND2
      port map(A => \I2.RAMDT4l5r_net_1\, B => 
        \I2.PIPE4_DTl18r_net_1\, Y => \I2.N313\);
    
    \I2.UN1_ERR_WORDS_RDY_0_SQMUXA_0_0_A5_1033\ : AND3FFT
      port map(A => \I2.BITCNTl2r_net_1\, B => 
        \I2.BITCNTl3r_net_1\, C => 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23152_\, Y => 
        \I2.ERR_WORDS_RDY_0_sqmuxa_1_adt_net_23155_\);
    
    \I2.N_4646_1_ADT_NET_19635__2836\ : NOR2
      port map(A => \I2.MIC_REG1L3R_ADT_NET_834596_RD1__381\, B
         => \I2.MIC_REG2L3R_ADT_NET_834020_RD1__453\, Y => 
        \I2.N_4646_1_ADT_NET_19635__185\);
    
    \I1.SSTATE_NS_0_IV_0_0L2R_1770\ : AND3FTT
      port map(A => \PULSE_0l0r_adt_net_834380_Rd1__net_1\, B => 
        \I1.N_321_adt_net_855540__net_1\, C => 
        \I1.sstatel8r_net_1\, Y => 
        \I1.sstate_nsl2r_adt_net_107620_\);
    
    \I2.LEADSRAM.M3\ : RAM256x9SST
      generic map(MEMORYFILE => "LEAD_SRAM_M3.mem")

      port map(DO8 => OPEN, DO7 => OPEN, DO6 => OPEN, DO5 => OPEN, 
        DO4 => OPEN, DO3 => OPEN, DO2 => OPEN, DO1 => 
        \I2.LSRAM_OUTl28r\, DO0 => \I2.LSRAM_OUTl27r\, WPE => 
        OPEN, RPE => OPEN, DOS => OPEN, WADDR7 => \GND\, WADDR6
         => \GND\, WADDR5 => \GND\, WADDR4 => \GND\, WADDR3 => 
        \GND\, WADDR2 => \I2.LSRAM_WADDRl2r_net_1\, WADDR1 => 
        \I2.LSRAM_WADDRl1r_net_1\, WADDR0 => 
        \I2.LSRAM_WADDRl0r_net_1\, RADDR7 => \GND\, RADDR6 => 
        \GND\, RADDR5 => \GND\, RADDR4 => \GND\, RADDR3 => \GND\, 
        RADDR2 => \I2.LSRAM_RADDRl2r_net_1\, RADDR1 => 
        \I2.LSRAM_RADDRl1r_net_1\, RADDR0 => 
        \I2.LSRAM_RADDRl0r_net_1\, DI8 => \GND\, DI7 => \GND\, 
        DI6 => \GND\, DI5 => \GND\, DI4 => 
        \I2.LSRAM_INl31r_net_1\, DI3 => \GND\, DI2 => 
        \I2.LSRAM_INl29r_net_1\, DI1 => \I2.LSRAM_INl28r_net_1\, 
        DI0 => \I2.LSRAM_INl27r_net_1\, WRB => 
        \I2.LSRAM_WR_net_1\, RDB => \I2.LSRAM_RD_net_1\, WBLKB
         => \GND\, RBLKB => \GND\, PARODD => \GND\, WCLKS => 
        CLK_c, RCLKS => CLK_c, DIS => \GND\);
    
    REGl171r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_72_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl171r\);
    
    \I2.DTESl25r\ : DFF
      port map(CLK => CLK_c, D => DTE_inl25r, Q => 
        \I2.DTESl25r_net_1\);
    
    \I1.REG_74_0_ivl287r\ : AO21
      port map(A => \REGl287r\, B => \I1.N_161\, C => 
        \I1.REG_74l287r_adt_net_122119_\, Y => \I1.REG_74l287r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I185_Y\ : XOR2FT
      port map(A => \I2.ADD_21x21_fast_I136_Y_0_o2_m4\, B => 
        \I2.ADD_21x21_fast_I185_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l15r\);
    
    \I1.REG_1_204\ : MUX2H
      port map(A => \REGl303r\, B => \I1.REG_74l303r\, S => 
        \I1.N_50_0_ADT_NET_1409__295\, Y => \I1.REG_1_204_net_1\);
    
    TDCDB_padl24r : IB33
      port map(PAD => TDCDB(24), Y => TDCDB_cl24r);
    
    \I3.UN1_STATE2_15_1_ADT_NET_1342__2857\ : OR2
      port map(A => \I3.STATE2_nsl0r_adt_net_136048_\, B => 
        \I3.un1_STATE2_15_1_adt_net_3723__net_1\, Y => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__251\);
    
    \I2.PIPE1_DT_42_1_ivl10r\ : OR3
      port map(A => \I2.PIPE1_DT_42l10r_adt_net_49942_\, B => 
        \I2.PIPE1_DT_42l10r_adt_net_49951_\, C => 
        \I2.PIPE1_DT_42l10r_adt_net_49952_\, Y => 
        \I2.PIPE1_DT_42l10r\);
    
    \I3.REG_44_i_o2l83r\ : NAND2
      port map(A => \I3.REGMAPl13r_net_1\, B => 
        \I3.STATE1_IPL8R_10\, Y => \I3.N_98\);
    
    \I2.un3_l2as_i_a2_0\ : AOI21
      port map(A => \I2.L2RF3_i\, B => \I2.L2RF2_net_1\, C => 
        \I2.L2AS_net_1\, Y => \I2.N_4482_0\);
    
    \I3.REG_1l5r\ : MUX2L
      port map(A => \I3.REG2l5r_net_1\, B => \I3.REG3l5r_net_1\, 
        S => \I3.un102_reg\, Y => REG_i_il5r);
    
    \I2.SUB8_2_0_0_SUB_21X21_FAST_I179_Y_2684\ : AND2FT
      port map(A => \I2.N303_0\, B => \I2.N350_864\, Y => 
        \I2.N481_adt_net_423940_\);
    
    \I2.DTO_16_1_iv_0_o2l8r\ : AO21FTT
      port map(A => \I2.N_4283_i_0_adt_net_854968__net_1\, B => 
        \I2.DT_TEMPl8r_net_1\, C => \I2.N_3967_adt_net_33418_\, Y
         => \I2.N_3967\);
    
    \I2.G_EVNT_NUM_931\ : MUX2L
      port map(A => \I2.G_EVNT_NUMl3r_net_1\, B => \I2.N_4343\, S
         => \I2.N_3769\, Y => \I2.G_EVNT_NUM_931_net_1\);
    
    \I2.un1_tdc_res_38_i\ : NOR2
      port map(A => \I2.N_4680_0\, B => REGl414r, Y => 
        \I2.N_4619_i_0\);
    
    \I1.REG_74_0_IV_I_A2L209R_2025\ : AND2
      port map(A => \REGl209r\, B => \I1.N_183_i_0\, Y => 
        \I1.N_1348_adt_net_129759_\);
    
    \I2.PIPE7_DTL27R_2785\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_78\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I175_Y\ : XOR2FT
      port map(A => \I2.N537_i\, B => 
        \I2.ADD_21x21_fast_I175_Y_0\, Y => \I2.un27_pipe5_dt0l5r\);
    
    \I2.OFFSET_37_3l0r\ : MUX2L
      port map(A => \I2.N_643\, B => \I2.N_635\, S => 
        \I2.PIPE7_DTL26R_350\, Y => \I2.N_651\);
    
    \I2.CRC32_12_0_0_x2l2r\ : XOR2FT
      port map(A => \I2.CRC32l2r_net_1\, B => \I2.N_4187_i_i\, Y
         => \I2.N_73_i_0_i_0\);
    
    \I2.BNCID_VECTra13_1\ : NOR2FT
      port map(A => \I2.TRGSERVL0R_465\, B => \I2.TRGSERVL1R_468\, 
        Y => \I2.BNCID_VECTra13_1_net_1\);
    
    \I1.REG_74_0_ivl399r\ : AO21
      port map(A => \REGl399r\, B => \I1.N_273\, C => 
        \I1.REG_74l399r_adt_net_110186_\, Y => \I1.REG_74l399r\);
    
    \I2.FCNTl1r\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_946_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.FCNTl1r_net_1\);
    
    \I2.DTO_16_1_IV_0L8R_1178\ : AND2FT
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        B => \I2.DT_TEMPl8r_net_1\, Y => 
        \I2.DTO_16_1l8r_adt_net_33478_\);
    
    \I3.REG_1_197\ : MUX2L
      port map(A => VDB_inl16r, B => \I3.REGl149r\, S => 
        \I3.REG_0_sqmuxa_2_adt_net_855300__net_1\, Y => 
        \I3.REG_1_197_0\);
    
    \I2.REG_1_n5\ : XOR2FT
      port map(A => \I2.N_3833_i_0\, B => \I2.REG_1_n5_0_net_1\, 
        Y => \I2.REG_1_n5_net_1\);
    
    REGl400r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_301_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl400r\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I136_Y_0_o2_m4\ : AND2
      port map(A => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_adt_net_56806_\, B => 
        \I2.N502_i_0_adt_net_490398_\, Y => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4\);
    
    \I2.MIC_REG3l2r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_319_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l2r_net_1\);
    
    COM_SER_pad : IB33
      port map(PAD => COM_SER, Y => COM_SER_c);
    
    \I2.PIPE4_DTl3r_adt_net_854548_\ : BFR
      port map(A => \I2.PIPE4_DTl3r_net_1\, Y => 
        \I2.PIPE4_DTl3r_adt_net_854548__net_1\);
    
    \I2.ADO_3l11r\ : MUX2H
      port map(A => \I2.ROFFSETl12r_net_1\, B => \I2.WOFFSETl12r\, 
        S => NOESRAME_c, Y => \I2.ADO_3l11r_net_1\);
    
    \I2.BNCID_VECTrff_9_256_0\ : AO21
      port map(A => \I2.BNCID_VECTwa13_1_net_1\, B => 
        \I2.BNCID_VECTrff_8_257_0_a2_0\, C => \I2.BNCID_VECTro_9\, 
        Y => \I2.BNCID_VECTrff_9_256_0_net_1\);
    
    \I2.CRC32_12_il23r\ : NOR2
      port map(A => \I2.N_2867_1\, B => \I2.N_129_i_0_i_0\, Y => 
        \I2.N_3940\);
    
    \I3.REGMAPL18R_3024\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un71_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPL18R_778\);
    
    \I2.N507_adt_net_347769_\ : AND3
      port map(A => \I2.N_128_135\, B => \I2.N_57\, C => 
        \I2.N_114_adt_net_275711_\, Y => 
        \I2.N507_adt_net_347769__net_1\);
    
    \I3.REGMAP_i_0_il38r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un171_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il38r_net_1\);
    
    \I1.REG_74_0_IV_0L264R_1959\ : AND2
      port map(A => \REGl264r\, B => 
        \I1.N_137_adt_net_854764__net_1\, Y => 
        \I1.REG_74l264r_adt_net_124371_\);
    
    \I3.REGMAPl47r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un216_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPl47r_net_1\);
    
    \I2.ADE_4l1r\ : MUX2H
      port map(A => \I2.WOFFSETl2r_adt_net_854984__net_1\, B => 
        \I2.ROFFSETl2r_net_1\, S => NOESRAME_c, Y => 
        \I2.ADE_4l1r_net_1\);
    
    \I1.REG_74_0_IVL195R_2039\ : AND2
      port map(A => \FBOUTl6r\, B => \I1.REG_4_sqmuxa\, Y => 
        \I1.REG_74l195r_adt_net_131011_\);
    
    \I3.REG_1_175\ : MUX2L
      port map(A => VDB_inl26r, B => REGl74r, S => 
        \I3.N_1935_adt_net_855316__net_1\, Y => \I3.REG_1_175_0\);
    
    \I3.REGMAPl7r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un33_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl7r_net_1\);
    
    \I2.MIC_REG1_301\ : MUX2L
      port map(A => \I2.MIC_REG1l1r_net_1\, B => 
        \I2.MIC_REG1l0r_net_1\, S => 
        \I2.MIC_REG1_0_sqmuxa_0_adt_net_855776__net_1\, Y => 
        \I2.MIC_REG1_301_net_1\);
    
    \I2.PIPE1_DT_1_sqmuxa_0_a3\ : AND3FFT
      port map(A => \I2.CHAINA_EN244_i_adt_net_855260__net_1\, B
         => \I2.N_3881\, C => \I2.STATE1L12R_646\, Y => 
        \I2.PIPE1_DT_1_sqmuxa\);
    
    \I3.un1_STATE1_13_1_adt_net_137902_\ : AO21FTT
      port map(A => \I3.N_277\, B => \I3.STATE1_ipl9r\, C => 
        \I3.STATE1_nsl3r_adt_net_136439_\, Y => 
        \I3.un1_STATE1_13_1_adt_net_137902__net_1\);
    
    \I3.un106_reg_ads_0_a2_0_a2_0_988\ : NOR2FT
      port map(A => \I3.VASl12r_net_1\, B => \I3.N_547_370\, Y
         => \I3.N_548_366\);
    
    \I2.EVNT_NUM_960\ : MUX2L
      port map(A => \I2.EVNT_NUMl3r_net_1\, B => 
        \I2.EVNT_NUM_n3_net_1\, S => \I2.N_3770\, Y => 
        \I2.EVNT_NUM_960_net_1\);
    
    \I2.PIPE9_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_288_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl19r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2595\ : AO21
      port map(A => \REGl271r\, B => \I3.REGMAPl31r_net_1\, C => 
        \I3.VDBoffa_31l2r_adt_net_164238_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164264_\);
    
    \I2.TDCDASl6r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl6r, Q => 
        \I2.TDCDASl6r_net_1\);
    
    \I2.CRC32l10r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_805_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l10r_net_1\);
    
    \I2.FID_7_0_ivl24r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl24r_net_1\, 
        C => \I2.FID_7l24r_adt_net_19123_\, Y => \I2.FID_7l24r\);
    
    \I3.un91_reg_ads_0_a2_0_a2\ : OR3
      port map(A => \I3.VASl4r_net_1\, B => \I3.VASl1r_net_1\, C
         => \I3.N_549_365\, Y => \I3.N_583\);
    
    \I5.COMMAND_4l8r\ : MUX2L
      port map(A => \I5.AIR_WDATAl8r_net_1\, B => REGl109r, S => 
        REGl7r, Y => \I5.COMMAND_4l8r_net_1\);
    
    \I2.G_EVNT_NUM_n6_i_a2\ : NOR2
      port map(A => \I2.N_4672\, B => \I2.G_EVNT_NUMl6r_net_1\, Y
         => \I2.N_280\);
    
    \I2.FID_7_0_IVL26R_983\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl26r_net_1\, 
        Y => \I2.FID_7l26r_adt_net_18927_\);
    
    \I3.TCNT2_n3\ : XOR2
      port map(A => \I3.TCNT2l3r_net_1\, B => \I3.TCNT2_c2\, Y
         => \I3.TCNT2_n3_net_1\);
    
    \I2.STATE2_NS_I_0_O2_0_0_M7_I_1003\ : OR2
      port map(A => \I2.ENDF_401\, B => \I2.TEMPF_393\, Y => 
        \I2.N_4273_adt_net_20927_\);
    
    \I2.PIPE7_DTL27R_2778\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTL27R_71\);
    
    \I1.REG_22_sqmuxa_adt_net_855492_\ : BFR
      port map(A => \I1.REG_22_sqmuxa\, Y => 
        \I1.REG_22_sqmuxa_adt_net_855492__net_1\);
    
    \I3.EFS\ : DFFS
      port map(CLK => CLK_c, D => EF_c, SET => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.EFS_net_1\);
    
    \I3.VDBOFFA_31_IV_0L2R_2599\ : OR3
      port map(A => \I3.VDBoffa_31l2r_adt_net_164267_\, B => 
        \I3.VDBoffa_31l2r_adt_net_164263_\, C => 
        \I3.VDBoffa_31l2r_adt_net_164264_\, Y => 
        \I3.VDBoffa_31l2r_adt_net_164270_\);
    
    \I3.PIPEA1_12l19r\ : AND2
      port map(A => DPR_cl19r, B => 
        \I3.N_243_4_adt_net_1290__adt_net_854496__net_1\, Y => 
        \I3.PIPEA1_12l19r_net_1\);
    
    \I1.REG_74_0_ivl186r\ : AO21
      port map(A => \REGl186r\, B => \I1.N_57_268\, C => 
        \I1.REG_74l186r_adt_net_131785_\, Y => \I1.REG_74l186r\);
    
    \I3.VDBI_10_I_M2L5R_2240\ : AND2FT
      port map(A => \I3.REGMAPL2R_737\, B => \I3.REGMAPL1R_724\, 
        Y => \I3.N_283_adt_net_143533_\);
    
    \I3.VDBoff_4_i_il5r\ : MUX2L
      port map(A => \I3.VDBoffbl5r_net_1\, B => 
        \I3.VDBoffal5r_net_1\, S => 
        \I3.N_178_adt_net_1360__net_1\, Y => \I3.N_77\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I142_Y_0_a2_1_1\ : AND2
      port map(A => \I2.N_67\, B => \I2.N_17_0\, Y => 
        \I2.N_108_0_adt_net_55153_\);
    
    \I2.PIPE1_DTl14r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_741_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl14r_net_1\);
    
    \I2.WREi_794\ : AO21
      port map(A => \I2.WREi_net_1\, B => 
        \I2.un1_DTO_cl_1_sqmuxa_2\, C => \I2.N_4203\, Y => 
        \I2.WREi_794_net_1\);
    
    \I2.CRC32l28r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_823_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l28r_net_1\);
    
    \I3.un29_reg_ads_0_a2_0_a2_0\ : AND2FT
      port map(A => \I3.VASl4r_net_1\, B => \I3.VASl2r_net_1\, Y
         => \I3.N_550\);
    
    \I3.un224_reg_ads_0_a2_3_a2_1\ : NAND2
      port map(A => \I3.N_552\, B => \I3.N_550\, Y => \I3.N_578\);
    
    \I2.ADEl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l9r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl9r);
    
    \I1.REG_74_8_0_o4_0l380r\ : NAND2
      port map(A => \I1.N_1366\, B => \I1.N_1367_i\, Y => 
        \I1.N_396\);
    
    \I2.CRC32_12_i_0_x2l31r\ : XOR2FT
      port map(A => \I2.CRC32l31r_net_1\, B => \I2.N_232_i_i\, Y
         => \I2.N_244_i_i_0\);
    
    \I3.VDBil19r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_359_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil19r_net_1\);
    
    \I1.REG_0_sqmuxa_i_0_o2_0_838\ : AND3FFT
      port map(A => \I1.BYTECNT_307_net_1\, B => 
        \I1.BYTECNT_308_net_1\, C => 
        \I1.N_304_adt_net_105325_Ra1_\, Y => \I1.N_304_RA1__216\);
    
    \I5.COMMAND_52\ : MUX2H
      port map(A => \I5.COMMANDl15r_net_1\, B => 
        \I5.COMMAND_4l15r_net_1\, S => \I5.sstate1l13r_net_1\, Y
         => \I5.COMMAND_52_net_1\);
    
    \I3.un17_reg_ads_0_a2_3_a3\ : NOR3
      port map(A => \I3.N_547\, B => \I3.N_551\, C => \I3.N_581\, 
        Y => \I3.un17_reg_ads_0_a2_3_a3_net_1\);
    
    \I1.sstate_ns_1_iv_0_i_o2l8r\ : AO21TTF
      port map(A => \I1.N_324\, B => \I1.BITCNTl2r_net_1\, C => 
        \I1.sstatel0r_net_1\, Y => \I1.N_368\);
    
    \I3.VDBi_31l31r\ : MUX2L
      port map(A => \I3.REGl164r\, B => \I3.VDBi_20l31r\, S => 
        \I3.REGMAPl17r_adt_net_854284__net_1\, Y => 
        \I3.VDBi_31l31r_net_1\);
    
    \I2.TRGSERV_2_I_18\ : XOR2
      port map(A => \I2.DWACT_ADD_CI_0_g_array_1_0l0r\, B => 
        \I2.TRGSERVl2r_net_1\, Y => \I2.TRGSERV_2l2r\);
    
    \I2.N434_adt_net_3677_\ : OAI21FTF
      port map(A => \I2.N457\, B => \I2.N327\, C => \I2.N326\, Y
         => \I2.N434_adt_net_3677__net_1\);
    
    \I3.VDBOFFB_30_IV_0L1R_2464\ : AO21
      port map(A => \REGl334r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l1r_adt_net_162888_\, Y => 
        \I3.VDBoffb_30l1r_adt_net_162929_\);
    
    \I2.LEAD_FLAG6_640_1603\ : NOR2FT
      port map(A => LEAD_FLAGl3r, B => \I2.N_4527\, Y => 
        \I2.LEAD_FLAG6_640_adt_net_64292_\);
    
    \I1.un1_sbyte13_2_i_i_a2_i\ : OR2FT
      port map(A => \I1.N_436_i_i\, B => 
        \I1.N_223_adt_net_108707_\, Y => \I1.N_223\);
    
    \I0.EV_RESF2\ : DFFC
      port map(CLK => CLK_c, D => \I0.EV_RESF1_net_1\, CLR => 
        \I0.un4_hwresi_i\, Q => \I0.EV_RESF2_net_1\);
    
    \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__2832\ : OR3FFT
      port map(A => \I2.N_2870\, B => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854628__net_1\, 
        C => \I2.un1_DTE_1_sqmuxa_2_1_adt_net_35789__net_1\, Y
         => \I2.UN1_DTE_1_SQMUXA_2_1_ADT_NET_775__176\);
    
    \I2.MIC_ERR_REGS_344\ : MUX2H
      port map(A => \I2.MIC_ERR_REGSl15r_net_1\, B => 
        \I2.MIC_ERR_REGSl16r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_344_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL9R_1467\ : AND2FT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855664__net_1\, 
        B => \I2.PIPE1_DT_12l9r_net_1\, Y => 
        \I2.PIPE1_DT_42l9r_adt_net_50183_\);
    
    \I2.un2_evnt_word_I_16_959\ : AND3
      port map(A => \I2.WOFFSETl0r_net_1\, B => \I2.WOFFSETl1r\, 
        C => \I2.WOFFSETl2r\, Y => \I2.DWACT_FINC_E_0L0R_337\);
    
    \I3.VDBml3r\ : MUX2L
      port map(A => \I3.VDBil3r_net_1\, B => \I3.N_145\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml3r_net_1\);
    
    \I3.PIPEBl22r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_101_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl22r_net_1\);
    
    IACKOUTB_pad : OB33PH
      port map(PAD => IACKOUTB, A => \VCC\);
    
    \I2.G_EVNT_NUMl9r\ : DFFC
      port map(CLK => CLK_c, D => \I2.G_EVNT_NUM_925_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.G_EVNT_NUMl9r_net_1\);
    
    \I2.W_ERR_WORDS_327\ : OA21TTF
      port map(A => \I2.W_ERR_WORDS_net_1\, B => 
        \I2.STATE1l1r_net_1\, C => \I2.STATE1l17r_net_1\, Y => 
        \I2.W_ERR_WORDS_327_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A4_0_1564\ : OA21
      port map(A => \I2.N_152_i_0_adt_net_610537_\, B => 
        \I2.N_152_i_0_adt_net_610543_\, C => \I2.N_20_i_0\, Y => 
        \I2.N_41_0_adt_net_55923_\);
    
    \I2.WOFFSET_13_il12r\ : AND2
      port map(A => \I2.I_73\, B => \I2.N_4262\, Y => \I2.N_4255\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I151_Y_I_A2_2_2695\ : AO21
      port map(A => \I2.PIPE4_DTL10R_792\, B => 
        \I2.N_152_i_0_adt_net_502367_\, C => \I2.RAMDT4L12R_829\, 
        Y => \I2.N_152_i_0_adt_net_502321_\);
    
    \I2.RAMAD1_662\ : MUX2L
      port map(A => \I2.RAMAD1_12l8r_net_1\, B => 
        \I2.RAMAD1l8r_net_1\, S => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__172\, Y => 
        \I2.RAMAD1_662_net_1\);
    
    \I2.FID_7_0_ivl22r\ : AO21
      port map(A => \I2.STATE3L3R_416\, B => \I2.DTESl22r_net_1\, 
        C => \I2.FID_7l22r_adt_net_19311_\, Y => \I2.FID_7l22r\);
    
    \I2.DTOSl11r\ : DFF
      port map(CLK => CLK_c, D => DTO_inl11r, Q => 
        \I2.DTOSl11r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I54_Y\ : AO21
      port map(A => \I2.N270_0\, B => \I2.N304_0_adt_net_87004_\, 
        C => \I2.N304_0_adt_net_86999_\, Y => \I2.N304_0\);
    
    \I2.N_3279_0_adt_net_855236_\ : BFR
      port map(A => \I2.N_3279_0\, Y => 
        \I2.N_3279_0_adt_net_855236__net_1\);
    
    \I3.VDBOFFB_30_IV_0L6R_2375\ : AO21
      port map(A => \REGl323r\, B => \I3.REGMAPl37r_net_1\, C => 
        \I3.VDBoffb_30l6r_adt_net_161942_\, Y => 
        \I3.VDBoffb_30l6r_adt_net_161980_\);
    
    \I2.DT_SRAMl26r\ : MUX2L
      port map(A => \I2.N_894\, B => \I2.PIPE2_DTl26r_net_1\, S
         => \I2.N_4646_1_ADT_NET_1645_RD1__27\, Y => 
        \I2.DT_SRAMl26r_net_1\);
    
    \I5.REG_1l437r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_20_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl437r);
    
    \I2.SUB9_1_ADD_18x18_fast_I94_un1_Y\ : AND2
      port map(A => \I2.N340\, B => \I2.N333\, Y => 
        \I2.I94_un1_Y\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_A2_2_1543\ : AO21
      port map(A => \I2.PIPE4_DTL6R_480\, B => 
        \I2.PIPE4_DTL7R_481\, C => \I2.RAMDT4L5R_810\, Y => 
        \I2.N_128_adt_net_54290_\);
    
    \I2.FID_7_0_IVL6R_1720\ : AND2
      port map(A => \I2.STATE3L2R_414\, B => \I2.DTOSl6r_net_1\, 
        Y => \I2.FID_7l6r_adt_net_92927_\);
    
    REGl346r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_247_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl346r\);
    
    \I2.TDCDASl0r\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDA_cl0r, Q => 
        \I2.TDCDASl0r_net_1\);
    
    \I2.MAJORITY_REG_IL0R_1748\ : OA21
      port map(A => \I2.MIC_REG3l0r_net_1\, B => 
        \I2.MIC_REG2l0r_net_1\, C => \I2.MIC_REG1l0r_net_1\, Y
         => \reg_il0r_adt_net_105174_\);
    
    \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854400_\ : BFR
      port map(A => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854404__net_1\, 
        Y => 
        \I1.PAGECNT_0l8r_adt_net_834720_Rd1__adt_net_854400__net_1\);
    
    \I3.VDBi_29_0_a2_0l9r_883\ : NOR3FTT
      port map(A => \I3.REGMAPL2R_737\, B => \I3.REGMAPL7R_460\, 
        C => \I3.N_1907_263\, Y => \I3.N_2040_261\);
    
    \I2.PIPE1_DT_42_1_ivl27r\ : OA21TTF
      port map(A => \I2.PIPE1_DT_42_3_0l28r\, B => 
        \I2.EVNT_NUMl11r_net_1\, C => 
        \I2.PIPE1_DT_42_1_iv_2_il27r\, Y => 
        \I2.PIPE1_DT_42_1_iv_i_0l27r\);
    
    \I3.PIPEA1l30r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEA1_328_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l30r_net_1\);
    
    \I3.un1_STATE2_11_0_0\ : OR2
      port map(A => \I3.un1_STATE2_15_1_adt_net_3723__net_1\, B
         => \I3.un1_STATE2_11_adt_net_153728_\, Y => 
        \I3.un1_STATE2_11\);
    
    \I3.VDBi_31l14r\ : MUX2L
      port map(A => \I3.REGl147r\, B => \I3.VDBi_20l14r\, S => 
        \I3.REGMAPl17r_adt_net_854288__net_1\, Y => 
        \I3.VDBi_31l14r_net_1\);
    
    \I3.REGMAPl15r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un60_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAP_i_0_il15r\);
    
    \I2.TOKENA_TIMOUT_2\ : AND3
      port map(A => \I2.N_3899\, B => \I2.TOKENA_CNTl1r_net_1\, C
         => \I2.TOKENA_CNTl0r_net_1\, Y => 
        \I2.TOKENA_TIMOUT_2_net_1\);
    
    \I2.RAMDT4L12R_3044\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_798\);
    
    \I3.VADm_0_a3l22r\ : AND2FT
      port map(A => \I3.N_264_0_adt_net_1653_Rd1__net_1\, B => 
        \I3.PIPEAl22r_net_1\, Y => \I3.VADml22r\);
    
    \I2.DTE_cl_0_sqmuxa_2_adt_net_19952_\ : MUX2L
      port map(A => \I2.NWPIPE5_577\, B => \I2.NWPIPE10_net_1\, S
         => \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_stt_m3_net_1\, Y
         => \I2.DTE_cl_0_sqmuxa_2_adt_net_19952__net_1\);
    
    \I2.DTO_16_1_IV_0_0L12R_1159\ : AO21
      port map(A => \I2.STATE2l4r_adt_net_855688__net_1\, B => 
        \I2.N_3966\, C => \I2.DTO_16_1l12r_adt_net_32622_\, Y => 
        \I2.DTO_16_1l12r_adt_net_32632_\);
    
    \I3.N_57_i_0_0_adt_net_854696_\ : BFR
      port map(A => \I3.N_57_i_0_0_adt_net_854700__net_1\, Y => 
        \I3.N_57_i_0_0_adt_net_854696__net_1\);
    
    \I2.MIC_ERR_REGS_376\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl48r_net_1\, B => 
        \I2.MIC_ERR_REGSl47r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_376_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL29R_1357\ : NAND3
      port map(A => \I2.N_3254\, B => 
        \I2.N_3234_adt_net_855652__net_1\, C => 
        \I2.PIPE1_DT_42_1l29r\, Y => 
        \I2.PIPE1_DT_42l29r_adt_net_45836_\);
    
    \I2.BNCID_VECT_tile_0_DIN_REG1l2r\ : DFF
      port map(CLK => CLK_c, D => \I2.BNC_IDl10r_net_1\, Q => 
        \I2.DIN_REG1l2r\);
    
    \I2.ADEl11r\ : DFFC
      port map(CLK => CLK_c, D => \I2.ADE_4l11r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => ADE_cl11r);
    
    LWORDB_pad : IOB33PH
      port map(PAD => LWORDB, A => \I3.VADml0r\, EN => 
        NOEAD_c_i_0, Y => LWORDB_in);
    
    \I2.PIPE1_DTl22r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_749_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl22r_net_1\);
    
    \I1.REG_17_sqmuxa_0_a2_0_a3_0_a2\ : NAND2
      port map(A => \I1.N_590_228\, B => 
        \I1.PAGECNTl9r_adt_net_854816__net_1\, Y => \I1.N_260\);
    
    \I2.OFFSET_37_7l2r\ : MUX2L
      port map(A => \I2.N_677\, B => \I2.N_653\, S => 
        \I2.PIPE7_DTL25R_683\, Y => \I2.N_685\);
    
    \I3.VDBm_0l10r\ : MUX2L
      port map(A => \I3.PIPEAl10r_net_1\, B => 
        \I3.PIPEBl10r_net_1\, S => \I3.BLTCYC_net_1\, Y => 
        \I3.N_152\);
    
    \I1.REG_74_2_0l404r_Rd1_\ : DFFS
      port map(CLK => CLK_c, D => \I1.REG_74_2_0l404r_Ra1_\, SET
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I1.REG_74_2_0l404r_Rd1__net_1\);
    
    \I2.SUB9_1_ADD_18x18_fast_I6_P0N\ : OR2
      port map(A => \I2.N_3545_i_i\, B => \I2.G_1\, Y => 
        \I2.N244\);
    
    \I1.SBYTE_8_0_IL6R_1754\ : OA21TTF
      port map(A => \I1.N_603_i\, B => \FBOUTl5r\, C => 
        \I1.N_337\, Y => \I1.N_206_adt_net_105994_\);
    
    \I5.BITCNT_84\ : MUX2H
      port map(A => \I5.BITCNTl2r_net_1\, B => 
        \I5.N_54_adt_net_9598_\, S => \I5.BITCNTe\, Y => 
        \I5.BITCNT_84_net_1\);
    
    \I2.TOKENB_CNTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.TOKENB_CNT_3l0r\, CLR => 
        \I2.un12_clear_stat_i\, Q => \I2.TOKENB_CNTl0r_net_1\);
    
    \I3.TCNT3_i_0_il0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT3_379_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT3_i_0_il0r_net_1\);
    
    \I2.DTO_16_1_IV_0L24R_1096\ : AO21
      port map(A => \I2.DTO_1l24r\, B => \I2.N_196_53\, C => 
        \I2.DTO_16_1l24r_adt_net_29854_\, Y => 
        \I2.DTO_16_1l24r_adt_net_29870_\);
    
    \I3.REGMAP_i_0_a2l52r_739\ : NOR3FFT
      port map(A => \I3.UN1_REGMAP_34_124\, B => 
        \I3.N_638_adt_net_134647_\, C => \I3.N_2017_119\, Y => 
        \I3.N_638_117\);
    
    \I3.REG_1_220\ : MUX2L
      port map(A => VDB_inl7r, B => REGl413r, S => 
        \I3.REG_0_sqmuxa_3\, Y => \I3.REG_1_220_0\);
    
    \I2.MIC_REG1_i_il6r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG1_307_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG1_i_il6r_net_1\);
    
    \I2.WOFFSETl9r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.WOFFSETl9r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WOFFSETl9r_Rd1__net_1\);
    
    \I2.PIPE8_DT_558\ : OAI21TTF
      port map(A => \I2.N_4707_i_0\, B => 
        \I2.PIPE8_DT_21_i_0_il30r\, C => 
        \I2.PIPE8_DT_558_adt_net_82590_\, Y => 
        \I2.PIPE8_DT_558_net_1\);
    
    \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_784\ : NOR3
      port map(A => \I2.N_4646_1_adt_net_19635__net_1\, B => 
        \I2.N_4646_1_adt_net_19637_Rd1__net_1\, C => 
        \I2.END_EVNT2_404\, Y => 
        \I2.STATE2_3_SQMUXA_0_A2_0_A2_0_A2_0_3_ADT_NET_19813__162\);
    
    \I2.MIC_ERR_REGS_361\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl33r_net_1\, B => 
        \I2.MIC_ERR_REGSl32r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855848__net_1\, Y => 
        \I2.MIC_ERR_REGS_361_net_1\);
    
    \I1.REG_74l220r_787\ : OR3
      port map(A => \I1.N_89_adt_net_128732_\, B => 
        \I1.N_97_6_adt_net_854712__net_1\, C => 
        \I1.N_89_adt_net_128736_\, Y => \I1.N_89_165\);
    
    \I3.N_243_4_adt_net_1290__adt_net_854500_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854512__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854500__net_1\);
    
    \I2.DT_SRAM_0l0r\ : MUX2L
      port map(A => \I2.PIPE10_DTl0r_net_1\, B => 
        \I2.PIPE5_DTl0r_net_1\, S => 
        \I2.REG_0l3r_adt_net_848__adt_net_854204__net_1\, Y => 
        \I2.N_868\);
    
    \I2.MIC_ERR_REGS_369\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl41r_net_1\, B => 
        \I2.MIC_ERR_REGSl40r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855844__net_1\, Y => 
        \I2.MIC_ERR_REGS_369_net_1\);
    
    \I2.DTO_16_1_IV_1L3R_1203\ : NOR2
      port map(A => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854608__net_1\, 
        B => \I2.DT_TEMPl3r_net_1\, Y => 
        \I2.DTO_16_1_iv_1l3r_adt_net_34602_\);
    
    DPR_padl17r : IB33
      port map(PAD => DPR(17), Y => DPR_cl17r);
    
    \I2.REG_1l38r_1767\ : DFFC
      port map(CLK => CLK_c, D => \I2.REG_1_n6_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => REGL38R_873);
    
    TDCDB_padl3r : IB33
      port map(PAD => TDCDB(3), Y => TDCDB_cl3r);
    
    \I1.SBYTE_8_0_a2_i_m2l2r\ : MUX2L
      port map(A => \FBOUTl1r\, B => REGl85r, S => 
        \I1.sstatel2r_net_1\, Y => \I1.N_1385\);
    
    \I1.PAGECNT_n6_i_i_a4_0_827\ : OR2FT
      port map(A => \I1.UN1_SBYTE13_1_I_1_209\, B => 
        \I1.N_656_496\, Y => \I1.N_473_205\);
    
    \I3.un1_STATE2_11_adt_net_1401_\ : NAND3FFT
      port map(A => DPR_cl29r, B => 
        \I3.un1_STATE2_11_adt_net_153679__net_1\, C => DPR_cl28r, 
        Y => \I3.un1_STATE2_11_adt_net_1401__net_1\);
    
    \I2.UN1_DTO_CL_1_SQMUXA_2_0_O2_1018\ : AO21FTF
      port map(A => \I2.N_4241_1\, B => \I2.STATE2l5r_net_1\, C
         => 
        \I2.DTO_cl_1_sqmuxa_adt_net_1022__adt_net_854604__net_1\, 
        Y => \I2.un1_DTO_cl_1_sqmuxa_2_adt_net_22202_\);
    
    \I3.VDBOFFB_30_IV_0L3R_2422\ : AND2
      port map(A => \REGl376r\, B => \I3.REGMAPl44r_net_1\, Y => 
        \I3.VDBoffb_30l3r_adt_net_162512_\);
    
    \I3.VDBoff_121\ : MUX2L
      port map(A => \I3.VDBoffl5r_net_1\, B => \I3.N_77\, S => 
        \I3.un1_REGMAP_34\, Y => \I3.VDBoff_121_net_1\);
    
    \I2.LSRAM_IN_408\ : MUX2L
      port map(A => \I2.PIPE5_DTl24r_net_1\, B => 
        \I2.LSRAM_INl24r_net_1\, S => 
        \I2.LEAD_FLAG6_0_sqmuxa_1_1\, Y => 
        \I2.LSRAM_IN_408_net_1\);
    
    \I1.BITCNTlde_i_a2_0_a4\ : AO21
      port map(A => \I1.N_329\, B => \I1.N_346\, C => 
        \PULSEl0r_adt_net_854536__net_1\, Y => \I1.N_457\);
    
    \I2.WPAGEl13r\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_950_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEl13r_net_1\);
    
    \I2.REG_1_n6_0\ : XOR2FT
      port map(A => \I2.un8_evread_1_adt_net_855784__net_1\, B
         => REGl38r, Y => \I2.REG_1_n6_0_net_1\);
    
    \I2.MSERCLKS\ : DFFC
      port map(CLK => CLK_c, D => \I2.MSERCLKF1_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I2.MSERCLKS_net_1\);
    
    \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__2764\ : NAND3FFT
      port map(A => \I2.ENDF_net_1\, B => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_20149__net_1\, C => 
        \I2.STATE2_3_sqmuxa_0_a2_0_a2_0_a2_0_3_net_1\, Y => 
        \I2.DTO_16_1_IV_0_A2_2_0L21R_ADT_NET_1014__47\);
    
    \I3.VDBml30r\ : MUX2L
      port map(A => \I3.VDBil30r_net_1\, B => \I3.N_172\, S => 
        \I3.SINGCYC_net_1\, Y => \I3.VDBml30r_net_1\);
    
    \I0.REG_1_3\ : OR2
      port map(A => REGl27r, B => TICKL0R_558, Y => 
        \I0.REG_1_3_net_1\);
    
    \I1.REG_1_252\ : MUX2H
      port map(A => \REGl351r\, B => \I1.REG_74l351r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_252_net_1\);
    
    \I1.BITCNT_316\ : MUX2L
      port map(A => \I1.BITCNTl1r_net_1\, B => \I1.N_416\, S => 
        \I1.N_68\, Y => \I1.BITCNT_316_net_1\);
    
    \I3.VDBi_57_iv_0_0_a2_16l0r\ : AND3FFT
      port map(A => \I3.N_2017\, B => 
        \I3.REGMAPl9r_adt_net_854308__net_1\, C => \I3.N_590\, Y
         => \I3.N_2036\);
    
    \I2.LSRAM_RD\ : MUX2L
      port map(A => LSRAM_FL_RD, B => \I2.LSRAM_RDi_net_1\, S => 
        FLUSH, Y => \I2.LSRAM_RD_net_1\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2280\ : AO21
      port map(A => \I3.N_2037\, B => \I3.N_132\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146422_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146447_\);
    
    \I1.REG_74_0_iv_i_a3l205r\ : OR2
      port map(A => \I1.N_181\, B => \I1.REG_5_sqmuxa\, Y => 
        \I1.N_183_i_0\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I136_Y_0_O2_M2_E_1569\ : 
        AND3
      port map(A => \I2.ADD_21x21_fast_I140_Y_0_a2_0_0_0\, B => 
        \I2.N_20_i_0\, C => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_N_6_i_adt_net_56543_\, Y
         => \I2.ADD_21x21_fast_I136_Y_0_o2_N_6_i_adt_net_56545_\);
    
    \I2.ROFFSET_n6\ : NOR2
      port map(A => 
        \I2.N_1170_adt_net_1217__adt_net_855696__net_1\, B => 
        \I2.ROFFSET_n6_tz_i\, Y => \I2.ROFFSET_n6_net_1\);
    
    \I2.PIPE8_DT_21_I_1L28R_1673\ : OAI21FTF
      port map(A => \I2.PIPE7_DTl30r_adt_net_855172__net_1\, B
         => \I2.PIPE7_DTl28r_net_1\, C => \I2.NWPIPE7_689\, Y => 
        \I2.PIPE8_DT_21_i_1l28r_adt_net_82784_\);
    
    \I2.DTO_9_IVL22R_1104\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996__net_1\, 
        B => \I2.G_EVNT_NUMl6r_net_1\, Y => 
        \I2.DTO_9l22r_adt_net_30286_\);
    
    \I1.REG_74_0_IVL276R_1947\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_14_sqmuxa_adt_net_855436__net_1\, Y => 
        \I1.REG_74l276r_adt_net_123302_\);
    
    \I2.PIPE1_DTl3r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.PIPE1_DT_730_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.PIPE1_DTl3r_net_1\);
    
    \I2.TOKENTOA_RES\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => 
        \I2.TOKENTOA_RES_648_net_1\, CLR => CLEAR_STAT_i_0, Q => 
        \I2.TOKENTOA_RES_net_1\);
    
    \I2.PIPE6_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DT_473_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE6_DTl19r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I173_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l10r_net_1\, B => 
        \I2.PIPE4_DTl3r_adt_net_854544__net_1\, Y => 
        \I2.ADD_21x21_fast_I173_Y_0_0\);
    
    \I2.SUB9_1_ADD_18x18_fast_I30_Y\ : AND2FT
      port map(A => \I2.SUB8l14r_adt_net_855568__net_1\, B => 
        \I2.N295_adt_net_68996_\, Y => \I2.N295\);
    
    \I3.VDBi_23l1r_adt_net_145526_\ : AND2
      port map(A => REGl49r, B => 
        \I3.REGMAPl9r_adt_net_854332__net_1\, Y => 
        \I3.VDBi_23l1r_adt_net_145526__net_1\);
    
    \I1.REG_9_sqmuxa_0_a2_1_0_a2\ : OR2
      port map(A => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__382\, 
        B => \I1.REG_74_1_380_M8_I_0_RD1__336\, Y => \I1.N_1169\);
    
    \I1.REG_74_1_0_il188r\ : NAND3FFT
      port map(A => 
        \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_2_0_ADT_NET_1417_RD1__198\, 
        B => \I1.REG_74_4_i_a2_404_N_4_i_adt_net_1465__net_1\, C
         => \I1.REG_74_9_0_o4_a0_2l372r\, Y => 
        \I1.REG_74_4_i_a2_404_N_4_i\);
    
    \I1.REG_74_0_IVL342R_1871\ : AND2
      port map(A => \FBOUTl1r\, B => 
        \I1.REG_23_sqmuxa_adt_net_855512__net_1\, Y => 
        \I1.REG_74l342r_adt_net_116842_\);
    
    \I3.TCNT2_i_0_il0r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT2_396_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT2_i_0_il0r_net_1\);
    
    \I2.PIPE7_DTl19r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl19r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl19r_net_1\);
    
    \I1.REG_1_254\ : MUX2H
      port map(A => \REGl353r\, B => \I1.REG_74l353r\, S => 
        \I1.N_50_0_ADT_NET_1409__20\, Y => \I1.REG_1_254_net_1\);
    
    \I2.UN1_CHAIN_RDY_1_SQMUXA_I_1708\ : AO21FTT
      port map(A => \I2.CHAIN_ERRS_net_1\, B => \I2.STATEe_ipl2r\, 
        C => \I2.N_3494_adt_net_90556_\, Y => 
        \I2.N_3494_adt_net_90563_\);
    
    \I2.DT_TEMP_766\ : MUX2L
      port map(A => \I2.DT_TEMP_7l5r_net_1\, B => 
        \I2.DT_TEMPl5r_net_1\, S => 
        \I2.UN1_STATE2_3_SQMUXA_1_ADT_NET_839__28\, Y => 
        \I2.DT_TEMP_766_net_1\);
    
    \I2.DTO_16_1_iv_0_o7l29r\ : AO21FTT
      port map(A => \I2.N_4283_i_0\, B => \I2.DT_TEMPl29r_net_1\, 
        C => \I2.N_4159_adt_net_28676_\, Y => \I2.N_4159\);
    
    \I3.VDBOFFA_31_IV_I_A2_IL6R_2522\ : AO21
      port map(A => \REGl267r\, B => \I3.REGMAP_i_0_il30r_net_1\, 
        C => \I3.N_2070_adt_net_163474_\, Y => 
        \I3.N_2070_adt_net_163503_\);
    
    \I2.REG_1l81r\ : DFFC
      port map(CLK => MROK_c, D => \VCC\, CLR => \I2.un3_hwres_i\, 
        Q => REGl81r);
    
    REGl366r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_267_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl366r\);
    
    \I2.STATE2l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.STATE2_nsl2r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE2l3r_net_1\);
    
    \I3.VDBOFFB_30_IV_0L2R_2454\ : OR3
      port map(A => \I3.VDBoffb_30l2r_adt_net_162745_\, B => 
        \I3.VDBoffb_30l2r_adt_net_162739_\, C => 
        \I3.VDBoffb_30l2r_adt_net_162740_\, Y => 
        \I3.VDBoffb_30l2r_adt_net_162749_\);
    
    DPR_padl12r : IB33
      port map(PAD => DPR(12), Y => DPR_cl12r);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I173_Y_0\ : XOR2
      port map(A => \I2.RAMDT4l3r_net_1\, B => 
        \I2.PIPE4_DTl3r_adt_net_854544__net_1\, Y => 
        \I2.ADD_21x21_fast_I173_Y_0\);
    
    \I2.PIPE7_DTl20r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE6_DTl20r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE7_DTl20r_net_1\);
    
    \I2.DT_TEMP_768\ : MUX2H
      port map(A => \I2.DT_TEMPl7r_net_1\, B => 
        \I2.DT_TEMP_7l7r_net_1\, S => 
        \I2.un1_STATE2_3_sqmuxa_1_adt_net_839__net_1\, Y => 
        \I2.DT_TEMP_768_net_1\);
    
    \I2.PIPE9_DT_294\ : MUX2L
      port map(A => \I2.PIPE9_DTl25r_net_1\, B => 
        \I2.PIPE8_DTl25r_net_1\, S => \I2.NWPIPE8_I_0_I_0_0_5\, Y
         => \I2.PIPE9_DT_294_net_1\);
    
    \I2.PIPE1_DT_42_1_IVL15R_1429\ : AND2
      port map(A => \I2.STATE1l3r_net_1\, B => 
        \I2.MIC_ERR_REGSl31r_net_1\, Y => 
        \I2.PIPE1_DT_42l15r_adt_net_48697_\);
    
    \I2.EVNT_WORDl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_WORD_713_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_WORDl0r_net_1\);
    
    \I2.ADO_3l0r\ : MUX2L
      port map(A => \I2.WOFFSETl1r_adt_net_854992__net_1\, B => 
        \I2.ROFFSETl1r_net_1\, S => NOESRAME_c, Y => 
        \I2.ADO_3l0r_net_1\);
    
    \I2.STATEE_ILLEGAL_1029\ : AO21
      port map(A => \I2.STATEe_ipl1r\, B => \I2.N_3450\, C => 
        \I2.N_3457_ip_adt_net_23079_\, Y => 
        \I2.N_3457_ip_adt_net_23080_\);
    
    \I3.PIPEAl30r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEA_261_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEAl30r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I171_Y\ : XOR2FT
      port map(A => \I2.N_85_0\, B => 
        \I2.ADD_21x21_fast_I171_Y_0_0\, Y => 
        \I2.un27_pipe5_dt1l1r\);
    
    \I5.REG_1l439r\ : DFFC
      port map(CLK => CLK_c, D => \I5.REG_1_22_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl439r);
    
    \I3.VDBOFFB_30_IV_0L0R_2475\ : AND2
      port map(A => \REGl349r\, B => \I3.REGMAPl41r_net_1\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163078_\);
    
    \I2.CRC32_12_i_m2l4r\ : MUX2L
      port map(A => \I2.DT_TEMPl4r_net_1\, B => 
        \I2.DT_SRAMl4r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854440__net_1\, Y => 
        \I2.N_3955_i_i\);
    
    \I3.REG_1l66r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_167_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl66r);
    
    \I1.REG_74_0_IVL308R_1910\ : AND2
      port map(A => \I1.FBOUTl7r_net_1\, B => 
        \I1.REG_18_sqmuxa_adt_net_855476__net_1\, Y => 
        \I1.REG_74l308r_adt_net_120180_\);
    
    \I3.REGMAPl39r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un176_reg_ads_0_a2_0_a3_net_1\, Q => 
        \I3.REGMAPl39r_net_1\);
    
    \I2.SUB9_585\ : MUX2H
      port map(A => \I2.SUB9_i_0_il17r\, B => \I2.SUB9_1l17r\, S
         => \I2.SUB9_0_sqmuxa_0\, Y => \I2.SUB9_585_net_1\);
    
    \I1.REG_0_sqmuxa_i_0_a4_1_905\ : NAND2
      port map(A => \I1.N_598_23\, B => 
        \I1.sstate_ns_il5r_adt_net_107266_\, Y => 
        \I1.N_435_1_283\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I37_P0N\ : OR2FT
      port map(A => \I2.LSRAM_OUTl16r\, B => 
        \I2.PIPE7_DTl16r_net_1\, Y => \I2.N279\);
    
    \I2.RMIC_i\ : OR2
      port map(A => \HWRES_3_ADT_NET_738__17\, B => PULSEL4R_15, 
        Y => \I2.un8_hwres_i\);
    
    \I3.un1_STATE2_13_adt_net_1333__adt_net_854652_\ : BFR
      port map(A => \I3.un1_STATE2_13_adt_net_1333__net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_1333__adt_net_854652__net_1\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2282\ : AO21FTT
      port map(A => \I3.N_2017\, B => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146304_\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146420_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146450_\);
    
    \I5.sstate1se_9_i_0_m4\ : MUX2L
      port map(A => \I5.sstate1l4r_net_1\, B => 
        \I5.sstate1l3r_net_1\, S => TICKL0R_558, Y => \I5.N_96\);
    
    \I1.REG_74_i_o2_i_2l364r\ : AND3FTT
      port map(A => \I1.N_97_2\, B => \I1.N_273_9\, C => 
        \I1.N_273_10\, Y => \I1.N_57_9_i\);
    
    \I3.STATE1_nsl2r_adt_net_134736_\ : NOR3FFT
      port map(A => \I3.N_2083\, B => \I3.N_1641\, C => 
        \I3.STATE1_tr24_i_0_a3_28_tz_i\, Y => 
        \I3.STATE1_nsl2r_adt_net_134736__net_1\);
    
    \I2.TOKOUT_FL_1537\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.TOKOUT_FL_674_net_1\, 
        CLR => CLEAR_STAT_i_0, Q => \I2.TOKOUT_FL_644\);
    
    \I2.CRC32l27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.CRC32_822_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.CRC32l27r_net_1\);
    
    \I2.DTEST_FIFO_645\ : AO21FTT
      port map(A => \I2.STATE3l5r_net_1\, B => DTEST_FIFO, C => 
        \I2.STATE3l6r_net_1\, Y => \I2.DTEST_FIFO_645_net_1\);
    
    \I1.BYTECNT_310\ : MUX2H
      port map(A => \I1.BYTECNT_i_0_il4r_net_1\, B => \I1.N_1381\, 
        S => \I1.N_1383_224\, Y => \I1.BYTECNT_310_net_1\);
    
    \I2.MIC_ERR_REGSl39r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_368_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl39r_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I119_Y_I_O4_1583\ : AND2
      port map(A => \I2.RAMDT4L5R_821\, B => 
        \I2.N_3_adt_net_940__net_1\, Y => \I2.N_3_adt_net_59496_\);
    
    \I5.DATA_1_sqmuxa_2_0_a2_0_a2\ : OR2FT
      port map(A => TICKL0R_556, B => \I5.N_70\, Y => 
        \I5.DATA_1_sqmuxa_2\);
    
    \I2.un28_sram_empty_6_0\ : MUX2L
      port map(A => \I2.N_624\, B => \I2.N_623\, S => 
        \I2.RPAGEL14R_612\, Y => \I2.N_625\);
    
    ADE_padl5r : OB33PH
      port map(PAD => ADE(5), A => ADE_cl5r);
    
    \I3.PIPEA1_324\ : MUX2L
      port map(A => \I3.PIPEA1l26r_net_1\, B => 
        \I3.PIPEA1_12l26r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, Y => 
        \I3.PIPEA1_324_net_1\);
    
    \I3.un1_REGMAP_34_5_0_a2_i_o2_i_a2_2_o2\ : NOR3FTT
      port map(A => \I3.N_2086_adt_net_134541_\, B => 
        \I3.REGMAP_I_0_IL42R_531\, C => \I3.REGMAPL41R_530\, Y
         => \I3.N_2086\);
    
    \I5.un1_sstate2_3_0\ : OR2
      port map(A => \I5.sstate2l4r_net_1\, B => 
        \I5.un1_sstate2_3_0_adt_net_11182_\, Y => 
        \I5.un1_sstate2_3_0_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I152_Y_0_o2\ : AO21
      port map(A => \I2.N_2360_tz_tz\, B => 
        \I2.N507_adt_net_56246__net_1\, C => 
        \I2.N507_adt_net_347771__net_1\, Y => 
        \I2.N_147_0_adt_net_604832_\);
    
    \I3.VAS_70\ : MUX2L
      port map(A => VAD_inl8r, B => \I3.VASl8r_net_1\, S => 
        \I3.VSEL_0\, Y => \I3.VAS_70_net_1\);
    
    \I2.un2_evnt_word_I_24\ : XOR2
      port map(A => \I2.WOFFSETl5r\, B => \I2.N_39\, Y => 
        \I2.I_24\);
    
    \I2.PIPE6_DT_0_sqmuxa_i_m2_0\ : MUX2L
      port map(A => LEAD_FLAGl3r, B => LEAD_FLAGl1r, S => 
        \I2.PIPE5_DTL22R_666\, Y => \I2.N_4543\);
    
    \I3.un1_MYBERRi_1_sqmuxa_0_0\ : AO21
      port map(A => \I3.DSS_9\, B => \I3.STATE1_ipl4r\, C => 
        \I3.un1_MYBERRi_1_sqmuxa_adt_net_161480_\, Y => 
        \I3.un1_MYBERRi_1_sqmuxa\);
    
    \I2.DTO_9_IV_0L20R_1115\ : AND2
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_855004__net_1\, 
        B => \I2.G_EVNT_NUMl4r_net_1\, Y => 
        \I2.DTO_9l20r_adt_net_30718_\);
    
    \I3.PIPEBl2r\ : DFFC
      port map(CLK => CLK_c, D => \I3.PIPEB_81_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I3.PIPEBl2r_net_1\);
    
    \I2.DTE_21_1_IV_0L19R_1263\ : AND2
      port map(A => \I2.STATE2l1r_adt_net_855116__net_1\, B => 
        \I2.L_LUT_net_1\, Y => \I2.DTE_21_1l19r_adt_net_37709_\);
    
    DTE_padl17r : IOB33PH
      port map(PAD => DTE(17), A => \I2.DTE_1l17r\, EN => 
        \I2.N_4178_i_0_1\, Y => DTE_inl17r);
    
    DTO_padl20r : IOB33PH
      port map(PAD => DTO(20), A => \I2.DTO_1l20r\, EN => 
        \I2.N_4239_i_0_1\, Y => DTO_inl20r);
    
    \I2.PIPE1_DT_12l30r\ : OA21
      port map(A => \I2.un3_tdcgda1_1_adt_net_21664__net_1\, B
         => \I2.TDCDASl28r_net_1\, C => \I2.TDCDASl30r_net_1\, Y
         => \I2.PIPE1_DT_12l30r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I138_Y_0_0_1581\ : AND3
      port map(A => \I2.N_2358_tz_tz_adt_net_55567_\, B => 
        \I2.N_53_0\, C => 
        \I2.ADD_21x21_fast_I136_Y_0_o2_m4_e_i_1\, Y => 
        \I2.ADD_21x21_fast_I138_Y_0_0_0_adt_net_58684_\);
    
    \I1.REG_3_sqmuxa_0_a2_0_818_899\ : NAND2FT
      port map(A => \I1.PAGECNTL9R_244\, B => 
        \I1.N_238_Rd1__net_1\, Y => \I1.N_254_277\);
    
    \I3.VDBil23r\ : DFFC
      port map(CLK => CLK_c, D => \I3.VDBi_363_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I3.VDBil23r_net_1\);
    
    \I2.WOFFSET_839\ : MUX2L
      port map(A => \I2.WOFFSETl12r_Rd1__net_1\, B => 
        \I2.N_4255_Rd1__net_1\, S => 
        \I2.N_2828_adt_net_1062__adt_net_835304_Rd1__net_1\, Y
         => \I2.WOFFSETl12r\);
    
    \I4.bcnt_7\ : MUX2H
      port map(A => \I4.bcnt_i_0_il2r_net_1\, B => \I4.I_9\, S
         => \I4.STATE1l1r_net_1\, Y => \I4.bcnt_7_net_1\);
    
    \I2.DTO_16_1_iv_0_0l0r\ : OA21FTF
      port map(A => \I2.N_182_ADT_NET_1007__386\, B => 
        \I2.DT_SRAMl0r_net_1\, C => 
        \I2.DTO_16_1_iv_0_0_1l0r_net_1\, Y => \I2.DTO_16_1_ivl0r\);
    
    \I2.PIPE9_DTl31r_1560\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_300_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTL31R_667\);
    
    \I1.ISCK_0_sqmuxa_0_0_a2_0\ : AND3FFT
      port map(A => \I1.SSTATEL2R_758\, B => \I1.sstatel1r_net_1\, 
        C => \I1.N_628_adt_net_107115_\, Y => \I1.N_628\);
    
    TDCDB_padl20r : IB33
      port map(PAD => TDCDB(20), Y => TDCDB_cl20r);
    
    \I5.UN1_SSTATE2_3_0_923\ : AOI21TTF
      port map(A => REGl117r, B => \I5.AIR_START_net_1\, C => 
        \I5.sstate2l3r_net_1\, Y => 
        \I5.un1_sstate2_3_0_adt_net_11182_\);
    
    \I3.REG_1l67r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_168_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl67r);
    
    \I2.L2ARR_944\ : XOR2FT
      port map(A => \I2.N_4482_0\, B => \I2.L2ARRl0r_net_1\, Y
         => \I2.L2ARR_944_net_1\);
    
    \I2.FCNTl2r_1493\ : DFFS
      port map(CLK => \I2.CLK_tdc\, D => \I2.FCNT_945_net_1\, SET
         => CLEAR_STAT_i_0, Q => \I2.FCNTL2R_600\);
    
    \I2.PIPE1_DT_42_1_IVL0R_1524\ : AO21FTT
      port map(A => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855656__net_1\, 
        B => \I2.PIPE1_DT_12l0r_net_1\, C => 
        \I2.PIPE1_DT_42l0r_adt_net_52239_\, Y => 
        \I2.PIPE1_DT_42l0r_adt_net_52248_\);
    
    \I1.REG_16_sqmuxa_0_a2_m3_e_716\ : NAND3FFT
      port map(A => 
        \I1.un110_bitcnt_7_0_a2_0_a3_0_a2_2_0_adt_net_1417_Rd1__net_1\, 
        B => \I1.N_253_97\, C => \I1.REG_74_1_i_a2_a0_2l404r\, Y
         => \I1.REG_16_SQMUXA_94\);
    
    \I3.STATE1_TR24_59_1_I_A2_0_A2_0_A2_1_A2_2080\ : NOR3
      port map(A => \I3.REGMAPl23r_net_1\, B => 
        \I3.REGMAPL28R_535\, C => \I3.REGMAP_I_0_IL19R_534\, Y
         => \I3.N_68_adt_net_134367_\);
    
    \I2.EVNT_REJ\ : DFFC
      port map(CLK => CLK_c, D => \I2.EVNT_REJ_646_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.EVNT_REJ_net_1\);
    
    \I3.UN68_REG_ADS_0_A2_3_A3_2650\ : NOR3
      port map(A => \I3.LWORDS_net_1\, B => \I3.N_558\, C => 
        \I3.N_581\, Y => 
        \I3.un68_reg_ads_0_a2_3_a3_adt_net_166224_\);
    
    \I2.SUB9_1_ADD_18x18_fast_I146_Y\ : XOR2
      port map(A => \I2.N466\, B => \I2.ADD_18x18_fast_I146_Y_0\, 
        Y => \I2.SUB9_1l9r\);
    
    \I2.CRC32_12_i_0_m2l31r\ : MUX2L
      port map(A => \I2.DT_TEMPl31r_net_1\, B => 
        \I2.DT_SRAMl31r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854188__net_1\, Y => 
        \I2.N_232_i_i\);
    
    \I2.DTE_21_1l17r_Rd1_\ : DFFC
      port map(CLK => CLK_c, D => \I2.DTE_21_1l17r\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.DTE_21_1l17r_Rd1__net_1\);
    
    \I2.END_CHAINB1_709\ : AO21
      port map(A => \I2.STATE1l6r_net_1\, B => 
        \I2.END_CHAINB1_709_adt_net_2397__net_1\, C => 
        \I2.END_CHAINB1_709_adt_net_53463_\, Y => 
        \I2.END_CHAINB1_709_net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I152_Y_0_O2_2712\ : AND3
      port map(A => \I2.N_63\, B => \I2.N_33_adt_net_55020_\, C
         => \I2.N_147_0_adt_net_604832_\, Y => 
        \I2.N_147_0_adt_net_604875_\);
    
    \I2.PIPE5_DTl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE5_DT_697_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE5_DTl21r_net_1\);
    
    \I2.PIPE4_DTl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl0r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DTl0r_net_1\);
    
    \I2.MIC_ERR_REGSl21r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_350_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl21r_net_1\);
    
    \I2.RAMDT4l10r\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl10r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4l10r_net_1\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I139_Y_I_A4_2689\ : 
        OAI21FTT
      port map(A => \I2.N_2358_tz_tz\, B => 
        \I2.N522_0_adt_net_329169_\, C => 
        \I2.N522_0_adt_net_384644_\, Y => 
        \I2.N_96_0_adt_net_469923_\);
    
    \I1.REG_74_0_ivl169r\ : AO21
      port map(A => \REGl169r\, B => \I1.N_41\, C => 
        \I1.REG_74l169r_adt_net_133321_\, Y => \I1.REG_74l169r\);
    
    \I3.REG_1l89r\ : DFFC
      port map(CLK => CLK_c, D => \I3.REG_1_270_0\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => REGl89r);
    
    \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__2827\ : OAI21TTF
      port map(A => 
        \I2.un3_tdcgda1_1_adt_net_821__adt_net_855096__net_1\, B
         => 
        \I2.PIPE1_DT_2_sqmuxa_adt_net_803__adt_net_855660__net_1\, 
        C => \I2.FIRST_TDC_1_sqmuxa_net_1\, Y => 
        \I2.UN1_FIRST_TDC_1_SQMUXA_0_ADT_NET_1038__171\);
    
    \I3.STATE1l5r\ : DFFC
      port map(CLK => CLK_c, D => \I3.STATE1_nsl5r\, CLR => 
        \I3.N_1311_0\, Q => \I3.STATE1_ipl5r\);
    
    \I1.SBYTE_8_0_a2_il2r\ : AND2
      port map(A => \I1.N_371_i\, B => \I1.N_1385\, Y => 
        \I1.N_190\);
    
    VAD_padl11r : IOB33PH
      port map(PAD => VAD(11), A => \I3.VADml11r\, EN => 
        NOEAD_c_i_0, Y => VAD_inl11r);
    
    \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880_\ : BFR
      port map(A => \I5.SENS_ADDR_1_sqmuxa_1_0_net_1\, Y => 
        \I5.SENS_ADDR_1_sqmuxa_1_0_adt_net_855880__net_1\);
    
    \I3.VDBOFFB_30_IV_0L0R_2487\ : AO21
      port map(A => \REGl333r\, B => \I3.REGMAPl39r_net_1\, C => 
        \I3.VDBoffb_30l0r_adt_net_163098_\, Y => 
        \I3.VDBoffb_30l0r_adt_net_163124_\);
    
    \I3.PIPEA1l29r\ : DFFS
      port map(CLK => CLK_c, D => \I3.PIPEA1_327_net_1\, SET => 
        CLEAR_STAT_i_0, Q => \I3.PIPEA1l29r_net_1\);
    
    \I3.VDBOFFA_31_IV_0L0R_2624\ : AND2
      port map(A => \REGl165r\, B => \I3.REGMAPl18r_net_1\, Y => 
        \I3.VDBoffa_31l0r_adt_net_164618_\);
    
    \I3.VDBI_57_IV_0_0L6R_2233\ : AND2
      port map(A => \I3.STATE1_ipl0r_adt_net_854360__net_1\, B
         => \I3.VDBoffl6r_net_1\, Y => 
        \I3.VDBi_57l6r_adt_net_143384_\);
    
    \I2.BNCID_VECTror_adt_net_48231_\ : AO21
      port map(A => \I2.BNCID_VECTra12_1_net_1\, B => 
        \I2.BNCID_VECTro_0\, C => 
        \I2.BNCID_VECTror_adt_net_48223__net_1\, Y => 
        \I2.BNCID_VECTror_adt_net_48231__net_1\);
    
    \I2.PIPE4_DT_I_IL1R_2957\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE3_DTl1r_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.PIPE4_DT_I_IL1R_474\);
    
    \I2.PIPE2_DTl27r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl27r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl27r_net_1\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I91_Y\ : AO21FTT
      port map(A => \I2.N303_0\, B => \I2.N306_i_i\, C => 
        \I2.N302_0\, Y => \I2.N345\);
    
    \I2.N_2838_i_0_a2_0_a2_0_a2\ : NAND2FT
      port map(A => 
        \I2.DTO_16_1_iv_0_a2_2_0l21r_adt_net_1014__adt_net_854996__net_1\, 
        B => \I2.N_4184\, Y => \I2.N_2838_i_0\);
    
    \I1.REG_1_99\ : MUX2H
      port map(A => \REGl198r\, B => \I1.N_1337\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855412__net_1\, Y => 
        \I1.REG_1_99_net_1\);
    
    \I1.REG_1_175\ : MUX2H
      port map(A => \REGl274r\, B => \I1.REG_74l274r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y => 
        \I1.REG_1_175_net_1\);
    
    LED_G_pad : OB33PH
      port map(PAD => LED_G, A => LED_G_c);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I153_Y_I_O4_1554\ : AO21
      port map(A => \I2.PIPE4_DTl15r_net_1\, B => 
        \I2.PIPE4_DTL13R_642\, C => \I2.RAMDT4L5R_819\, Y => 
        \I2.N_33_adt_net_55020_\);
    
    \I3.VDBI_57_0_IVL17R_2180\ : AO21
      port map(A => \I3.VDBil17r_net_1\, B => 
        \I3.N_1910_0_adt_net_854336__net_1\, C => 
        \I3.VDBi_57l17r_adt_net_139627_\, Y => 
        \I3.VDBi_57l17r_adt_net_139631_\);
    
    \I2.L2TYPE_4_IL13R_1619\ : AND2
      port map(A => \I2.L2TYPE_i_0_il13r\, B => 
        \I2.N_4439_adt_net_67071_\, Y => 
        \I2.N_4439_adt_net_67114_\);
    
    \I2.WPAGEl12r\ : DFFC
      port map(CLK => CLK_c, D => \I2.WPAGE_951_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.WPAGEl12r_net_1\);
    
    \I3.STATE1_ipl3r_adt_net_854364_\ : BFR
      port map(A => \I3.STATE1_ipl3r_adt_net_854368__net_1\, Y
         => \I3.STATE1_ipl3r_adt_net_854364__net_1\);
    
    \I3.STATE1_ipl0r_adt_net_854360_\ : BFR
      port map(A => \I3.STATE1_ipl0r_net_1\, Y => 
        \I3.STATE1_ipl0r_adt_net_854360__net_1\);
    
    \I2.SUB9l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.SUB9_568_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.SUB9l0r_net_1\);
    
    \I2.SUB8_520_2703\ : NOR3FTT
      port map(A => \I2.SUB8_1_sqmuxa_0_adt_net_855136__net_1\, B
         => \I2.SUB_21x21_fast_I213_Y_0\, C => \I2.N298_0\, Y => 
        \I2.SUB8_520_adt_net_531407_\);
    
    \I2.UN27_PIPE5_DT_1_ADD_21X21_FAST_I138_Y_0_1582\ : OA21FTF
      port map(A => \I2.N_20_i_0\, B => \I2.N_70_0\, C => 
        \I2.ADD_21x21_fast_I138_Y_0_0_0\, Y => 
        \I2.N513_i_0_adt_net_58712_\);
    
    \I1.LUT_3006\ : DFFC
      port map(CLK => CLK_c, D => \I1.LUT_55_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \I1.LUT_760\);
    
    \I2.END_EVNT5_1144\ : DFFC
      port map(CLK => CLK_c, D => \I2.END_EVNT4_net_1\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.END_EVNT5_406\);
    
    \I1.REG_16_sqmuxa_0_a2_m3_e_2\ : AND3FFT
      port map(A => \I1.UN110_BITCNT_7_0_A2_0_A3_0_A2_1_RD1__458\, 
        B => \PULSEl0r\, C => \I1.REG_74_2_0l404r_Rd1__net_1\, Y
         => \I1.REG_74_1_i_a2_a0_2l404r\);
    
    \I2.PIPE10_DT_621\ : MUX2L
      port map(A => \I2.PIPE10_DTl16r_net_1\, B => \I2.N_3802\, S
         => \I2.NWPIPE9_0_net_1\, Y => \I2.PIPE10_DT_621_net_1\);
    
    \I2.MIC_ERR_REGS_356\ : MUX2L
      port map(A => \I2.MIC_ERR_REGSl28r_net_1\, B => 
        \I2.MIC_ERR_REGSl27r_net_1\, S => 
        \I2.MIC_REG1_1_sqmuxa_0_adt_net_855852__net_1\, Y => 
        \I2.MIC_ERR_REGS_356_net_1\);
    
    \I3.UN12_TCNT3_2642\ : AND3FFT
      port map(A => \I3.TCNT3_i_0_il2r_net_1\, B => 
        \I3.TCNT3l1r_net_1\, C => \I3.un12_tcnt3_adt_net_165616_\, 
        Y => \I3.un12_tcnt3_adt_net_165620_\);
    
    \I3.un1_STATE2_13_adt_net_150833_\ : AND3FFT
      port map(A => \I3.N_203\, B => DTEST_FIFO, C => 
        \I3.STATE2l4r_net_1\, Y => 
        \I3.un1_STATE2_13_adt_net_150833__net_1\);
    
    \I2.END_EVNT1_1_sqmuxa_1_0_o2_0\ : NOR3
      port map(A => \I2.N_3280\, B => \I2.STATE1l14r_net_1\, C
         => \I2.STATE1l4r_net_1\, Y => \I2.N_3279_0\);
    
    \I2.CRC32_12_i_m2l0r\ : MUX2L
      port map(A => \I2.DT_TEMPl0r_net_1\, B => 
        \I2.DT_SRAMl0r_net_1\, S => 
        \I2.N_4667_1_adt_net_1046__adt_net_854188__net_1\, Y => 
        \I2.N_3954_i_i\);
    
    \I1.REG_1_177\ : MUX2H
      port map(A => \REGl276r\, B => \I1.REG_74l276r_net_1\, S
         => \I1.N_50_0_adt_net_1409__adt_net_855448__net_1\, Y
         => \I1.REG_1_177_net_1\);
    
    \I2.STATE1l3r\ : DFFC
      port map(CLK => \I2.CLK_tdc\, D => \I2.N_154\, CLR => 
        CLEAR_STAT_i_0, Q => \I2.STATE1l3r_net_1\);
    
    \I2.RAMDT4L12R_2817\ : DFFC
      port map(CLK => CLK_c, D => RAMDT_inl12r, CLR => 
        CLEAR_STAT_i_0, Q => \I2.RAMDT4L12R_145\);
    
    \I2.SUB8_516\ : MUX2H
      port map(A => \I2.SUB8l13r_adt_net_855564__net_1\, B => 
        \I2.SUB8_2l13r\, S => 
        \I2.SUB8_1_sqmuxa_0_adt_net_855140__net_1\, Y => 
        \I2.SUB8_516_net_1\);
    
    \I2.MIC_ERR_REGSl0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_ERR_REGS_329_net_1\, 
        CLR => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_ERR_REGSl0r_net_1\);
    
    \I2.PIPE2_DTl23r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE1_DTl23r_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE2_DTl23r_net_1\);
    
    \I2.RAMAD1_12l5r\ : MUX2L
      port map(A => \I2.TDCDASl3r_net_1\, B => 
        \I2.TDCDBSl3r_net_1\, S => 
        \I2.STATE1l12r_adt_net_855180__net_1\, Y => 
        \I2.RAMAD1_12l5r_net_1\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I176_Y_0\ : XOR2
      port map(A => \I2.RAMDT4L5R_139\, B => 
        \I2.PIPE4_DTl6r_net_1\, Y => \I2.ADD_21x21_fast_I176_Y_0\);
    
    \I2.un27_pipe5_dt_0_ADD_21x21_fast_I16_P0N_i_o2\ : OR2
      port map(A => \I2.RAMDT4L5R_139\, B => 
        \I2.PIPE4_DTl16r_net_1\, Y => \I2.N_65\);
    
    \I5.AIR_PULSE_3\ : MUX2L
      port map(A => \I5.AIR_PULSE_net_1\, B => \I5.N_459\, S => 
        \I5.un1_sstate2_3_0_net_1\, Y => \I5.AIR_PULSE_3_net_1\);
    
    \I2.MIC_REG3l0r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_317_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l0r_net_1\);
    
    \I3.REGMAPL29R_3017\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un126_reg_ads_0_a2_1_a3_net_1\, Q => 
        \I3.REGMAPL29R_771\);
    
    \I2.LEAD_FLAG6_0_sqmuxa_1_0_a4_0_a2_1\ : NOR2
      port map(A => END_FLUSH_559, B => \I2.LEAD_FLAG6_0_sqmuxa\, 
        Y => \I2.LEAD_FLAG6_0_sqmuxa_1_1\);
    
    \I2.FIRST_TDC_1_sqmuxa_1_0\ : OR2FT
      port map(A => \I2.STATE1L12R_647\, B => 
        \I2.END_CHAINA1_1_sqmuxa_3\, Y => 
        \I2.NWPIPE1_4_sqmuxa_1_0\);
    
    \I2.OFFSET_37_9l3r\ : MUX2L
      port map(A => \REGl392r\, B => \REGl328r\, S => 
        \I2.PIPE7_DTL27R_81\, Y => \I2.N_702\);
    
    \I3.VDBI_57_IV_0_0_O2_0_7L0R_2283\ : OR3
      port map(A => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146447_\, B => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146448_\, C => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146432_\, Y => 
        \I3.VDBi_57_iv_0_0_o2_0_7_il0r_adt_net_146451_\);
    
    \I2.SUB8_2_0_0_SUB_21x21_fast_I55_Y\ : AND2
      port map(A => \I2.N267_0\, B => \I2.N270_0\, Y => 
        \I2.N305_0\);
    
    \I3.VDBI_57_IV_0_0L2R_2263\ : AO21
      port map(A => \I3.PIPEAl2r_net_1\, B => \I3.N_90_i_0\, C
         => \I3.VDBi_57l2r_adt_net_145362_\, Y => 
        \I3.VDBi_57l2r_adt_net_145379_\);
    
    \I2.ADE_4l4r\ : MUX2H
      port map(A => \I2.WOFFSETl5r\, B => \I2.ROFFSETl5r_net_1\, 
        S => NOESRAME_c, Y => \I2.ADE_4l4r_net_1\);
    
    \I2.un27_pipe5_dt_1_ADD_21x21_fast_I153_Y_i_a4_0\ : NAND3FFT
      port map(A => \I2.N_152_i_0_adt_net_4117__net_1\, B => 
        \I2.N519_0\, C => \I2.N_163_0\, Y => \I2.N_86_i_0\);
    
    \I1.REG_74l196r\ : OR2
      port map(A => \I1.REG_3_sqmuxa\, B => 
        \I1.N_65_adt_net_1433__net_1\, Y => \I1.N_65\);
    
    DPR_padl18r : IB33
      port map(PAD => DPR(18), Y => DPR_cl18r);
    
    \I1.REG_74_24_404_m3_e\ : OR2
      port map(A => \I1.PAGECNT_0l7r_adt_net_835112_Rd1__net_1\, 
        B => \I1.REG_74_1_a0_0l228r_adt_net_854832__net_1\, Y => 
        \I1.REG_74_24_404_m3_e_net_1\);
    
    REGl295r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_196_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl295r\);
    
    \I2.PIPE9_DTl31r\ : DFFC
      port map(CLK => CLK_c, D => \I2.PIPE9_DT_300_net_1\, CLR
         => CLEAR_STAT_i_0, Q => \I2.PIPE9_DTl31r_net_1\);
    
    \I1.REG_74_0_IVL382R_1811\ : AND2
      port map(A => \FBOUTl1r\, B => \I1.REG_28_sqmuxa\, Y => 
        \I1.REG_74l382r_adt_net_111835_\);
    
    REGl298r : DFFC
      port map(CLK => CLK_c, D => \I1.REG_1_199_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => \REGl298r\);
    
    \I2.REG_1_c13_i\ : AOI21FTT
      port map(A => \I2.un8_evread_1_adt_net_855796__net_1\, B
         => \I2.N_3859\, C => \I2.N_138\, Y => \I2.N_3842_i_0\);
    
    \I2.TRGSERV_2_I_21\ : AND2
      port map(A => \I2.DWACT_ADD_CI_0_g_array_1_0l0r\, B => 
        \I2.TRGSERVl2r_net_1\, Y => 
        \I2.DWACT_ADD_CI_0_g_array_12_0l0r\);
    
    \I2.un1_STATE1_40_1_adt_net_812__adt_net_854572_\ : BFR
      port map(A => \I2.un1_STATE1_40_1_adt_net_812__net_1\, Y
         => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854572__net_1\);
    
    \I2.MIC_REG3l3r\ : DFFC
      port map(CLK => CLK_c, D => \I2.MIC_REG3_320_net_1\, CLR
         => \HWRES_3_adt_net_738__net_1\, Q => 
        \I2.MIC_REG3l3r_net_1\);
    
    \I1.PAGECNTl9r_adt_net_854816_\ : BFR
      port map(A => \I1.PAGECNTL9R_246\, Y => 
        \I1.PAGECNTl9r_adt_net_854816__net_1\);
    
    VDB_pad_il31r : OAI21FTT
      port map(A => \I3.N_290\, B => \I3.LWORDS_net_1\, C => 
        NOEAD_c, Y => NOE32R_c_i_0);
    
    \I3.N_243_4_adt_net_1290__adt_net_854476_\ : BFR
      port map(A => 
        \I3.N_243_4_adt_net_1290__adt_net_854492__net_1\, Y => 
        \I3.N_243_4_adt_net_1290__adt_net_854476__net_1\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I151_Y_I_A4_0_1552\ : OA21
      port map(A => \I2.N_152_i_adt_net_54886_\, B => 
        \I2.N_152_i_adt_net_54890_\, C => \I2.N_20_i\, Y => 
        \I2.N_41_adt_net_54984_\);
    
    \I2.UN27_PIPE5_DT_0_ADD_21X21_FAST_I142_Y_0_A2_1_2667\ : OR2
      port map(A => \I2.N_107_adt_net_276024_\, B => \I2.N_28\, Y
         => \I2.N_107_adt_net_256839_\);
    
    \I2.PIPE8_DT_21_e_0l4r\ : NAND2FT
      port map(A => \I2.NWPIPE7_689\, B => 
        \I2.N_587_adt_net_1201__adt_net_855168__net_1\, Y => 
        \I2.N_4707_i_0\);
    
    \I3.REGMAPl14r\ : DFF
      port map(CLK => CLK_c, D => 
        \I3.un57_reg_ads_0_a2_3_a3_net_1\, Q => 
        \I3.REGMAPl14r_net_1\);
    
    \I2.PIPE1_DT_750\ : MUX2L
      port map(A => \I2.PIPE1_DTl23r_net_1\, B => 
        \I2.PIPE1_DT_42l23r\, S => 
        \I2.un1_STATE1_40_1_adt_net_812__adt_net_854568__net_1\, 
        Y => \I2.PIPE1_DT_750_net_1\);
    
    \I2.TDCDBSl31r_1241\ : DFF
      port map(CLK => \I2.CLK_tdc\, D => TDCDB_cl31r, Q => 
        \I2.TDCDBSL31R_503\);
    
    \I2.L2TYPE_4_IL6R_1630\ : NAND2
      port map(A => \I2.N_4456\, B => \I2.N_4460\, Y => 
        \I2.N_4446_adt_net_67934_\);
    
    \I3.TCNT2_i_0_il4r\ : DFFC
      port map(CLK => CLK_c, D => \I3.TCNT2_392_net_1\, CLR => 
        \HWRES_3_adt_net_738__net_1\, Q => 
        \I3.TCNT2_i_0_il4r_net_1\);
    
    \I3.PIPEA1_323\ : MUX2L
      port map(A => \I3.PIPEA1l25r_net_1\, B => 
        \I3.PIPEA1_12l25r_net_1\, S => 
        \I3.UN1_STATE2_15_1_ADT_NET_1342__250\, Y => 
        \I3.PIPEA1_323_net_1\);
    
    \I3.VDBi_29l9r_adt_net_1596_\ : AO21FTT
      port map(A => LOAD_RES_1, B => \I3.N_2040_261\, C => 
        \I3.VDBi_29l9r_adt_net_142020__net_1\, Y => 
        \I3.VDBi_29l9r_adt_net_1596__net_1\);
    
    \I2.DT_SRAMl14r\ : MUX2L
      port map(A => \I2.N_882\, B => \I2.PIPE2_DTl14r_net_1\, S
         => \I2.N_4646_1_adt_net_1645_Rd1__adt_net_855672__net_1\, 
        Y => \I2.DT_SRAMl14r_net_1\);
    
    \I1.REG_1_184\ : MUX2H
      port map(A => \REGl283r\, B => \I1.REG_74l283r\, S => 
        \I1.N_50_0_adt_net_1409__adt_net_855472__net_1\, Y => 
        \I1.REG_1_184_net_1\);
    

end DEF_ARCH; 
