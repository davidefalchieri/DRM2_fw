----------------------------------------------------------------------------------
-- Company		: OCST Co.,Ltd.
-- Engineer		: RyuShinHyung
-- 
-- Create Date	: 02/23/2005
-- Design Name	: 
-- Module Name	: DEC8B10B - RTL
-- Project Name	: Fiber Optic Application
--
-- Revision
-- Revision 0.01 - File Created
--          1.00 - publishing on the opencores.org
--          1.01 - eliminate needing the VECTLIB.vhd in the original revision.(20110424)
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEC8B10B is
	port
	(
		CLK_IN : IN STD_LOGIC;
		ENCODE_IN : in STD_LOGIC_VECTOR(9 downto 0);
		CTRL_OUT : out STD_LOGIC;
		DATA_OUT : out STD_LOGIC_VECTOR(7 downto 0)
	);
end DEC8B10B;

architecture RTL of DEC8B10B is

constant DEC8b10bERR : std_logic_vector := "100000000";
type TYPE_DEC8b10b is array (0 to 1023) of std_logic_vector (8 downto 0); -- Ctrl & Value
signal TBL_DEC8b10b : TYPE_DEC8b10b:=
	(
		DEC8b10bERR,	-- "0000000000" 
		DEC8b10bERR,	-- "0000000001" 
		DEC8b10bERR,	-- "0000000010" 
		DEC8b10bERR,	-- "0000000011" 
		DEC8b10bERR,	-- "0000000100" 
		DEC8b10bERR,	-- "0000000101" 
		DEC8b10bERR,	-- "0000000110" 
		DEC8b10bERR,	-- "0000000111" 
		DEC8b10bERR,	-- "0000001000" 
		DEC8b10bERR,	-- "0000001001" 
		DEC8b10bERR,	-- "0000001010" 
		DEC8b10bERR,	-- "0000001011" 
		DEC8b10bERR,	-- "0000001100" 
		DEC8b10bERR,	-- "0000001101" 
		DEC8b10bERR,	-- "0000001110" 
		DEC8b10bERR,	-- "0000001111" 
		DEC8b10bERR,	-- "0000010000" 
		DEC8b10bERR,	-- "0000010001" 
		DEC8b10bERR,	-- "0000010010" 
		DEC8b10bERR,	-- "0000010011" 
		DEC8b10bERR,	-- "0000010100" 
		DEC8b10bERR,	-- "0000010101" 
		DEC8b10bERR,	-- "0000010110" 
		DEC8b10bERR,	-- "0000010111" 
		DEC8b10bERR,	-- "0000011000" 
		DEC8b10bERR,	-- "0000011001" 
		DEC8b10bERR,	-- "0000011010" 
		DEC8b10bERR,	-- "0000011011" 
		DEC8b10bERR,	-- "0000011100" 
		DEC8b10bERR,	-- "0000011101" 
		DEC8b10bERR,	-- "0000011110" 
		DEC8b10bERR,	-- "0000011111" 
		DEC8b10bERR,	-- "0000100000" 
		DEC8b10bERR,	-- "0000100001" 
		DEC8b10bERR,	-- "0000100010" 
		DEC8b10bERR,	-- "0000100011" 
		DEC8b10bERR,	-- "0000100100" 
		DEC8b10bERR,	-- "0000100101" 
		DEC8b10bERR,	-- "0000100110" 
		DEC8b10bERR,	-- "0000100111" 
		DEC8b10bERR,	-- "0000101000" 
		DEC8b10bERR,	-- "0000101001" 
		DEC8b10bERR,	-- "0000101010" 
		DEC8b10bERR,	-- "0000101011" 
		DEC8b10bERR,	-- "0000101100" 
		DEC8b10bERR,	-- "0000101101" 
		DEC8b10bERR,	-- "0000101110" 
		DEC8b10bERR,	-- "0000101111" 
		DEC8b10bERR,	-- "0000110000" 
		DEC8b10bERR,	-- "0000110001" 
		DEC8b10bERR,	-- "0000110010" 
		DEC8b10bERR,	-- "0000110011" 
		DEC8b10bERR,	-- "0000110100" 
		DEC8b10bERR,	-- "0000110101" 
		DEC8b10bERR,	-- "0000110110" 
		DEC8b10bERR,	-- "0000110111" 
		DEC8b10bERR,	-- "0000111000" 
		DEC8b10bERR,	-- "0000111001" 
		DEC8b10bERR,	-- "0000111010" 
		DEC8b10bERR,	-- "0000111011" 
		DEC8b10bERR,	-- "0000111100" 
		DEC8b10bERR,	-- "0000111101" 
		DEC8b10bERR,	-- "0000111110" 
		DEC8b10bERR,	-- "0000111111" 
		DEC8b10bERR,	-- "0001000000" 
		DEC8b10bERR,	-- "0001000001" 
		DEC8b10bERR,	-- "0001000010" 
		DEC8b10bERR,	-- "0001000011" 
		DEC8b10bERR,	-- "0001000100" 
		DEC8b10bERR,	-- "0001000101" 
		DEC8b10bERR,	-- "0001000110" 
		DEC8b10bERR,	-- "0001000111" 
		DEC8b10bERR,	-- "0001001000" 
		DEC8b10bERR,	-- "0001001001" 
		DEC8b10bERR,	-- "0001001010" 
		"011101011",	-- "0001001011", -D11.7+, [1,1]
		DEC8b10bERR,	-- "0001001100" 
		"011101101",	-- "0001001101", -D13.7+, [2,2]
		"011101110",	-- "0001001110", -D14.7+, [3,3]
		DEC8b10bERR,	-- "0001001111" 
		DEC8b10bERR,	-- "0001010000" 
		DEC8b10bERR,	-- "0001010001" 
		DEC8b10bERR,	-- "0001010010" 
		"111110011",	-- "0001010011", -K19.7+, [4,1]
		DEC8b10bERR,	-- "0001010100" 
		"111110101",	-- "0001010101", -K21.7+, [5,2]
		"111110110",	-- "0001010110", -K22.7+, [6,3]
		"111110111",	-- "0001010111", +K23.7+, [7,4]
		DEC8b10bERR,	-- "0001011000" 
		"111111001",	-- "0001011001", -K25.7+, [8,5]
		"111111010",	-- "0001011010", -K26.7+, [9,6]
		"111111011",	-- "0001011011", +K27.7+, [10,7]
		DEC8b10bERR,	-- "0001011100" 
		"111111101",	-- "0001011101", +K29.7+, [11,8]
		"111111110",	-- "0001011110", +K30.7+, [12,9]
		DEC8b10bERR,	-- "0001011111" 
		DEC8b10bERR,	-- "0001100000" 
		DEC8b10bERR,	-- "0001100001" 
		DEC8b10bERR,	-- "0001100010" 
		"111100011",	-- "0001100011", -K3.7+, [13,10]
		DEC8b10bERR,	-- "0001100100" 
		"111100101",	-- "0001100101", -K5.7+, [14,11]
		"111100110",	-- "0001100110", -K6.7+, [15,12]
		"111101000",	-- "0001100111", +K8.7+, [16,13]
		DEC8b10bERR,	-- "0001101000" 
		"111101001",	-- "0001101001", -K9.7+, [17,14]
		"111101010",	-- "0001101010", -K10.7+, [18,15]
		"111100100",	-- "0001101011", +K4.7+, [19,16]
		"111101100",	-- "0001101100", -K12.7+, [20,17]
		"111100010",	-- "0001101101", +K2.7+, [21,18]
		"111100001",	-- "0001101110", +K1.7+, [22,19]
		DEC8b10bERR,	-- "0001101111" 
		DEC8b10bERR,	-- "0001110000" 
		"111110001",	-- "0001110001", -K17.7+, [23,20]
		"111110010",	-- "0001110010", -K18.7+, [24,21]
		"111111000",	-- "0001110011", +K24.7+, [25,22]
		"111110100",	-- "0001110100", -K20.7+, [26,23]
		"111111111",	-- "0001110101", +K31.7+, [27,24]
		"111110000",	-- "0001110110", +K16.7+, [28,25]
		DEC8b10bERR,	-- "0001110111" 
		"111100111",	-- "0001111000", -K7.7+, [29,26]
		"111100000",	-- "0001111001", +K0.7+, [30,27]
		"111101111",	-- "0001111010", +K15.7+, [31,28]
		DEC8b10bERR,	-- "0001111011" 
		"111111100",	-- "0001111100", +K28.7+, [32,29]
		DEC8b10bERR,	-- "0001111101" 
		DEC8b10bERR,	-- "0001111110" 
		DEC8b10bERR,	-- "0001111111" 
		DEC8b10bERR,	-- "0010000000" 
		DEC8b10bERR,	-- "0010000001" 
		DEC8b10bERR,	-- "0010000010" 
		DEC8b10bERR,	-- "0010000011" 
		DEC8b10bERR,	-- "0010000100" 
		DEC8b10bERR,	-- "0010000101" 
		DEC8b10bERR,	-- "0010000110" 
		DEC8b10bERR,	-- "0010000111" 
		DEC8b10bERR,	-- "0010001000" 
		DEC8b10bERR,	-- "0010001001" 
		DEC8b10bERR,	-- "0010001010" 
		"000001011",	-- "0010001011", -D11.0+, [33,4]
		DEC8b10bERR,	-- "0010001100" 
		"000001101",	-- "0010001101", -D13.0+, [34,5]
		"000001110",	-- "0010001110", -D14.0+, [35,6]
		DEC8b10bERR,	-- "0010001111" 
		DEC8b10bERR,	-- "0010010000" 
		DEC8b10bERR,	-- "0010010001" 
		DEC8b10bERR,	-- "0010010010" 
		"000010011",	-- "0010010011", -D19.0+, [36,7]
		DEC8b10bERR,	-- "0010010100" 
		"000010101",	-- "0010010101", -D21.0+, [37,8]
		"000010110",	-- "0010010110", -D22.0+, [38,9]
		"000010111",	-- "0010010111", +D23.0+, [39,10]
		DEC8b10bERR,	-- "0010011000" 
		"000011001",	-- "0010011001", -D25.0+, [40,11]
		"000011010",	-- "0010011010", -D26.0+, [41,12]
		"000011011",	-- "0010011011", +D27.0+, [42,13]
		"000011100",	-- "0010011100", -D28.0+, [43,14]
		"000011101",	-- "0010011101", +D29.0+, [44,15]
		"000011110",	-- "0010011110", +D30.0+, [45,16]
		DEC8b10bERR,	-- "0010011111" 
		DEC8b10bERR,	-- "0010100000" 
		DEC8b10bERR,	-- "0010100001" 
		DEC8b10bERR,	-- "0010100010" 
		"000000011",	-- "0010100011", -D3.0+, [46,17]
		DEC8b10bERR,	-- "0010100100" 
		"000000101",	-- "0010100101", -D5.0+, [47,18]
		"000000110",	-- "0010100110", -D6.0+, [48,19]
		"000001000",	-- "0010100111", +D8.0+, [49,20]
		DEC8b10bERR,	-- "0010101000" 
		"000001001",	-- "0010101001", -D9.0+, [50,21]
		"000001010",	-- "0010101010", -D10.0+, [51,22]
		"000000100",	-- "0010101011", +D4.0+, [52,23]
		"000001100",	-- "0010101100", -D12.0+, [53,24]
		"000000010",	-- "0010101101", +D2.0+, [54,25]
		"000000001",	-- "0010101110", +D1.0+, [55,26]
		DEC8b10bERR,	-- "0010101111" 
		DEC8b10bERR,	-- "0010110000" 
		"000010001",	-- "0010110001", -D17.0+, [56,27]
		"000010010",	-- "0010110010", -D18.0+, [57,28]
		"000011000",	-- "0010110011", +D24.0+, [58,29]
		"000010100",	-- "0010110100", -D20.0+, [59,30]
		"000011111",	-- "0010110101", +D31.0+, [60,31]
		"000010000",	-- "0010110110", +D16.0+, [61,32]
		DEC8b10bERR,	-- "0010110111" 
		"000000111",	-- "0010111000", -D7.0+, [62,33]
		"000000000",	-- "0010111001", +D0.0+, [63,34]
		"000001111",	-- "0010111010", +D15.0+, [64,35]
		DEC8b10bERR,	-- "0010111011" 
		"100011100",	-- "0010111100", +K28.0+, [65,30]
		DEC8b10bERR,	-- "0010111101" 
		DEC8b10bERR,	-- "0010111110" 
		DEC8b10bERR,	-- "0010111111" 
		DEC8b10bERR,	-- "0011000000" 
		DEC8b10bERR,	-- "0011000001" 
		DEC8b10bERR,	-- "0011000010" 
		"101111100",	-- "0011000011", -K28.3+, [66,31]
		DEC8b10bERR,	-- "0011000100" 
		"001101111",	-- "0011000101", -D15.3+, [67,36]
		"001100000",	-- "0011000110", -D0.3+, [68,37]
		"001100111",	-- "0011000111", +D7.3+, [69,38]
		DEC8b10bERR,	-- "0011001000" 
		"001110000",	-- "0011001001", -D16.3+, [70,39]
		"001111111",	-- "0011001010", -D31.3+, [71,40]
		"001101011",	-- "0011001011", +D11.3+, [72,41]
		"001111000",	-- "0011001100", -D24.3+, [73,42]
		"001101101",	-- "0011001101", +D13.3+, [74,43]
		"001101110",	-- "0011001110", +D14.3+, [75,44]
		DEC8b10bERR,	-- "0011001111" 
		DEC8b10bERR,	-- "0011010000" 
		"001100001",	-- "0011010001", -D1.3+, [76,45]
		"001100010",	-- "0011010010", -D2.3+, [77,46]
		"001110011",	-- "0011010011", +D19.3+, [78,47]
		"001100100",	-- "0011010100", -D4.3+, [79,48]
		"001110101",	-- "0011010101", +D21.3+, [80,49]
		"001110110",	-- "0011010110", +D22.3+, [81,50]
		DEC8b10bERR,	-- "0011010111" 
		"001101000",	-- "0011011000", -D8.3+, [82,51]
		"001111001",	-- "0011011001", +D25.3+, [83,52]
		"001111010",	-- "0011011010", +D26.3+, [84,53]
		DEC8b10bERR,	-- "0011011011" 
		"001111100",	-- "0011011100", +D28.3+, [85,54]
		DEC8b10bERR,	-- "0011011101" 
		DEC8b10bERR,	-- "0011011110" 
		DEC8b10bERR,	-- "0011011111" 
		DEC8b10bERR,	-- "0011100000" 
		"001111110",	-- "0011100001", -D30.3+, [86,55]
		"001111101",	-- "0011100010", -D29.3+, [87,56]
		"001100011",	-- "0011100011", +D3.3+, [88,57]
		"001111011",	-- "0011100100", -D27.3+, [89,58]
		"001100101",	-- "0011100101", +D5.3+, [90,59]
		"001100110",	-- "0011100110", +D6.3+, [91,60]
		DEC8b10bERR,	-- "0011100111" 
		"001110111",	-- "0011101000", -D23.3+, [92,61]
		"001101001",	-- "0011101001", +D9.3+, [93,62]
		"001101010",	-- "0011101010", +D10.3+, [94,63]
		DEC8b10bERR,	-- "0011101011" 
		"001101100",	-- "0011101100", +D12.3+, [95,64]
		DEC8b10bERR,	-- "0011101101" 
		DEC8b10bERR,	-- "0011101110" 
		DEC8b10bERR,	-- "0011101111" 
		DEC8b10bERR,	-- "0011110000" 
		"001110001",	-- "0011110001", +D17.3+, [96,65]
		"001110010",	-- "0011110010", +D18.3+, [97,66]
		DEC8b10bERR,	-- "0011110011" 
		"001110100",	-- "0011110100", +D20.3+, [98,67]
		DEC8b10bERR,	-- "0011110101" 
		DEC8b10bERR,	-- "0011110110" 
		DEC8b10bERR,	-- "0011110111" 
		DEC8b10bERR,	-- "0011111000" 
		DEC8b10bERR,	-- "0011111001" 
		DEC8b10bERR,	-- "0011111010" 
		DEC8b10bERR,	-- "0011111011" 
		DEC8b10bERR,	-- "0011111100" 
		DEC8b10bERR,	-- "0011111101" 
		DEC8b10bERR,	-- "0011111110" 
		DEC8b10bERR,	-- "0011111111" 
		DEC8b10bERR,	-- "0100000000" 
		DEC8b10bERR,	-- "0100000001" 
		DEC8b10bERR,	-- "0100000010" 
		DEC8b10bERR,	-- "0100000011" 
		DEC8b10bERR,	-- "0100000100" 
		DEC8b10bERR,	-- "0100000101" 
		DEC8b10bERR,	-- "0100000110" 
		DEC8b10bERR,	-- "0100000111" 
		DEC8b10bERR,	-- "0100001000" 
		DEC8b10bERR,	-- "0100001001" 
		DEC8b10bERR,	-- "0100001010" 
		"010001011",	-- "0100001011", -D11.4+, [99,68]
		DEC8b10bERR,	-- "0100001100" 
		"010001101",	-- "0100001101", -D13.4+, [100,69]
		"010001110",	-- "0100001110", -D14.4+, [101,70]
		DEC8b10bERR,	-- "0100001111" 
		DEC8b10bERR,	-- "0100010000" 
		DEC8b10bERR,	-- "0100010001" 
		DEC8b10bERR,	-- "0100010010" 
		"010010011",	-- "0100010011", -D19.4+, [102,71]
		DEC8b10bERR,	-- "0100010100" 
		"010010101",	-- "0100010101", -D21.4+, [103,72]
		"010010110",	-- "0100010110", -D22.4+, [104,73]
		"010010111",	-- "0100010111", +D23.4+, [105,74]
		DEC8b10bERR,	-- "0100011000" 
		"010011001",	-- "0100011001", -D25.4+, [106,75]
		"010011010",	-- "0100011010", -D26.4+, [107,76]
		"010011011",	-- "0100011011", +D27.4+, [108,77]
		"010011100",	-- "0100011100", -D28.4+, [109,78]
		"010011101",	-- "0100011101", +D29.4+, [110,79]
		"010011110",	-- "0100011110", +D30.4+, [111,80]
		DEC8b10bERR,	-- "0100011111" 
		DEC8b10bERR,	-- "0100100000" 
		DEC8b10bERR,	-- "0100100001" 
		DEC8b10bERR,	-- "0100100010" 
		"010000011",	-- "0100100011", -D3.4+, [112,81]
		DEC8b10bERR,	-- "0100100100" 
		"010000101",	-- "0100100101", -D5.4+, [113,82]
		"010000110",	-- "0100100110", -D6.4+, [114,83]
		"010001000",	-- "0100100111", +D8.4+, [115,84]
		DEC8b10bERR,	-- "0100101000" 
		"010001001",	-- "0100101001", -D9.4+, [116,85]
		"010001010",	-- "0100101010", -D10.4+, [117,86]
		"010000100",	-- "0100101011", +D4.4+, [118,87]
		"010001100",	-- "0100101100", -D12.4+, [119,88]
		"010000010",	-- "0100101101", +D2.4+, [120,89]
		"010000001",	-- "0100101110", +D1.4+, [121,90]
		DEC8b10bERR,	-- "0100101111" 
		DEC8b10bERR,	-- "0100110000" 
		"010010001",	-- "0100110001", -D17.4+, [122,91]
		"010010010",	-- "0100110010", -D18.4+, [123,92]
		"010011000",	-- "0100110011", +D24.4+, [124,93]
		"010010100",	-- "0100110100", -D20.4+, [125,94]
		"010011111",	-- "0100110101", +D31.4+, [126,95]
		"010010000",	-- "0100110110", +D16.4+, [127,96]
		DEC8b10bERR,	-- "0100110111" 
		"010000111",	-- "0100111000", -D7.4+, [128,97]
		"010000000",	-- "0100111001", +D0.4+, [129,98]
		"010001111",	-- "0100111010", +D15.4+, [130,99]
		DEC8b10bERR,	-- "0100111011" 
		"110011100",	-- "0100111100", +K28.4+, [131,32]
		DEC8b10bERR,	-- "0100111101" 
		DEC8b10bERR,	-- "0100111110" 
		DEC8b10bERR,	-- "0100111111" 
		DEC8b10bERR,	-- "0101000000" 
		DEC8b10bERR,	-- "0101000001" 
		DEC8b10bERR,	-- "0101000010" 
		"101011100",	-- "0101000011", -K28.2+, [132,33]
		DEC8b10bERR,	-- "0101000100" 
		"010101111",	-- "0101000101", -D15.5+, [133,100]
		"010100000",	-- "0101000110", -D0.5+, [134,101]
		"010100111",	-- "0101000111", +D7.5+, [135,102]
		DEC8b10bERR,	-- "0101001000" 
		"010110000",	-- "0101001001", -D16.5+, [136,103]
		"010111111",	-- "0101001010", -D31.5+, [137,104]
		"010101011",	-- "0101001011", +D11.5+, [138,105]
		"010111000",	-- "0101001100", -D24.5+, [139,106]
		"010101101",	-- "0101001101", +D13.5+, [140,107]
		"010101110",	-- "0101001110", +D14.5+, [141,108]
		DEC8b10bERR,	-- "0101001111" 
		DEC8b10bERR,	-- "0101010000" 
		"010100001",	-- "0101010001", -D1.5+, [142,109]
		"010100010",	-- "0101010010", -D2.5+, [143,110]
		"010110011",	-- "0101010011", +D19.5+, [144,111]
		"010100100",	-- "0101010100", -D4.5+, [145,112]
		"010110101",	-- "0101010101", +D21.5+, [146,113]
		"010110110",	-- "0101010110", +D22.5+, [147,114]
		"010110111",	-- "0101010111", +D23.5-, [148,115]
		"010101000",	-- "0101011000", -D8.5+, [149,116]
		"010111001",	-- "0101011001", +D25.5+, [150,117]
		"010111010",	-- "0101011010", +D26.5+, [151,118]
		"010111011",	-- "0101011011", +D27.5-, [152,119]
		"010111100",	-- "0101011100", +D28.5+, [153,120]
		"010111101",	-- "0101011101", +D29.5-, [154,121]
		"010111110",	-- "0101011110", +D30.5-, [155,122]
		DEC8b10bERR,	-- "0101011111" 
		DEC8b10bERR,	-- "0101100000" 
		"010111110",	-- "0101100001", -D30.5+, [156,123]
		"010111101",	-- "0101100010", -D29.5+, [157,124]
		"010100011",	-- "0101100011", +D3.5+, [158,125]
		"010111011",	-- "0101100100", -D27.5+, [159,126]
		"010100101",	-- "0101100101", +D5.5+, [160,127]
		"010100110",	-- "0101100110", +D6.5+, [161,128]
		"010101000",	-- "0101100111", +D8.5-, [162,129]
		"010110111",	-- "0101101000", -D23.5+, [163,130]
		"010101001",	-- "0101101001", +D9.5+, [164,131]
		"010101010",	-- "0101101010", +D10.5+, [165,132]
		"010100100",	-- "0101101011", +D4.5-, [166,133]
		"010101100",	-- "0101101100", +D12.5+, [167,134]
		"010100010",	-- "0101101101", +D2.5-, [168,135]
		"010100001",	-- "0101101110", +D1.5-, [169,136]
		DEC8b10bERR,	-- "0101101111" 
		DEC8b10bERR,	-- "0101110000" 
		"010110001",	-- "0101110001", +D17.5+, [170,137]
		"010110010",	-- "0101110010", +D18.5+, [171,138]
		"010111000",	-- "0101110011", +D24.5-, [172,139]
		"010110100",	-- "0101110100", +D20.5+, [173,140]
		"010111111",	-- "0101110101", +D31.5-, [174,141]
		"010110000",	-- "0101110110", +D16.5-, [175,142]
		DEC8b10bERR,	-- "0101110111" 
		"010100111",	-- "0101111000", -D7.5-, [176,143]
		"010100000",	-- "0101111001", +D0.5-, [177,144]
		"010101111",	-- "0101111010", +D15.5-, [178,145]
		DEC8b10bERR,	-- "0101111011" 
		"110111100",	-- "0101111100", +K28.5-, [179,34]
		DEC8b10bERR,	-- "0101111101" 
		DEC8b10bERR,	-- "0101111110" 
		DEC8b10bERR,	-- "0101111111" 
		DEC8b10bERR,	-- "0110000000" 
		DEC8b10bERR,	-- "0110000001" 
		DEC8b10bERR,	-- "0110000010" 
		"100111100",	-- "0110000011", -K28.1+, [180,35]
		DEC8b10bERR,	-- "0110000100" 
		"011001111",	-- "0110000101", -D15.6+, [181,146]
		"011000000",	-- "0110000110", -D0.6+, [182,147]
		"011000111",	-- "0110000111", +D7.6+, [183,148]
		DEC8b10bERR,	-- "0110001000" 
		"011010000",	-- "0110001001", -D16.6+, [184,149]
		"011011111",	-- "0110001010", -D31.6+, [185,150]
		"011001011",	-- "0110001011", +D11.6+, [186,151]
		"011011000",	-- "0110001100", -D24.6+, [187,152]
		"011001101",	-- "0110001101", +D13.6+, [188,153]
		"011001110",	-- "0110001110", +D14.6+, [189,154]
		DEC8b10bERR,	-- "0110001111" 
		DEC8b10bERR,	-- "0110010000" 
		"011000001",	-- "0110010001", -D1.6+, [190,155]
		"011000010",	-- "0110010010", -D2.6+, [191,156]
		"011010011",	-- "0110010011", +D19.6+, [192,157]
		"011000100",	-- "0110010100", -D4.6+, [193,158]
		"011010101",	-- "0110010101", +D21.6+, [194,159]
		"011010110",	-- "0110010110", +D22.6+, [195,160]
		"011010111",	-- "0110010111", +D23.6-, [196,161]
		"011001000",	-- "0110011000", -D8.6+, [197,162]
		"011011001",	-- "0110011001", +D25.6+, [198,163]
		"011011010",	-- "0110011010", +D26.6+, [199,164]
		"011011011",	-- "0110011011", +D27.6-, [200,165]
		"011011100",	-- "0110011100", +D28.6+, [201,166]
		"011011101",	-- "0110011101", +D29.6-, [202,167]
		"011011110",	-- "0110011110", +D30.6-, [203,168]
		DEC8b10bERR,	-- "0110011111" 
		DEC8b10bERR,	-- "0110100000" 
		"011011110",	-- "0110100001", -D30.6+, [204,169]
		"011011101",	-- "0110100010", -D29.6+, [205,170]
		"011000011",	-- "0110100011", +D3.6+, [206,171]
		"011011011",	-- "0110100100", -D27.6+, [207,172]
		"011000101",	-- "0110100101", +D5.6+, [208,173]
		"011000110",	-- "0110100110", +D6.6+, [209,174]
		"011001000",	-- "0110100111", +D8.6-, [210,175]
		"011010111",	-- "0110101000", -D23.6+, [211,176]
		"011001001",	-- "0110101001", +D9.6+, [212,177]
		"011001010",	-- "0110101010", +D10.6+, [213,178]
		"011000100",	-- "0110101011", +D4.6-, [214,179]
		"011001100",	-- "0110101100", +D12.6+, [215,180]
		"011000010",	-- "0110101101", +D2.6-, [216,181]
		"011000001",	-- "0110101110", +D1.6-, [217,182]
		DEC8b10bERR,	-- "0110101111" 
		DEC8b10bERR,	-- "0110110000" 
		"011010001",	-- "0110110001", +D17.6+, [218,183]
		"011010010",	-- "0110110010", +D18.6+, [219,184]
		"011011000",	-- "0110110011", +D24.6-, [220,185]
		"011010100",	-- "0110110100", +D20.6+, [221,186]
		"011011111",	-- "0110110101", +D31.6-, [222,187]
		"011010000",	-- "0110110110", +D16.6-, [223,188]
		DEC8b10bERR,	-- "0110110111" 
		"011000111",	-- "0110111000", -D7.6-, [224,189]
		"011000000",	-- "0110111001", +D0.6-, [225,190]
		"011001111",	-- "0110111010", +D15.6-, [226,191]
		DEC8b10bERR,	-- "0110111011" 
		"111011100",	-- "0110111100", +K28.6-, [227,36]
		DEC8b10bERR,	-- "0110111101" 
		DEC8b10bERR,	-- "0110111110" 
		DEC8b10bERR,	-- "0110111111" 
		DEC8b10bERR,	-- "0111000000" 
		DEC8b10bERR,	-- "0111000001" 
		DEC8b10bERR,	-- "0111000010" 
		DEC8b10bERR,	-- "0111000011" 
		DEC8b10bERR,	-- "0111000100" 
		"011101111",	-- "0111000101", -D15.7-, [228,192]
		"011100000",	-- "0111000110", -D0.7-, [229,193]
		"011100111",	-- "0111000111", +D7.7-, [230,194]
		DEC8b10bERR,	-- "0111001000" 
		"011110000",	-- "0111001001", -D16.7-, [231,195]
		"011111111",	-- "0111001010", -D31.7-, [232,196]
		"011101011",	-- "0111001011", +D11.7-, [233,197]
		"011111000",	-- "0111001100", -D24.7-, [234,198]
		"011101101",	-- "0111001101", +D13.7-, [235,199]
		"011101110",	-- "0111001110", +D14.7-, [236,200]
		DEC8b10bERR,	-- "0111001111" 
		DEC8b10bERR,	-- "0111010000" 
		"011100001",	-- "0111010001", -D1.7-, [237,201]
		"011100010",	-- "0111010010", -D2.7-, [238,202]
		"011110011",	-- "0111010011", +D19.7-, [239,203]
		"011100100",	-- "0111010100", -D4.7-, [240,204]
		"011110101",	-- "0111010101", +D21.7-, [241,205]
		"011110110",	-- "0111010110", +D22.7-, [242,206]
		DEC8b10bERR,	-- "0111010111" 
		"011101000",	-- "0111011000", -D8.7-, [243,207]
		"011111001",	-- "0111011001", +D25.7-, [244,208]
		"011111010",	-- "0111011010", +D26.7-, [245,209]
		DEC8b10bERR,	-- "0111011011" 
		"011111100",	-- "0111011100", +D28.7-, [246,210]
		DEC8b10bERR,	-- "0111011101" 
		DEC8b10bERR,	-- "0111011110" 
		DEC8b10bERR,	-- "0111011111" 
		DEC8b10bERR,	-- "0111100000" 
		"011111110",	-- "0111100001", -D30.7-, [247,211]
		"011111101",	-- "0111100010", -D29.7-, [248,212]
		"011100011",	-- "0111100011", +D3.7-, [249,213]
		"011111011",	-- "0111100100", -D27.7-, [250,214]
		"011100101",	-- "0111100101", +D5.7-, [251,215]
		"011100110",	-- "0111100110", +D6.7-, [252,216]
		DEC8b10bERR,	-- "0111100111" 
		"011110111",	-- "0111101000", -D23.7-, [253,217]
		"011101001",	-- "0111101001", +D9.7-, [254,218]
		"011101010",	-- "0111101010", +D10.7-, [255,219]
		DEC8b10bERR,	-- "0111101011" 
		"011101100",	-- "0111101100", +D12.7-, [256,220]
		DEC8b10bERR,	-- "0111101101" 
		DEC8b10bERR,	-- "0111101110" 
		DEC8b10bERR,	-- "0111101111" 
		DEC8b10bERR,	-- "0111110000" 
		DEC8b10bERR,	-- "0111110001" 
		DEC8b10bERR,	-- "0111110010" 
		DEC8b10bERR,	-- "0111110011" 
		DEC8b10bERR,	-- "0111110100" 
		DEC8b10bERR,	-- "0111110101" 
		DEC8b10bERR,	-- "0111110110" 
		DEC8b10bERR,	-- "0111110111" 
		DEC8b10bERR,	-- "0111111000" 
		DEC8b10bERR,	-- "0111111001" 
		DEC8b10bERR,	-- "0111111010" 
		DEC8b10bERR,	-- "0111111011" 
		DEC8b10bERR,	-- "0111111100" 
		DEC8b10bERR,	-- "0111111101" 
		DEC8b10bERR,	-- "0111111110" 
		DEC8b10bERR,	-- "0111111111" 
		DEC8b10bERR,	-- "1000000000" 
		DEC8b10bERR,	-- "1000000001" 
		DEC8b10bERR,	-- "1000000010" 
		DEC8b10bERR,	-- "1000000011" 
		DEC8b10bERR,	-- "1000000100" 
		DEC8b10bERR,	-- "1000000101" 
		DEC8b10bERR,	-- "1000000110" 
		DEC8b10bERR,	-- "1000000111" 
		DEC8b10bERR,	-- "1000001000" 
		DEC8b10bERR,	-- "1000001001" 
		DEC8b10bERR,	-- "1000001010" 
		DEC8b10bERR,	-- "1000001011" 
		DEC8b10bERR,	-- "1000001100" 
		DEC8b10bERR,	-- "1000001101" 
		DEC8b10bERR,	-- "1000001110" 
		DEC8b10bERR,	-- "1000001111" 
		DEC8b10bERR,	-- "1000010000" 
		DEC8b10bERR,	-- "1000010001" 
		DEC8b10bERR,	-- "1000010010" 
		"011110011",	-- "1000010011", -D19.7+, [257,221]
		DEC8b10bERR,	-- "1000010100" 
		"011110101",	-- "1000010101", -D21.7+, [258,222]
		"011110110",	-- "1000010110", -D22.7+, [259,223]
		"011110111",	-- "1000010111", +D23.7+, [260,224]
		DEC8b10bERR,	-- "1000011000" 
		"011111001",	-- "1000011001", -D25.7+, [261,225]
		"011111010",	-- "1000011010", -D26.7+, [262,226]
		"011111011",	-- "1000011011", +D27.7+, [263,227]
		"011111100",	-- "1000011100", -D28.7+, [264,228]
		"011111101",	-- "1000011101", +D29.7+, [265,229]
		"011111110",	-- "1000011110", +D30.7+, [266,230]
		DEC8b10bERR,	-- "1000011111" 
		DEC8b10bERR,	-- "1000100000" 
		DEC8b10bERR,	-- "1000100001" 
		DEC8b10bERR,	-- "1000100010" 
		"011100011",	-- "1000100011", -D3.7+, [267,231]
		DEC8b10bERR,	-- "1000100100" 
		"011100101",	-- "1000100101", -D5.7+, [268,232]
		"011100110",	-- "1000100110", -D6.7+, [269,233]
		"011101000",	-- "1000100111", +D8.7+, [270,234]
		DEC8b10bERR,	-- "1000101000" 
		"011101001",	-- "1000101001", -D9.7+, [271,235]
		"011101010",	-- "1000101010", -D10.7+, [272,236]
		"011100100",	-- "1000101011", +D4.7+, [273,237]
		"011101100",	-- "1000101100", -D12.7+, [274,238]
		"011100010",	-- "1000101101", +D2.7+, [275,239]
		"011100001",	-- "1000101110", +D1.7+, [276,240]
		DEC8b10bERR,	-- "1000101111" 
		DEC8b10bERR,	-- "1000110000" 
		"011110001",	-- "1000110001", -D17.7+, [277,241]
		"011110010",	-- "1000110010", -D18.7+, [278,242]
		"011111000",	-- "1000110011", +D24.7+, [279,243]
		"011110100",	-- "1000110100", -D20.7+, [280,244]
		"011111111",	-- "1000110101", +D31.7+, [281,245]
		"011110000",	-- "1000110110", +D16.7+, [282,246]
		DEC8b10bERR,	-- "1000110111" 
		"011100111",	-- "1000111000", -D7.7+, [283,247]
		"011100000",	-- "1000111001", +D0.7+, [284,248]
		"011101111",	-- "1000111010", +D15.7+, [285,249]
		DEC8b10bERR,	-- "1000111011" 
		DEC8b10bERR,	-- "1000111100" 
		DEC8b10bERR,	-- "1000111101" 
		DEC8b10bERR,	-- "1000111110" 
		DEC8b10bERR,	-- "1000111111" 
		DEC8b10bERR,	-- "1001000000" 
		DEC8b10bERR,	-- "1001000001" 
		DEC8b10bERR,	-- "1001000010" 
		"111011100",	-- "1001000011", -K28.6+, [286,37]
		DEC8b10bERR,	-- "1001000100" 
		"000101111",	-- "1001000101", -D15.1+, [287,250]
		"000100000",	-- "1001000110", -D0.1+, [288,251]
		"000100111",	-- "1001000111", +D7.1+, [289,252]
		DEC8b10bERR,	-- "1001001000" 
		"000110000",	-- "1001001001", -D16.1+, [290,253]
		"000111111",	-- "1001001010", -D31.1+, [291,254]
		"000101011",	-- "1001001011", +D11.1+, [292,255]
		"000111000",	-- "1001001100", -D24.1+, [293,256]
		"000101101",	-- "1001001101", +D13.1+, [294,257]
		"000101110",	-- "1001001110", +D14.1+, [295,258]
		DEC8b10bERR,	-- "1001001111" 
		DEC8b10bERR,	-- "1001010000" 
		"000100001",	-- "1001010001", -D1.1+, [296,259]
		"000100010",	-- "1001010010", -D2.1+, [297,260]
		"000110011",	-- "1001010011", +D19.1+, [298,261]
		"000100100",	-- "1001010100", -D4.1+, [299,262]
		"000110101",	-- "1001010101", +D21.1+, [300,263]
		"000110110",	-- "1001010110", +D22.1+, [301,264]
		"000110111",	-- "1001010111", +D23.1-, [302,265]
		"000101000",	-- "1001011000", -D8.1+, [303,266]
		"000111001",	-- "1001011001", +D25.1+, [304,267]
		"000111010",	-- "1001011010", +D26.1+, [305,268]
		"000111011",	-- "1001011011", +D27.1-, [306,269]
		"000111100",	-- "1001011100", +D28.1+, [307,270]
		"000111101",	-- "1001011101", +D29.1-, [308,271]
		"000111110",	-- "1001011110", +D30.1-, [309,272]
		DEC8b10bERR,	-- "1001011111" 
		DEC8b10bERR,	-- "1001100000" 
		"000111110",	-- "1001100001", -D30.1+, [310,273]
		"000111101",	-- "1001100010", -D29.1+, [311,274]
		"000100011",	-- "1001100011", +D3.1+, [312,275]
		"000111011",	-- "1001100100", -D27.1+, [313,276]
		"000100101",	-- "1001100101", +D5.1+, [314,277]
		"000100110",	-- "1001100110", +D6.1+, [315,278]
		"000101000",	-- "1001100111", +D8.1-, [316,279]
		"000110111",	-- "1001101000", -D23.1+, [317,280]
		"000101001",	-- "1001101001", +D9.1+, [318,281]
		"000101010",	-- "1001101010", +D10.1+, [319,282]
		"000100100",	-- "1001101011", +D4.1-, [320,283]
		"000101100",	-- "1001101100", +D12.1+, [321,284]
		"000100010",	-- "1001101101", +D2.1-, [322,285]
		"000100001",	-- "1001101110", +D1.1-, [323,286]
		DEC8b10bERR,	-- "1001101111" 
		DEC8b10bERR,	-- "1001110000" 
		"000110001",	-- "1001110001", +D17.1+, [324,287]
		"000110010",	-- "1001110010", +D18.1+, [325,288]
		"000111000",	-- "1001110011", +D24.1-, [326,289]
		"000110100",	-- "1001110100", +D20.1+, [327,290]
		"000111111",	-- "1001110101", +D31.1-, [328,291]
		"000110000",	-- "1001110110", +D16.1-, [329,292]
		DEC8b10bERR,	-- "1001110111" 
		"000100111",	-- "1001111000", -D7.1-, [330,293]
		"000100000",	-- "1001111001", +D0.1-, [331,294]
		"000101111",	-- "1001111010", +D15.1-, [332,295]
		DEC8b10bERR,	-- "1001111011" 
		"100111100",	-- "1001111100", +K28.1-, [333,38]
		DEC8b10bERR,	-- "1001111101" 
		DEC8b10bERR,	-- "1001111110" 
		DEC8b10bERR,	-- "1001111111" 
		DEC8b10bERR,	-- "1010000000" 
		DEC8b10bERR,	-- "1010000001" 
		DEC8b10bERR,	-- "1010000010" 
		"110111100",	-- "1010000011", -K28.5+, [334,39]
		DEC8b10bERR,	-- "1010000100" 
		"001001111",	-- "1010000101", -D15.2+, [335,296]
		"001000000",	-- "1010000110", -D0.2+, [336,297]
		"001000111",	-- "1010000111", +D7.2+, [337,298]
		DEC8b10bERR,	-- "1010001000" 
		"001010000",	-- "1010001001", -D16.2+, [338,299]
		"001011111",	-- "1010001010", -D31.2+, [339,300]
		"001001011",	-- "1010001011", +D11.2+, [340,301]
		"001011000",	-- "1010001100", -D24.2+, [341,302]
		"001001101",	-- "1010001101", +D13.2+, [342,303]
		"001001110",	-- "1010001110", +D14.2+, [343,304]
		DEC8b10bERR,	-- "1010001111" 
		DEC8b10bERR,	-- "1010010000" 
		"001000001",	-- "1010010001", -D1.2+, [344,305]
		"001000010",	-- "1010010010", -D2.2+, [345,306]
		"001010011",	-- "1010010011", +D19.2+, [346,307]
		"001000100",	-- "1010010100", -D4.2+, [347,308]
		"001010101",	-- "1010010101", +D21.2+, [348,309]
		"001010110",	-- "1010010110", +D22.2+, [349,310]
		"001010111",	-- "1010010111", +D23.2-, [350,311]
		"001001000",	-- "1010011000", -D8.2+, [351,312]
		"001011001",	-- "1010011001", +D25.2+, [352,313]
		"001011010",	-- "1010011010", +D26.2+, [353,314]
		"001011011",	-- "1010011011", +D27.2-, [354,315]
		"001011100",	-- "1010011100", +D28.2+, [355,316]
		"001011101",	-- "1010011101", +D29.2-, [356,317]
		"001011110",	-- "1010011110", +D30.2-, [357,318]
		DEC8b10bERR,	-- "1010011111" 
		DEC8b10bERR,	-- "1010100000" 
		"001011110",	-- "1010100001", -D30.2+, [358,319]
		"001011101",	-- "1010100010", -D29.2+, [359,320]
		"001000011",	-- "1010100011", +D3.2+, [360,321]
		"001011011",	-- "1010100100", -D27.2+, [361,322]
		"001000101",	-- "1010100101", +D5.2+, [362,323]
		"001000110",	-- "1010100110", +D6.2+, [363,324]
		"001001000",	-- "1010100111", +D8.2-, [364,325]
		"001010111",	-- "1010101000", -D23.2+, [365,326]
		"001001001",	-- "1010101001", +D9.2+, [366,327]
		"001001010",	-- "1010101010", +D10.2+, [367,328]
		"001000100",	-- "1010101011", +D4.2-, [368,329]
		"001001100",	-- "1010101100", +D12.2+, [369,330]
		"001000010",	-- "1010101101", +D2.2-, [370,331]
		"001000001",	-- "1010101110", +D1.2-, [371,332]
		DEC8b10bERR,	-- "1010101111" 
		DEC8b10bERR,	-- "1010110000" 
		"001010001",	-- "1010110001", +D17.2+, [372,333]
		"001010010",	-- "1010110010", +D18.2+, [373,334]
		"001011000",	-- "1010110011", +D24.2-, [374,335]
		"001010100",	-- "1010110100", +D20.2+, [375,336]
		"001011111",	-- "1010110101", +D31.2-, [376,337]
		"001010000",	-- "1010110110", +D16.2-, [377,338]
		DEC8b10bERR,	-- "1010110111" 
		"001000111",	-- "1010111000", -D7.2-, [378,339]
		"001000000",	-- "1010111001", +D0.2-, [379,340]
		"001001111",	-- "1010111010", +D15.2-, [380,341]
		DEC8b10bERR,	-- "1010111011" 
		"101011100",	-- "1010111100", +K28.2-, [381,40]
		DEC8b10bERR,	-- "1010111101" 
		DEC8b10bERR,	-- "1010111110" 
		DEC8b10bERR,	-- "1010111111" 
		DEC8b10bERR,	-- "1011000000" 
		DEC8b10bERR,	-- "1011000001" 
		DEC8b10bERR,	-- "1011000010" 
		"110011100",	-- "1011000011", -K28.4-, [382,41]
		DEC8b10bERR,	-- "1011000100" 
		"010001111",	-- "1011000101", -D15.4-, [383,342]
		"010000000",	-- "1011000110", -D0.4-, [384,343]
		"010000111",	-- "1011000111", +D7.4-, [385,344]
		DEC8b10bERR,	-- "1011001000" 
		"010010000",	-- "1011001001", -D16.4-, [386,345]
		"010011111",	-- "1011001010", -D31.4-, [387,346]
		"010001011",	-- "1011001011", +D11.4-, [388,347]
		"010011000",	-- "1011001100", -D24.4-, [389,348]
		"010001101",	-- "1011001101", +D13.4-, [390,349]
		"010001110",	-- "1011001110", +D14.4-, [391,350]
		DEC8b10bERR,	-- "1011001111" 
		DEC8b10bERR,	-- "1011010000" 
		"010000001",	-- "1011010001", -D1.4-, [392,351]
		"010000010",	-- "1011010010", -D2.4-, [393,352]
		"010010011",	-- "1011010011", +D19.4-, [394,353]
		"010000100",	-- "1011010100", -D4.4-, [395,354]
		"010010101",	-- "1011010101", +D21.4-, [396,355]
		"010010110",	-- "1011010110", +D22.4-, [397,356]
		DEC8b10bERR,	-- "1011010111" 
		"010001000",	-- "1011011000", -D8.4-, [398,357]
		"010011001",	-- "1011011001", +D25.4-, [399,358]
		"010011010",	-- "1011011010", +D26.4-, [400,359]
		DEC8b10bERR,	-- "1011011011" 
		"010011100",	-- "1011011100", +D28.4-, [401,360]
		DEC8b10bERR,	-- "1011011101" 
		DEC8b10bERR,	-- "1011011110" 
		DEC8b10bERR,	-- "1011011111" 
		DEC8b10bERR,	-- "1011100000" 
		"010011110",	-- "1011100001", -D30.4-, [402,361]
		"010011101",	-- "1011100010", -D29.4-, [403,362]
		"010000011",	-- "1011100011", +D3.4-, [404,363]
		"010011011",	-- "1011100100", -D27.4-, [405,364]
		"010000101",	-- "1011100101", +D5.4-, [406,365]
		"010000110",	-- "1011100110", +D6.4-, [407,366]
		DEC8b10bERR,	-- "1011100111" 
		"010010111",	-- "1011101000", -D23.4-, [408,367]
		"010001001",	-- "1011101001", +D9.4-, [409,368]
		"010001010",	-- "1011101010", +D10.4-, [410,369]
		DEC8b10bERR,	-- "1011101011" 
		"010001100",	-- "1011101100", +D12.4-, [411,370]
		DEC8b10bERR,	-- "1011101101" 
		DEC8b10bERR,	-- "1011101110" 
		DEC8b10bERR,	-- "1011101111" 
		DEC8b10bERR,	-- "1011110000" 
		"010010001",	-- "1011110001", +D17.4-, [412,371]
		"010010010",	-- "1011110010", +D18.4-, [413,372]
		DEC8b10bERR,	-- "1011110011" 
		"010010100",	-- "1011110100", +D20.4-, [414,373]
		DEC8b10bERR,	-- "1011110101" 
		DEC8b10bERR,	-- "1011110110" 
		DEC8b10bERR,	-- "1011110111" 
		DEC8b10bERR,	-- "1011111000" 
		DEC8b10bERR,	-- "1011111001" 
		DEC8b10bERR,	-- "1011111010" 
		DEC8b10bERR,	-- "1011111011" 
		DEC8b10bERR,	-- "1011111100" 
		DEC8b10bERR,	-- "1011111101" 
		DEC8b10bERR,	-- "1011111110" 
		DEC8b10bERR,	-- "1011111111" 
		DEC8b10bERR,	-- "1100000000" 
		DEC8b10bERR,	-- "1100000001" 
		DEC8b10bERR,	-- "1100000010" 
		DEC8b10bERR,	-- "1100000011" 
		DEC8b10bERR,	-- "1100000100" 
		DEC8b10bERR,	-- "1100000101" 
		DEC8b10bERR,	-- "1100000110" 
		DEC8b10bERR,	-- "1100000111" 
		DEC8b10bERR,	-- "1100001000" 
		DEC8b10bERR,	-- "1100001001" 
		DEC8b10bERR,	-- "1100001010" 
		"001101011",	-- "1100001011", -D11.3-, [415,374]
		DEC8b10bERR,	-- "1100001100" 
		"001101101",	-- "1100001101", -D13.3-, [416,375]
		"001101110",	-- "1100001110", -D14.3-, [417,376]
		DEC8b10bERR,	-- "1100001111" 
		DEC8b10bERR,	-- "1100010000" 
		DEC8b10bERR,	-- "1100010001" 
		DEC8b10bERR,	-- "1100010010" 
		"001110011",	-- "1100010011", -D19.3-, [418,377]
		DEC8b10bERR,	-- "1100010100" 
		"001110101",	-- "1100010101", -D21.3-, [419,378]
		"001110110",	-- "1100010110", -D22.3-, [420,379]
		"001110111",	-- "1100010111", +D23.3-, [421,380]
		DEC8b10bERR,	-- "1100011000" 
		"001111001",	-- "1100011001", -D25.3-, [422,381]
		"001111010",	-- "1100011010", -D26.3-, [423,382]
		"001111011",	-- "1100011011", +D27.3-, [424,383]
		"001111100",	-- "1100011100", -D28.3-, [425,384]
		"001111101",	-- "1100011101", +D29.3-, [426,385]
		"001111110",	-- "1100011110", +D30.3-, [427,386]
		DEC8b10bERR,	-- "1100011111" 
		DEC8b10bERR,	-- "1100100000" 
		DEC8b10bERR,	-- "1100100001" 
		DEC8b10bERR,	-- "1100100010" 
		"001100011",	-- "1100100011", -D3.3-, [428,387]
		DEC8b10bERR,	-- "1100100100" 
		"001100101",	-- "1100100101", -D5.3-, [429,388]
		"001100110",	-- "1100100110", -D6.3-, [430,389]
		"001101000",	-- "1100100111", +D8.3-, [431,390]
		DEC8b10bERR,	-- "1100101000" 
		"001101001",	-- "1100101001", -D9.3-, [432,391]
		"001101010",	-- "1100101010", -D10.3-, [433,392]
		"001100100",	-- "1100101011", +D4.3-, [434,393]
		"001101100",	-- "1100101100", -D12.3-, [435,394]
		"001100010",	-- "1100101101", +D2.3-, [436,395]
		"001100001",	-- "1100101110", +D1.3-, [437,396]
		DEC8b10bERR,	-- "1100101111" 
		DEC8b10bERR,	-- "1100110000" 
		"001110001",	-- "1100110001", -D17.3-, [438,397]
		"001110010",	-- "1100110010", -D18.3-, [439,398]
		"001111000",	-- "1100110011", +D24.3-, [440,399]
		"001110100",	-- "1100110100", -D20.3-, [441,400]
		"001111111",	-- "1100110101", +D31.3-, [442,401]
		"001110000",	-- "1100110110", +D16.3-, [443,402]
		DEC8b10bERR,	-- "1100110111" 
		"001100111",	-- "1100111000", -D7.3-, [444,403]
		"001100000",	-- "1100111001", +D0.3-, [445,404]
		"001101111",	-- "1100111010", +D15.3-, [446,405]
		DEC8b10bERR,	-- "1100111011" 
		"101111100",	-- "1100111100", +K28.3-, [447,42]
		DEC8b10bERR,	-- "1100111101" 
		DEC8b10bERR,	-- "1100111110" 
		DEC8b10bERR,	-- "1100111111" 
		DEC8b10bERR,	-- "1101000000" 
		DEC8b10bERR,	-- "1101000001" 
		DEC8b10bERR,	-- "1101000010" 
		"100011100",	-- "1101000011", -K28.0-, [448,43]
		DEC8b10bERR,	-- "1101000100" 
		"000001111",	-- "1101000101", -D15.0-, [449,406]
		"000000000",	-- "1101000110", -D0.0-, [450,407]
		"000000111",	-- "1101000111", +D7.0-, [451,408]
		DEC8b10bERR,	-- "1101001000" 
		"000010000",	-- "1101001001", -D16.0-, [452,409]
		"000011111",	-- "1101001010", -D31.0-, [453,410]
		"000001011",	-- "1101001011", +D11.0-, [454,411]
		"000011000",	-- "1101001100", -D24.0-, [455,412]
		"000001101",	-- "1101001101", +D13.0-, [456,413]
		"000001110",	-- "1101001110", +D14.0-, [457,414]
		DEC8b10bERR,	-- "1101001111" 
		DEC8b10bERR,	-- "1101010000" 
		"000000001",	-- "1101010001", -D1.0-, [458,415]
		"000000010",	-- "1101010010", -D2.0-, [459,416]
		"000010011",	-- "1101010011", +D19.0-, [460,417]
		"000000100",	-- "1101010100", -D4.0-, [461,418]
		"000010101",	-- "1101010101", +D21.0-, [462,419]
		"000010110",	-- "1101010110", +D22.0-, [463,420]
		DEC8b10bERR,	-- "1101010111" 
		"000001000",	-- "1101011000", -D8.0-, [464,421]
		"000011001",	-- "1101011001", +D25.0-, [465,422]
		"000011010",	-- "1101011010", +D26.0-, [466,423]
		DEC8b10bERR,	-- "1101011011" 
		"000011100",	-- "1101011100", +D28.0-, [467,424]
		DEC8b10bERR,	-- "1101011101" 
		DEC8b10bERR,	-- "1101011110" 
		DEC8b10bERR,	-- "1101011111" 
		DEC8b10bERR,	-- "1101100000" 
		"000011110",	-- "1101100001", -D30.0-, [468,425]
		"000011101",	-- "1101100010", -D29.0-, [469,426]
		"000000011",	-- "1101100011", +D3.0-, [470,427]
		"000011011",	-- "1101100100", -D27.0-, [471,428]
		"000000101",	-- "1101100101", +D5.0-, [472,429]
		"000000110",	-- "1101100110", +D6.0-, [473,430]
		DEC8b10bERR,	-- "1101100111" 
		"000010111",	-- "1101101000", -D23.0-, [474,431]
		"000001001",	-- "1101101001", +D9.0-, [475,432]
		"000001010",	-- "1101101010", +D10.0-, [476,433]
		DEC8b10bERR,	-- "1101101011" 
		"000001100",	-- "1101101100", +D12.0-, [477,434]
		DEC8b10bERR,	-- "1101101101" 
		DEC8b10bERR,	-- "1101101110" 
		DEC8b10bERR,	-- "1101101111" 
		DEC8b10bERR,	-- "1101110000" 
		"000010001",	-- "1101110001", +D17.0-, [478,435]
		"000010010",	-- "1101110010", +D18.0-, [479,436]
		DEC8b10bERR,	-- "1101110011" 
		"000010100",	-- "1101110100", +D20.0-, [480,437]
		DEC8b10bERR,	-- "1101110101" 
		DEC8b10bERR,	-- "1101110110" 
		DEC8b10bERR,	-- "1101110111" 
		DEC8b10bERR,	-- "1101111000" 
		DEC8b10bERR,	-- "1101111001" 
		DEC8b10bERR,	-- "1101111010" 
		DEC8b10bERR,	-- "1101111011" 
		DEC8b10bERR,	-- "1101111100" 
		DEC8b10bERR,	-- "1101111101" 
		DEC8b10bERR,	-- "1101111110" 
		DEC8b10bERR,	-- "1101111111" 
		DEC8b10bERR,	-- "1110000000" 
		DEC8b10bERR,	-- "1110000001" 
		DEC8b10bERR,	-- "1110000010" 
		"111111100",	-- "1110000011", -K28.7-, [481,44]
		DEC8b10bERR,	-- "1110000100" 
		"111101111",	-- "1110000101", -K15.7-, [482,45]
		"111100000",	-- "1110000110", -K0.7-, [483,46]
		"111100111",	-- "1110000111", +K7.7-, [484,47]
		DEC8b10bERR,	-- "1110001000" 
		"111110000",	-- "1110001001", -K16.7-, [485,48]
		"111111111",	-- "1110001010", -K31.7-, [486,49]
		"111101011",	-- "1110001011", +K11.7-, [487,50]
		"111111000",	-- "1110001100", -K24.7-, [488,51]
		"111101101",	-- "1110001101", +K13.7-, [489,52]
		"111101110",	-- "1110001110", +K14.7-, [490,53]
		DEC8b10bERR,	-- "1110001111" 
		DEC8b10bERR,	-- "1110010000" 
		"111100001",	-- "1110010001", -K1.7-, [491,54]
		"111100010",	-- "1110010010", -K2.7-, [492,55]
		"111110011",	-- "1110010011", +K19.7-, [493,56]
		"111100100",	-- "1110010100", -K4.7-, [494,57]
		"111110101",	-- "1110010101", +K21.7-, [495,58]
		"111110110",	-- "1110010110", +K22.7-, [496,59]
		DEC8b10bERR,	-- "1110010111" 
		"111101000",	-- "1110011000", -K8.7-, [497,60]
		"111111001",	-- "1110011001", +K25.7-, [498,61]
		"111111010",	-- "1110011010", +K26.7-, [499,62]
		DEC8b10bERR,	-- "1110011011" 
		DEC8b10bERR,	-- "1110011100" 
		DEC8b10bERR,	-- "1110011101" 
		DEC8b10bERR,	-- "1110011110" 
		DEC8b10bERR,	-- "1110011111" 
		DEC8b10bERR,	-- "1110100000" 
		"111111110",	-- "1110100001", -K30.7-, [500,63]
		"111111101",	-- "1110100010", -K29.7-, [501,64]
		"111100011",	-- "1110100011", +K3.7-, [502,65]
		"111111011",	-- "1110100100", -K27.7-, [503,66]
		"111100101",	-- "1110100101", +K5.7-, [504,67]
		"111100110",	-- "1110100110", +K6.7-, [505,68]
		DEC8b10bERR,	-- "1110100111" 
		"111110111",	-- "1110101000", -K23.7-, [506,69]
		"111101001",	-- "1110101001", +K9.7-, [507,70]
		"111101010",	-- "1110101010", +K10.7-, [508,71]
		DEC8b10bERR,	-- "1110101011" 
		"111101100",	-- "1110101100", +K12.7-, [509,72]
		DEC8b10bERR,	-- "1110101101" 
		DEC8b10bERR,	-- "1110101110" 
		DEC8b10bERR,	-- "1110101111" 
		DEC8b10bERR,	-- "1110110000" 
		"011110001",	-- "1110110001", +D17.7-, [510,438]
		"011110010",	-- "1110110010", +D18.7-, [511,439]
		DEC8b10bERR,	-- "1110110011" 
		"011110100",	-- "1110110100", +D20.7-, [512,440]
		DEC8b10bERR,	-- "1110110101" 
		DEC8b10bERR,	-- "1110110110" 
		DEC8b10bERR,	-- "1110110111" 
		DEC8b10bERR,	-- "1110111000" 
		DEC8b10bERR,	-- "1110111001" 
		DEC8b10bERR,	-- "1110111010" 
		DEC8b10bERR,	-- "1110111011" 
		DEC8b10bERR,	-- "1110111100" 
		DEC8b10bERR,	-- "1110111101" 
		DEC8b10bERR,	-- "1110111110" 
		DEC8b10bERR,	-- "1110111111" 
		DEC8b10bERR,	-- "1111000000" 
		DEC8b10bERR,	-- "1111000001" 
		DEC8b10bERR,	-- "1111000010" 
		DEC8b10bERR,	-- "1111000011" 
		DEC8b10bERR,	-- "1111000100" 
		DEC8b10bERR,	-- "1111000101" 
		DEC8b10bERR,	-- "1111000110" 
		DEC8b10bERR,	-- "1111000111" 
		DEC8b10bERR,	-- "1111001000" 
		DEC8b10bERR,	-- "1111001001" 
		DEC8b10bERR,	-- "1111001010" 
		DEC8b10bERR,	-- "1111001011" 
		DEC8b10bERR,	-- "1111001100" 
		DEC8b10bERR,	-- "1111001101" 
		DEC8b10bERR,	-- "1111001110" 
		DEC8b10bERR,	-- "1111001111" 
		DEC8b10bERR,	-- "1111010000" 
		DEC8b10bERR,	-- "1111010001" 
		DEC8b10bERR,	-- "1111010010" 
		DEC8b10bERR,	-- "1111010011" 
		DEC8b10bERR,	-- "1111010100" 
		DEC8b10bERR,	-- "1111010101" 
		DEC8b10bERR,	-- "1111010110" 
		DEC8b10bERR,	-- "1111010111" 
		DEC8b10bERR,	-- "1111011000" 
		DEC8b10bERR,	-- "1111011001" 
		DEC8b10bERR,	-- "1111011010" 
		DEC8b10bERR,	-- "1111011011" 
		DEC8b10bERR,	-- "1111011100" 
		DEC8b10bERR,	-- "1111011101" 
		DEC8b10bERR,	-- "1111011110" 
		DEC8b10bERR,	-- "1111011111" 
		DEC8b10bERR,	-- "1111100000" 
		DEC8b10bERR,	-- "1111100001" 
		DEC8b10bERR,	-- "1111100010" 
		DEC8b10bERR,	-- "1111100011" 
		DEC8b10bERR,	-- "1111100100" 
		DEC8b10bERR,	-- "1111100101" 
		DEC8b10bERR,	-- "1111100110" 
		DEC8b10bERR,	-- "1111100111" 
		DEC8b10bERR,	-- "1111101000" 
		DEC8b10bERR,	-- "1111101001" 
		DEC8b10bERR,	-- "1111101010" 
		DEC8b10bERR,	-- "1111101011" 
		DEC8b10bERR,	-- "1111101100" 
		DEC8b10bERR,	-- "1111101101" 
		DEC8b10bERR,	-- "1111101110" 
		DEC8b10bERR,	-- "1111101111" 
		DEC8b10bERR,	-- "1111110000" 
		DEC8b10bERR,	-- "1111110001" 
		DEC8b10bERR,	-- "1111110010" 
		DEC8b10bERR,	-- "1111110011" 
		DEC8b10bERR,	-- "1111110100" 
		DEC8b10bERR,	-- "1111110101" 
		DEC8b10bERR,	-- "1111110110" 
		DEC8b10bERR,	-- "1111110111" 
		DEC8b10bERR,	-- "1111111000" 
		DEC8b10bERR,	-- "1111111001" 
		DEC8b10bERR,	-- "1111111010" 
		DEC8b10bERR,	-- "1111111011" 
		DEC8b10bERR,	-- "1111111100" 
		DEC8b10bERR,	-- "1111111101" 
		DEC8b10bERR,	-- "1111111110" 
		DEC8b10bERR 	-- "1111111111" 
	);


signal DECODE : std_logic_vector (8 downto 0);

begin

	CTRL_OUT <= DECODE(8);
	DATA_OUT <= DECODE(7 downto 0);
	
	process (CLK_IN)
	begin
		if(CLK_IN = '1' and CLK_IN'event)
		then
			DECODE <= TBL_DEC8B10B(conv_integer(ENCODE_IN));
		end if;
	end process;

end RTL;

