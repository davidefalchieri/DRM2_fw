-- Company:              CAEN SpA - Viareggio - Italy
-- Model:                   VX1392 -  ALICE Local Triiger Module
-- FPGA Proj. Name: vx1392ltm
-- Device:                 Actel APA600
-- Author:                  Colombini
-- Date:                     10:23:49 16/01/2008
-- ----------------------------------------------------------------------------
-- Module:         
-- Description:     
-- ****************************************************************************
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.2 (Build 37)

-- ############################################################################
-- Revision History:
-- ############################################################################
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE work.v1392pkg.all;

LIBRARY ltm_libr;

ENTITY v1392ltm IS
   PORT( 
      ALICLK      : IN     std_logic;
      AMB         : IN     std_logic_vector ( 5 DOWNTO 0);
      ASB         : IN     std_logic;
      BERRVME     : IN     std_logic;
      BNCRES      : IN     std_logic;
      DS0B        : IN     std_logic;
      DS1B        : IN     std_logic;
      EVRES       : IN     std_logic;
      F_SO        : IN     std_logic;
      GA          : IN     std_logic_vector ( 3 DOWNTO 0);
      IACKB       : IN     std_logic;
      IACKINB     : IN     std_logic;
      L0          : IN     std_logic;
      L1A         : IN     std_logic;
      L1R         : IN     std_logic;
      L2A         : IN     std_logic;
      L2R         : IN     std_logic;
      LCLK        : IN     std_logic;
      LOS         : IN     std_logic;
      NLBPCKE     : IN     std_logic;
      NLBPCKR     : IN     std_logic;
      NPWON       : IN     std_logic;
      PSM_SP0     : IN     std_logic;
      PSM_SP1     : IN     std_logic;
      PSM_SP2     : IN     std_logic;
      PSM_SP3     : IN     std_logic;
      PSM_SP4     : IN     std_logic;
      PSM_SP5     : IN     std_logic;
      SPULSE0     : IN     std_logic;
      SPULSE1     : IN     std_logic;
      SPULSE2     : IN     std_logic;
      SYSRESB     : IN     std_logic;
      WRITEB      : IN     std_logic;
      nLBRDY      : IN     std_logic;                       -- Pilotaggio led rosso vicino a conn. TDC (su pannello)
      ADLTC       : OUT    std_logic;
      AE_PDL      : OUT    std_logic_vector (47 DOWNTO 0);
      APACLK0     : OUT    std_logic;
      DIR_CTTM    : OUT    std_logic_vector (7 DOWNTO 0);
      FCS         : OUT    std_logic;
      F_SCK       : OUT    std_logic;
      F_SI        : OUT    std_logic;
      IACKOUTB    : OUT    std_logic;
      INTR1       : OUT    std_logic;
      INTR2       : OUT    std_logic;
      LED         : OUT    display_stream;
      LTM_BUSY    : OUT    std_logic;
      LTM_DRDY    : OUT    std_logic;
      MD_PDL      : OUT    std_logic;
      MYBERR      : OUT    std_logic;
      NDTKIN      : OUT    std_logic;
      NLBCLR      : OUT    std_logic;
      NLBCS       : OUT    std_logic;
      NLBRD       : OUT    std_logic;
      NLBRES      : OUT    std_logic;
      NLBWAIT     : OUT    std_logic;
      NOE16R      : OUT    std_logic;
      NOE16W      : OUT    std_logic;
      NOE32R      : OUT    std_logic;
      NOE32W      : OUT    std_logic;
      NOE64R      : OUT    std_logic;
      NOEAD       : OUT    std_logic;
      NOEDTK      : OUT    std_logic;                       -- Pilotaggio led verde vicino a conn. TDC (su pannello)
      NSELCLK     : OUT    std_logic;
      PSM_RES     : OUT    std_logic;
      P_PDL       : OUT    std_logic_vector (7 DOWNTO 1);
      RSELA0      : OUT    std_logic;
      RSELA1      : OUT    std_logic;
      RSELB0      : OUT    std_logic;
      RSELB1      : OUT    std_logic;
      RSELC0      : OUT    std_logic;
      RSELC1      : OUT    std_logic;
      RSELD0      : OUT    std_logic;
      RSELD1      : OUT    std_logic;
      SCL0        : OUT    std_logic;
      SCL1        : OUT    std_logic;
      SCLK_DAC    : OUT    std_logic;
      SCLK_PDL    : OUT    std_logic;
      SDIN_DAC    : OUT    std_logic;
      SELCLK      : OUT    std_logic;
      SI_PDL      : OUT    std_logic;
      SYNC        : OUT    std_logic_vector (15 DOWNTO 0);
      TST         : OUT    std_logic_vector (15 DOWNTO 0);
      nLBAS       : OUT    std_logic;                       -- Pilotaggio led rosso vicino a conn. TDC (su pannello)
      LB          : INOUT  std_logic_vector (31 DOWNTO 0);
      LBSP        : INOUT  std_logic_vector (31 DOWNTO 0);
      LWORDB      : INOUT  std_logic;
      NCYC_RELOAD : INOUT  std_logic;
      NLBLAST     : INOUT  std_logic;
      SDA0        : INOUT  std_logic;
      SDA1        : INOUT  std_logic;
      SP_PDL      : INOUT  std_logic_vector (47 DOWNTO 0);
      VAD         : INOUT  std_logic_vector (31 DOWNTO 1);
      VDB         : INOUT  std_logic_vector (31 DOWNTO 0)
   );

-- Declarations

END v1392ltm ;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE work.v1392pkg.all;


ARCHITECTURE struct OF v1392ltm IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL ACLK        : std_logic;
   SIGNAL BNC_RES     : std_logic;
   SIGNAL CHANNEL     : std_logic_vector(2 DOWNTO 0);
   SIGNAL CHIP_ADDR   : std_logic_vector(2 DOWNTO 0);
   SIGNAL CLEAR       : std_logic;
   SIGNAL CLK         : std_logic;
   SIGNAL CROMWAD     : std_logic_vector(8 DOWNTO 0);
   SIGNAL CROMWDT     : std_logic_vector(7 DOWNTO 0);
   SIGNAL DACCFG_DT   : std_logic_vector(15 DOWNTO 0);
   SIGNAL DACCFG_RAD  : std_logic_vector( 3 DOWNTO 0);
   SIGNAL DACCFG_WAD  : std_logic_vector( 3 DOWNTO 0);
   SIGNAL DACCFG_WDT  : std_logic_vector(15 DOWNTO 0);
   SIGNAL DACCFG_nRD  : std_logic;
   SIGNAL DACCFG_nWR  : std_logic;
   SIGNAL DAC_REFRESH : std_logic;
   SIGNAL DEBUG       : debug_stream;
   SIGNAL DL7         : std_logic;                        -- Pilotaggio led rosso vicino a ALICLK (su pannello)
   SIGNAL DPR         : std_logic_vector(31 DOWNTO 0);
   SIGNAL DPR_P       : std_logic_vector(3 DOWNTO 0);
   SIGNAL DTEST_FIFO  : std_logic;
   SIGNAL EF          : std_logic;
   SIGNAL EVRDY       : std_logic;
   SIGNAL EVREAD      : std_logic;
   SIGNAL EV_RES      : std_logic;
   SIGNAL FBOUT       : std_logic_vector(7 DOWNTO 0);
   SIGNAL FF          : std_logic;
   SIGNAL FWIMG2LOAD  : std_logic;
   SIGNAL HWCLEAR     : std_logic;
   SIGNAL HWRES       : std_logic;
   SIGNAL I2C_CHAIN   : std_logic;
   SIGNAL I2C_RACK    : std_logic;
   SIGNAL I2C_RDATA   : std_logic_vector(9 DOWNTO 0);
   SIGNAL I2C_RREQ    : std_logic;
   SIGNAL LOAD_RES    : std_logic;
   SIGNAL NRDMEB      : std_logic;
   SIGNAL OR_RACK     : std_logic;
   SIGNAL OR_RADDR    : std_logic_vector(5 DOWNTO 0);
   SIGNAL OR_RDATA    : std_logic_vector(9 DOWNTO 0);
   SIGNAL OR_RREQ     : std_logic;
   SIGNAL PAE         : std_logic;
   SIGNAL PAF         : std_logic;
   SIGNAL PDLCFG_DT   : std_logic_vector(7 DOWNTO 0);
   SIGNAL PDLCFG_RAD  : std_logic_vector(5 DOWNTO 0);
   SIGNAL PDLCFG_WAD  : std_logic_vector(5 DOWNTO 0);
   SIGNAL PDLCFG_WDT  : std_logic_vector(7 DOWNTO 0);
   SIGNAL PDLCFG_nRD  : std_logic;
   SIGNAL PDLCFG_nWR  : std_logic;
   SIGNAL PDL_RACK    : std_logic;
   SIGNAL PDL_RADDR   : std_logic_vector(5 DOWNTO 0);
   SIGNAL PDL_RDATA   : std_logic_vector(7 DOWNTO 0);
   SIGNAL PDL_RREQ    : std_logic;
   SIGNAL PON_LOAD    : std_logic;
   SIGNAL PULSE       : reg_pulse;
   SIGNAL RAMAD_VME   : std_logic_vector(8 DOWNTO 0);
   SIGNAL RAMDT       : std_logic_vector(7 DOWNTO 0);
   SIGNAL RAMRD       : std_logic;
   SIGNAL REG         : reg_stream;
   SIGNAL RUN         : std_logic;
   SIGNAL SM_SIDE     : std_logic;
   SIGNAL TICK        : tick_pulses;
   SIGNAL TRIGLED     : std_logic;
   SIGNAL VDD         : std_logic;
   SIGNAL WDOGTO      : std_logic;
   SIGNAL WRCROM      : std_logic;
   SIGNAL dout        : std_logic;
   SIGNAL dout1       : std_logic;

   -- Implicit buffer signal declarations
   SIGNAL NOEDTK_internal : std_logic;

   -- Component Declarations
   COMPONENT CLK_INTERF
   PORT (
      CLK     : IN     std_logic;
      HWRES   : IN     std_logic;
      LOS     : IN     std_logic;
      PULSE   : IN     reg_pulse;
      TICK    : IN     tick_pulses;
      NSELCLK : OUT    std_logic;
      RSELA0  : OUT    std_logic;
      RSELA1  : OUT    std_logic;
      RSELB0  : OUT    std_logic;
      RSELB1  : OUT    std_logic;
      RSELC0  : OUT    std_logic;
      RSELC1  : OUT    std_logic;
      RSELD0  : OUT    std_logic;
      RSELD1  : OUT    std_logic;
      SELCLK  : OUT    std_logic;
      DEBUG   : INOUT  debug_stream;
      REG     : INOUT  reg_stream
   );
   END COMPONENT;
   COMPONENT CROM
   PORT (
      DI     : IN     std_logic_vector (7 DOWNTO 0);
      RADDR  : IN     std_logic_vector (8 DOWNTO 0);
      RCLOCK : IN     std_logic;
      RDB    : IN     std_logic;
      WADDR  : IN     std_logic_vector (8 DOWNTO 0);
      WCLOCK : IN     std_logic;
      WRB    : IN     std_logic;
      DO     : OUT    std_logic_vector (7 DOWNTO 0);
      PO     : OUT    std_logic
   );
   END COMPONENT;
   COMPONENT DACCFG
   PORT (
      DI     : IN     std_logic_vector (15 DOWNTO 0);
      RADDR  : IN     std_logic_vector (3 DOWNTO 0);
      RCLOCK : IN     std_logic;
      RDB    : IN     std_logic;
      WADDR  : IN     std_logic_vector (3 DOWNTO 0);
      WCLOCK : IN     std_logic;
      WRB    : IN     std_logic;
      DO     : OUT    std_logic_vector (15 DOWNTO 0);
      PO     : OUT    std_logic_vector (1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT DAC_INTERF
   GENERIC (
      G_SIM_ON : boolean      -- Fast SPI
   );
   PORT (
      CLK         : IN     std_logic;
      DACCFG_DT   : IN     std_logic_vector (15 DOWNTO 0);
      DAC_REFRESH : IN     std_logic;
      HWRES       : IN     std_logic;
      PULSE       : IN     reg_pulse;
      TICK        : IN     tick_pulses;
      DACCFG_RAD  : OUT    std_logic_vector ( 3 DOWNTO 0);
      DACCFG_nRD  : OUT    std_logic;
      SCLK_DAC    : OUT    std_logic;
      SDIN_DAC    : OUT    std_logic;
      SYNC        : OUT    std_logic_vector (15 DOWNTO 0);
      DEBUG       : INOUT  debug_stream;
      REG         : INOUT  reg_stream
   );
   END COMPONENT;
   COMPONENT I2C_INTERF_LTM
   PORT (
      CHANNEL   : IN     std_logic_vector (2 DOWNTO 0);
      CHIP_ADDR : IN     std_logic_vector (2 DOWNTO 0);
      CLK       : IN     std_logic;
      HWRES     : IN     std_logic;
      I2C_CHAIN : IN     std_logic;
      I2C_RREQ  : IN     std_logic;
      PULSE     : IN     reg_pulse;
      TICK      : IN     tick_pulses;
      I2C_RACK  : OUT    std_logic;
      I2C_RDATA : OUT    std_logic_vector (9 DOWNTO 0);
      SCLA      : OUT    std_logic;
      SCLB      : OUT    std_logic;
      DEBUG     : INOUT  debug_stream;
      REG       : INOUT  reg_stream;
      SDAA      : INOUT  std_logic;
      SDAB      : INOUT  std_logic
   );
   END COMPONENT;
   COMPONENT PDLCFG
   PORT (
      DI     : IN     std_logic_vector (7 DOWNTO 0);
      RADDR  : IN     std_logic_vector (5 DOWNTO 0);
      RCLOCK : IN     std_logic;
      RDB    : IN     std_logic;
      WADDR  : IN     std_logic_vector (5 DOWNTO 0);
      WCLOCK : IN     std_logic;
      WRB    : IN     std_logic;
      DO     : OUT    std_logic_vector (7 DOWNTO 0);
      PO     : OUT    std_logic
   );
   END COMPONENT;
   COMPONENT RESET_MOD
   GENERIC (
      G_SIM_ON : boolean      -- TRUE=Fast simulation
   );
   PORT (
      ACLK      : IN     std_logic;
      BNC_RESIN : IN     std_logic;
      CLK       : IN     std_logic;
      EV_RESIN  : IN     std_logic;
      LOAD_RES  : IN     std_logic;
      NPWON     : IN     std_logic;
      PULSE     : IN     reg_pulse;
      SYSRESB   : IN     std_logic;
      WDOGTO    : IN     std_logic;
      BNC_RES   : OUT    std_logic;
      CLEAR     : OUT    std_logic;
      EV_RES    : OUT    std_logic;
      HWCLEAR   : OUT    std_logic;
      HWRES     : OUT    std_logic;
      PON_LOAD  : OUT    std_logic;
      RUN       : OUT    std_logic;
      TICK      : OUT    tick_pulses;
      DEBUG     : INOUT  debug_stream;
      REG       : INOUT  reg_stream
   );
   END COMPONENT;
   COMPONENT ROC32
   GENERIC (
      SimCfg_NoADCEvent : boolean
   );
   PORT (
      ACLK        : IN     std_logic;
      BNC_RES     : IN     std_logic;
      CLEAR       : IN     std_logic;
      CLK         : IN     std_logic;
      EVREAD      : IN     std_logic;
      GA          : IN     std_logic_vector ( 3 DOWNTO 0);
      HWRES       : IN     std_logic;
      I2C_RACK    : IN     std_logic;
      I2C_RDATA   : IN     std_logic_vector (9 DOWNTO 0);
      L0          : IN     std_logic;
      L1A         : IN     std_logic;
      L1R         : IN     std_logic;
      L2A         : IN     std_logic;
      L2R         : IN     std_logic;
      NRDMEB      : IN     std_logic;
      OR_RACK     : IN     std_logic;
      OR_RDATA    : IN     std_logic_vector (9 DOWNTO 0);
      PDL_RACK    : IN     std_logic;
      PDL_RDATA   : IN     std_logic_vector (7 DOWNTO 0);
      PSM_SP0     : IN     std_logic;
      PSM_SP1     : IN     std_logic;
      PSM_SP2     : IN     std_logic;
      PSM_SP3     : IN     std_logic;
      PSM_SP4     : IN     std_logic;
      PSM_SP5     : IN     std_logic;
      PULSE       : IN     reg_pulse;
      SPULSE0     : IN     std_logic;
      SPULSE1     : IN     std_logic;
      SPULSE2     : IN     std_logic;
      TICK        : IN     tick_pulses;
      CHANNEL     : OUT    std_logic_vector (2 DOWNTO 0);
      CHIP_ADDR   : OUT    std_logic_vector (2 DOWNTO 0);
      DAC_REFRESH : OUT    std_logic;
      DPR         : OUT    std_logic_vector (31 DOWNTO 0);
      DPR_P       : OUT    std_logic_vector ( 3 DOWNTO 0);
      DTEST_FIFO  : OUT    std_logic;
      EF          : OUT    std_logic;
      EVRDY       : OUT    std_logic;
      I2C_CHAIN   : OUT    std_logic;
      I2C_RREQ    : OUT    std_logic;
      LTM_BUSY    : OUT    std_logic;
      LTM_DRDY    : OUT    std_logic;
      OR_RADDR    : OUT    std_logic_vector (5 DOWNTO 0);
      OR_RREQ     : OUT    std_logic;
      PAE         : OUT    std_logic;
      PAF         : OUT    std_logic;
      PDL_RADDR   : OUT    std_logic_vector (5 DOWNTO 0);
      PDL_RREQ    : OUT    std_logic;
      TRIGLED     : OUT    std_logic;
      ff          : OUT    std_logic;
      DEBUG       : INOUT  debug_stream;
      REG         : INOUT  reg_stream
   );
   END COMPONENT;
   COMPONENT SPI_INTERF
   GENERIC (
      G_SIM_ON       : boolean;      -- Fast SPI
      G_LOAD_DISABLE : boolean       -- Disable CRAM load
   );
   PORT (
      CLK         : IN     std_logic;
      FWIMG2LOAD  : IN     std_logic;
      F_SO        : IN     std_logic;
      HWCLEAR     : IN     std_logic;
      HWRES       : IN     std_logic;
      PON_LOAD    : IN     std_logic;
      PULSE       : IN     reg_pulse;
      TICK        : IN     tick_pulses;
      CROMWAD     : OUT    std_logic_vector (8 DOWNTO 0);
      CROMWDT     : OUT    std_logic_vector (7 DOWNTO 0);
      DACCFG_WAD  : OUT    std_logic_vector ( 3 DOWNTO 0);
      DACCFG_WDT  : OUT    std_logic_vector (15 DOWNTO 0);
      DACCFG_nWR  : OUT    std_logic;
      FBOUT       : OUT    std_logic_vector (7 DOWNTO 0);
      FCS         : OUT    std_logic;
      F_SCK       : OUT    std_logic;
      F_SI        : OUT    std_logic;
      LOAD_RES    : OUT    std_logic;
      PDLCFG_WAD  : OUT    std_logic_vector (5 DOWNTO 0);
      PDLCFG_WDT  : OUT    std_logic_vector (7 DOWNTO 0);
      PDLCFG_nWR  : OUT    std_logic;
      WRCROM      : OUT    std_logic;
      DEBUG       : INOUT  debug_stream;
      REG         : INOUT  reg_stream;
      nCYC_RELOAD : INOUT  std_logic
   );
   END COMPONENT;
   COMPONENT VINTERF
   PORT (
      ALICLK     : IN     std_logic;
      AMB        : IN     std_logic_vector ( 5 DOWNTO 0);
      ASB        : IN     std_logic;
      BERRVME    : IN     std_logic;
      CLEAR      : IN     std_logic;
      CLK        : IN     std_logic;
      DPR        : IN     std_logic_vector (31 DOWNTO 0);
      DPR_P      : IN     std_logic_vector ( 3 DOWNTO 0);
      DS0B       : IN     std_logic;
      DS1B       : IN     std_logic;
      DTEST_FIFO : IN     std_logic;
      EF         : IN     std_logic;
      EVRDY      : IN     std_logic;
      FBOUT      : IN     std_logic_vector (7 DOWNTO 0);
      GA         : IN     std_logic_vector ( 3 DOWNTO 0);
      HWCLEAR    : IN     std_logic;
      HWRES      : IN     std_logic;
      IACKB      : IN     std_logic;
      IACKINB    : IN     std_logic;
      LBSP       : IN     std_logic_vector (31 DOWNTO 0);
      OR_RADDR   : IN     std_logic_vector (5 DOWNTO 0);
      OR_RREQ    : IN     std_logic;
      PAE        : IN     std_logic;
      PAF        : IN     std_logic;
      RAMDT      : IN     std_logic_vector (7 DOWNTO 0);
      TICK       : IN     tick_pulses;
      WRITEB     : IN     std_logic;
      ff         : IN     std_logic;
      nLBPCKE    : IN     std_logic;
      nLBPCKR    : IN     std_logic;
      nLBRDY     : IN     std_logic;
      ADLTC      : OUT    std_logic;
      EVREAD     : OUT    std_logic;
      FWIMG2LOAD : OUT    std_logic;
      IACKOUTB   : OUT    std_logic;
      INTR1      : OUT    std_logic;
      INTR2      : OUT    std_logic;
      MYBERR     : OUT    std_logic;
      NDTKIN     : OUT    std_logic;
      NOE16R     : OUT    std_logic;
      NOE16W     : OUT    std_logic;
      NOE32R     : OUT    std_logic;
      NOE32W     : OUT    std_logic;
      NOE64R     : OUT    std_logic;
      NOEAD      : OUT    std_logic;
      NOEDTK     : OUT    std_logic;
      NRDMEB     : OUT    std_logic;
      OR_RACK    : OUT    std_logic;
      OR_RDATA   : OUT    std_logic_vector (9 DOWNTO 0);
      PULSE      : OUT    reg_pulse;
      RAMAD_VME  : OUT    std_logic_vector (8 DOWNTO 0);
      RAMRD      : OUT    std_logic;
      SM_SIDE    : OUT    std_logic;
      WDOGTO     : OUT    std_logic;
      nLBAS      : OUT    std_logic;
      nLBCLR     : OUT    std_logic;
      nLBCS      : OUT    std_logic;
      nLBLAST    : OUT    std_logic;
      nLBRD      : OUT    std_logic;
      nLBRES     : OUT    std_logic;
      nLBWAIT    : OUT    std_logic;
      DEBUG      : INOUT  debug_stream;
      LB         : INOUT  std_logic_vector (31 DOWNTO 0);
      LWORDB     : INOUT  std_logic;
      REG        : INOUT  reg_stream;
      VAD        : INOUT  std_logic_vector (31 DOWNTO 1);
      VDB        : INOUT  std_logic_vector (31 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT ctrl
   PORT (
      HWRES    : IN     std_logic ;
      CLK      : IN     std_logic ;
      DL1      : IN     std_logic ;                    -- Pilotaggio led rosso vicino a conn. TDC (su pannello)
      DL2      : IN     std_logic ;                    -- Pilotaggio led verde vicino a conn. TDC (su pannello)
      DL5      : IN     std_logic ;                    -- Pilotaggio led verde vicino a CTTM (non visibile su pannello)
      DL6      : IN     std_logic ;                    -- Pilotaggio led giallo vicino a CTTM (non visibile su pannello)
      DL7      : IN     std_logic ;                    -- Pilotaggio led rosso vicino a ALICLK (su pannello)
      DL8      : IN     std_logic ;                    -- Pilotaggio led giallo vicino a ALICLK (su pannello)
      DIR_CTTM : OUT    std_logic_vector (7 DOWNTO 0); -- CTTM LVDS Buffers dir ('0' = RX, '1' = TX)
      LED      : OUT    std_logic_vector (5 DOWNTO 0); -- LED driver
      PSM_RES  : OUT    std_logic ;                    -- Reset micro (active high)
      SP       : OUT    std_logic_vector (5 DOWNTO 0); -- Spare conn. w/ micro
      REG      : INOUT  reg_stream ;
      PULSE    : IN     reg_pulse ;
      DEBUG    : INOUT  debug_stream ;
      TICK     : IN     tick_pulses 
   );
   END COMPONENT;
   COMPONENT lbspare
   PORT (
      BNC_RES : IN     std_logic;
      EV_RES  : IN     std_logic;
      L0      : IN     std_logic;
      L1A     : IN     std_logic;
      L1R     : IN     std_logic;
      L2A     : IN     std_logic;
      L2R     : IN     std_logic;
      LOS     : IN     std_logic;
      RUN     : IN     std_logic;
      SM_SIDE : IN     std_logic;
      SPULSE0 : IN     std_logic;
      SPULSE1 : IN     std_logic;
      SPULSE2 : IN     std_logic;
      LBSP    : INOUT  std_logic_vector (31 DOWNTO 0);
      REG     : INOUT  reg_stream
   );
   END COMPONENT;
   COMPONENT pdl_interf
   PORT (
      CLEAR      : IN     std_logic;
      CLK        : IN     std_logic;
      HWRES      : IN     std_logic;
      LOAD_RES   : IN     std_logic;
      PDLCFG_DT  : IN     std_logic_vector (7 DOWNTO 0);
      PDL_RADDR  : IN     std_logic_vector (5 DOWNTO 0);
      PDL_RREQ   : IN     std_logic;
      PULSE      : IN     reg_pulse;
      TICK       : IN     tick_pulses;
      AE         : OUT    std_logic_vector (47 DOWNTO 0);
      MD         : OUT    std_logic;
      P          : OUT    std_logic_vector (7 DOWNTO 1);
      PDLCFG_RAD : OUT    std_logic_vector (5 DOWNTO 0);
      PDLCFG_nRD : OUT    std_logic;
      PDL_RACK   : OUT    std_logic;
      PDL_RDATA  : OUT    std_logic_vector (7 DOWNTO 0);
      SC         : OUT    std_logic;
      si         : OUT    std_logic;
      DEBUG      : INOUT  debug_stream;
      REG        : INOUT  reg_stream;
      SP0        : INOUT  std_logic_vector (47 DOWNTO 0)
   );
   END COMPONENT;


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 eb1
   -- eb1 1
   TST(0) <= DEBUG(0); 
   TST(1) <= DEBUG(1);
   TST(2) <= DEBUG(2);
   TST(3) <= DEBUG(3);
   TST(4) <= DEBUG(4);
   TST(5) <= DEBUG(5);
   TST(6) <= DEBUG(6);
   TST(7) <= DEBUG(7);
   TST(8) <= DEBUG(8);
   TST(9) <= DEBUG(9);
   TST(10) <= DEBUG(10);
   TST(11) <= DEBUG(11);
   TST(12) <= DEBUG(12);
   TST(13) <= DEBUG(13);
   TST(14) <= DEBUG(14);
   TST(15) <= DEBUG(15);


   -- ModuleWare code(v1.7) for instance 'I17' of 'inv'
   DL7 <= NOT(RUN);

   -- ModuleWare code(v1.7) for instance 'I19' of 'inv'
   dout1 <= NOT(TRIGLED);

   -- ModuleWare code(v1.7) for instance 'I12' of 'pbuf'
   i12seq_proc: PROCESS (ALICLK)
   BEGIN
      IF (ALICLK ='1' ) THEN
         ACLK <= '1';
      ELSIF (ALICLK ='H' ) THEN
         ACLK <= '1';
      ELSIF (ALICLK ='0' ) THEN
         ACLK <= '0';
      ELSIF (ALICLK ='L' ) THEN
         ACLK <= '0';
      ELSIF (ALICLK ='U' ) THEN
         ACLK <= 'U';
      ELSIF (ALICLK ='X' ) THEN
         ACLK <= 'X';
      ELSIF (ALICLK ='Z' ) THEN
         ACLK <= 'X';
      END IF;
   END PROCESS i12seq_proc;

   -- ModuleWare code(v1.7) for instance 'I13' of 'pbuf'
   i13seq_proc: PROCESS (LCLK)
   BEGIN
      IF (LCLK ='1' ) THEN
         CLK <= '1';
      ELSIF (LCLK ='H' ) THEN
         CLK <= '1';
      ELSIF (LCLK ='0' ) THEN
         CLK <= '0';
      ELSIF (LCLK ='L' ) THEN
         CLK <= '0';
      ELSIF (LCLK ='U' ) THEN
         CLK <= 'U';
      ELSIF (LCLK ='X' ) THEN
         CLK <= 'X';
      ELSIF (LCLK ='Z' ) THEN
         CLK <= 'X';
      END IF;
   END PROCESS i13seq_proc;

   -- ModuleWare code(v1.7) for instance 'I15' of 'pbuf'
   i15seq_proc: PROCESS (CLK)
   BEGIN
      IF (CLK ='1' ) THEN
         APACLK0 <= '1';
      ELSIF (CLK ='H' ) THEN
         APACLK0 <= '1';
      ELSIF (CLK ='0' ) THEN
         APACLK0 <= '0';
      ELSIF (CLK ='L' ) THEN
         APACLK0 <= '0';
      ELSIF (CLK ='U' ) THEN
         APACLK0 <= 'U';
      ELSIF (CLK ='X' ) THEN
         APACLK0 <= 'X';
      ELSIF (CLK ='Z' ) THEN
         APACLK0 <= 'X';
      END IF;
   END PROCESS i15seq_proc;

   -- ModuleWare code(v1.7) for instance 'I4' of 'vdd'
   VDD <= '1';

   -- ModuleWare code(v1.7) for instance 'I18' of 'vdd'
   dout <= '1';

   -- Instance port mappings.
   I9 : CLK_INTERF
      PORT MAP (
         CLK     => CLK,
         HWRES   => HWRES,
         RSELA0  => RSELA0,
         RSELA1  => RSELA1,
         RSELB0  => RSELB0,
         RSELB1  => RSELB1,
         RSELC0  => RSELC0,
         RSELC1  => RSELC1,
         RSELD0  => RSELD0,
         RSELD1  => RSELD1,
         SELCLK  => SELCLK,
         NSELCLK => NSELCLK,
         LOS     => LOS,
         REG     => REG,
         PULSE   => PULSE,
         TICK    => TICK,
         DEBUG   => DEBUG
      );
   I6 : CROM
      PORT MAP (
         DO     => RAMDT,
         RCLOCK => CLK,
         WCLOCK => CLK,
         DI     => CROMWDT,
         PO     => OPEN,
         WRB    => WRCROM,
         RDB    => RAMRD,
         WADDR  => CROMWAD,
         RADDR  => RAMAD_VME
      );
   I14 : DACCFG
      PORT MAP (
         DO     => DACCFG_DT,
         RCLOCK => CLK,
         WCLOCK => CLK,
         DI     => DACCFG_WDT,
         PO     => OPEN,
         WRB    => DACCFG_nWR,
         RDB    => DACCFG_nRD,
         WADDR  => DACCFG_WAD,
         RADDR  => DACCFG_RAD
      );
   I8 : DAC_INTERF
      GENERIC MAP (
         G_SIM_ON => TRUE         -- Fast SPI  -- DAV (was FALSE)
      )
      PORT MAP (
         CLK         => CLK,
         HWRES       => HWRES,
         SYNC        => SYNC,
         SDIN_DAC    => SDIN_DAC,
         SCLK_DAC    => SCLK_DAC,
         DAC_REFRESH => DAC_REFRESH,
         DACCFG_nRD  => DACCFG_nRD,
         DACCFG_DT   => DACCFG_DT,
         DACCFG_RAD  => DACCFG_RAD,
         REG         => REG,
         PULSE       => PULSE,
         TICK        => TICK,
         DEBUG       => DEBUG
      );
   I1 : I2C_INTERF_LTM
      PORT MAP (
         CLK       => CLK,
         HWRES     => HWRES,
         SDAA      => SDA0,
         SCLA      => SCL0,
         SDAB      => SDA1,
         SCLB      => SCL1,
         I2C_RDATA => I2C_RDATA,
         I2C_RREQ  => I2C_RREQ,
         I2C_RACK  => I2C_RACK,
         I2C_CHAIN => I2C_CHAIN,
         CHIP_ADDR => CHIP_ADDR,
         CHANNEL   => CHANNEL,
         REG       => REG,
         PULSE     => PULSE,
         TICK      => TICK,
         DEBUG     => DEBUG
      );
   I11 : PDLCFG
      PORT MAP (
         DO     => PDLCFG_DT,
         RCLOCK => CLK,
         WCLOCK => CLK,
         DI     => PDLCFG_WDT,
         PO     => OPEN,
         WRB    => PDLCFG_nWR,
         RDB    => PDLCFG_nRD,
         WADDR  => PDLCFG_WAD,
         RADDR  => PDLCFG_RAD
      );
   I0 : RESET_MOD
      GENERIC MAP (
         G_SIM_ON => TRUE         -- TRUE=Fast simulation  -- DAV (was FALSE)
      )
      PORT MAP (
         CLK       => CLK,
         ACLK      => ACLK,
         NPWON     => NPWON,
         SYSRESB   => SYSRESB,
         LOAD_RES  => LOAD_RES,
         WDOGTO    => WDOGTO,
         HWRES     => HWRES,
         CLEAR     => CLEAR,
         HWCLEAR   => HWCLEAR,
         RUN       => RUN,
         PON_LOAD  => PON_LOAD,
         BNC_RESIN => BNCRES,
         EV_RESIN  => EVRES,
         BNC_RES   => BNC_RES,
         EV_RES    => EV_RES,
         DEBUG     => DEBUG,
         PULSE     => PULSE,
         REG       => REG,
         TICK      => TICK
      );
   I10 : ROC32
      GENERIC MAP (
         SimCfg_NoADCEvent => TRUE  -- FALSE (DAV)
      )
      PORT MAP (
         CLK         => CLK,
         ACLK        => ACLK,
         HWRES       => HWRES,
         CLEAR       => CLEAR,
         GA          => GA,
         L0          => L0,
         L1A         => L1A,
         L1R         => L1R,
         L2A         => L2A,
         L2R         => L2R,
         BNC_RES     => BNC_RES,
         SPULSE0     => SPULSE0,
         SPULSE1     => SPULSE1,
         SPULSE2     => SPULSE2,
         LTM_DRDY    => LTM_DRDY,
         LTM_BUSY    => LTM_BUSY,
         I2C_RDATA   => I2C_RDATA,
         I2C_RREQ    => I2C_RREQ,
         I2C_RACK    => I2C_RACK,
         I2C_CHAIN   => I2C_CHAIN,
         CHIP_ADDR   => CHIP_ADDR,
         CHANNEL     => CHANNEL,
         PDL_RDATA   => PDL_RDATA,
         PDL_RADDR   => PDL_RADDR,
         PDL_RREQ    => PDL_RREQ,
         PDL_RACK    => PDL_RACK,
         OR_RDATA    => OR_RDATA,
         OR_RADDR    => OR_RADDR,
         OR_RREQ     => OR_RREQ,
         OR_RACK     => OR_RACK,
         DAC_REFRESH => DAC_REFRESH,
         PSM_SP0     => PSM_SP0,
         PSM_SP1     => PSM_SP1,
         PSM_SP2     => PSM_SP2,
         PSM_SP3     => PSM_SP3,
         PSM_SP4     => PSM_SP4,
         PSM_SP5     => PSM_SP5,
         DPR         => DPR,
         DPR_P       => DPR_P,
         NRDMEB      => NRDMEB,
         PAF         => PAF,
         PAE         => PAE,
         EF          => EF,
         ff          => FF,
         EVRDY       => EVRDY,
         EVREAD      => EVREAD,
         TRIGLED     => TRIGLED,
         DEBUG       => DEBUG,
         DTEST_FIFO  => DTEST_FIFO,
         REG         => REG,
         TICK        => TICK,
         PULSE       => PULSE
      );
   I5 : SPI_INTERF
      GENERIC MAP (
         G_SIM_ON       => TRUE,         -- Fast SPI  -- DAV (was false)
         G_LOAD_DISABLE => FALSE          -- Disable CRAM load
      )
      PORT MAP (
         CLK         => CLK,
         HWRES       => HWRES,
         HWCLEAR     => HWCLEAR,
         FCS         => FCS,
         nCYC_RELOAD => NCYC_RELOAD,
         F_SI        => F_SI,
         F_SO        => F_SO,
         F_SCK       => F_SCK,
         FBOUT       => FBOUT,
         LOAD_RES    => LOAD_RES,
         PON_LOAD    => PON_LOAD,
         FWIMG2LOAD  => FWIMG2LOAD,
         CROMWAD     => CROMWAD,
         CROMWDT     => CROMWDT,
         WRCROM      => WRCROM,
         PDLCFG_nWR  => PDLCFG_nWR,
         PDLCFG_WAD  => PDLCFG_WAD,
         PDLCFG_WDT  => PDLCFG_WDT,
         DACCFG_nWR  => DACCFG_nWR,
         DACCFG_WAD  => DACCFG_WAD,
         DACCFG_WDT  => DACCFG_WDT,
         REG         => REG,
         PULSE       => PULSE,
         DEBUG       => DEBUG,
         TICK        => TICK
      );
   I2 : VINTERF
      PORT MAP (
         CLK        => CLK,
         ALICLK     => ALICLK,
         HWRES      => HWRES,
         CLEAR      => CLEAR,
         HWCLEAR    => HWCLEAR,
         WDOGTO     => WDOGTO,
         ASB        => ASB,
         DS0B       => DS0B,
         DS1B       => DS1B,
         WRITEB     => WRITEB,
         IACKB      => IACKB,
         IACKINB    => IACKINB,
         IACKOUTB   => IACKOUTB,
         NDTKIN     => NDTKIN,
         NOEDTK     => NOEDTK_internal,
         BERRVME    => BERRVME,
         MYBERR     => MYBERR,
         LWORDB     => LWORDB,
         VAD        => VAD,
         VDB        => VDB,
         AMB        => AMB,
         GA         => GA,
         INTR1      => INTR1,
         INTR2      => INTR2,
         ADLTC      => ADLTC,
         NOE16R     => NOE16R,
         NOE16W     => NOE16W,
         NOE32R     => NOE32R,
         NOE32W     => NOE32W,
         NOE64R     => NOE64R,
         NOEAD      => NOEAD,
         DPR        => DPR,
         DPR_P      => DPR_P,
         NRDMEB     => NRDMEB,
         PAF        => PAF,
         PAE        => PAE,
         EF         => EF,
         ff         => FF,
         OR_RDATA   => OR_RDATA,
         OR_RADDR   => OR_RADDR,
         OR_RREQ    => OR_RREQ,
         OR_RACK    => OR_RACK,
         RAMDT      => RAMDT,
         RAMAD_VME  => RAMAD_VME,
         RAMRD      => RAMRD,
         EVRDY      => EVRDY,
         EVREAD     => EVREAD,
         DTEST_FIFO => DTEST_FIFO,
         nLBAS      => nLBAS,
         nLBCLR     => NLBCLR,
         nLBCS      => NLBCS,
         nLBLAST    => NLBLAST,
         nLBRD      => NLBRD,
         nLBRES     => NLBRES,
         nLBWAIT    => NLBWAIT,
         nLBPCKE    => NLBPCKE,
         nLBPCKR    => NLBPCKR,
         nLBRDY     => nLBRDY,
         LB         => LB,
         LBSP       => LBSP,
         SM_SIDE    => SM_SIDE,
         FBOUT      => FBOUT,
         DEBUG      => DEBUG,
         FWIMG2LOAD => FWIMG2LOAD,
         REG        => REG,
         PULSE      => PULSE,
         TICK       => TICK
      );
   I7 : ctrl
      PORT MAP (
         HWRES    => HWRES,
         CLK      => CLK,
         DL1      => nLBRDY,
         DL2      => NOEDTK_internal,
         DL5      => dout,
         DL6      => dout,
         DL7      => DL7,
         DL8      => dout1,
         DIR_CTTM => DIR_CTTM,
         LED      => LED,
         PSM_RES  => PSM_RES,
         SP       => OPEN,
         REG      => REG,
         PULSE    => PULSE,
         DEBUG    => DEBUG,
         TICK     => TICK
      );
   I16 : lbspare
      PORT MAP (
         RUN     => RUN,
         LOS     => LOS,
         SM_SIDE => SM_SIDE,
         L0      => L0,
         L1A     => L1A,
         L1R     => L1R,
         L2A     => L2A,
         L2R     => L2R,
         BNC_RES => BNC_RES,
         EV_RES  => EV_RES,
         SPULSE0 => SPULSE0,
         SPULSE1 => SPULSE1,
         SPULSE2 => SPULSE2,
         LBSP    => LBSP,
         REG     => REG
      );
   I3 : pdl_interf
      PORT MAP (
         CLK        => CLK,
         HWRES      => HWRES,
         CLEAR      => CLEAR,
         LOAD_RES   => LOAD_RES,
         SP0        => SP_PDL,
         AE         => AE_PDL,
         si         => SI_PDL,
         SC         => SCLK_PDL,
         MD         => MD_PDL,
         P          => P_PDL,
         PDL_RDATA  => PDL_RDATA,
         PDL_RADDR  => PDL_RADDR,
         PDL_RREQ   => PDL_RREQ,
         PDL_RACK   => PDL_RACK,
         PDLCFG_nRD => PDLCFG_nRD,
         PDLCFG_DT  => PDLCFG_DT,
         PDLCFG_RAD => PDLCFG_RAD,
         DEBUG      => DEBUG,
         REG        => REG,
         PULSE      => PULSE,
         TICK       => TICK
      );

   -- Implicit buffered output assignments
   NOEDTK <= NOEDTK_internal;

END struct;
